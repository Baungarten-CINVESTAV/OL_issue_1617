magic
tech sky130A
magscale 1 2
timestamp 1674174324
<< viali >>
rect 8327 37417 8361 37451
rect 16313 37417 16347 37451
rect 17693 37417 17727 37451
rect 38025 37349 38059 37383
rect 3157 37281 3191 37315
rect 3985 37281 4019 37315
rect 5733 37281 5767 37315
rect 10609 37281 10643 37315
rect 11713 37281 11747 37315
rect 14289 37281 14323 37315
rect 15577 37281 15611 37315
rect 18153 37281 18187 37315
rect 34345 37281 34379 37315
rect 3433 37213 3467 37247
rect 6009 37213 6043 37247
rect 8585 37213 8619 37247
rect 10885 37213 10919 37247
rect 11989 37213 12023 37247
rect 13277 37213 13311 37247
rect 15117 37213 15151 37247
rect 17049 37213 17083 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22017 37213 22051 37247
rect 24593 37213 24627 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 29745 37213 29779 37247
rect 31217 37213 31251 37247
rect 31677 37213 31711 37247
rect 32597 37213 32631 37247
rect 34897 37213 34931 37247
rect 36461 37213 36495 37247
rect 37565 37213 37599 37247
rect 38209 37213 38243 37247
rect 6561 37145 6595 37179
rect 1685 37077 1719 37111
rect 9137 37077 9171 37111
rect 13093 37077 13127 37111
rect 14933 37077 14967 37111
rect 16957 37077 16991 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 24777 37077 24811 37111
rect 25513 37077 25547 37111
rect 27353 37077 27387 37111
rect 29929 37077 29963 37111
rect 31033 37077 31067 37111
rect 32413 37077 32447 37111
rect 35081 37077 35115 37111
rect 36277 37077 36311 37111
rect 14749 36873 14783 36907
rect 17049 36873 17083 36907
rect 32505 36873 32539 36907
rect 38209 36873 38243 36907
rect 5825 36805 5859 36839
rect 10517 36805 10551 36839
rect 11989 36805 12023 36839
rect 1593 36737 1627 36771
rect 4905 36737 4939 36771
rect 10793 36737 10827 36771
rect 11713 36737 11747 36771
rect 14289 36737 14323 36771
rect 16865 36737 16899 36771
rect 28181 36737 28215 36771
rect 32321 36737 32355 36771
rect 37565 36737 37599 36771
rect 38025 36737 38059 36771
rect 1869 36669 1903 36703
rect 2881 36669 2915 36703
rect 4629 36669 4663 36703
rect 6561 36669 6595 36703
rect 8309 36669 8343 36703
rect 8585 36669 8619 36703
rect 9045 36669 9079 36703
rect 13461 36669 13495 36703
rect 27905 36669 27939 36703
rect 6009 36601 6043 36635
rect 31769 36601 31803 36635
rect 14105 36533 14139 36567
rect 15301 36533 15335 36567
rect 15853 36533 15887 36567
rect 25237 36533 25271 36567
rect 4077 36329 4111 36363
rect 16497 36329 16531 36363
rect 12081 36261 12115 36295
rect 13185 36261 13219 36295
rect 1685 36193 1719 36227
rect 10885 36193 10919 36227
rect 11529 36193 11563 36227
rect 12633 36193 12667 36227
rect 14841 36193 14875 36227
rect 15393 36193 15427 36227
rect 4261 36125 4295 36159
rect 6837 36125 6871 36159
rect 7297 36125 7331 36159
rect 8033 36125 8067 36159
rect 1961 36057 1995 36091
rect 4813 36057 4847 36091
rect 6561 36057 6595 36091
rect 8585 36057 8619 36091
rect 10609 36057 10643 36091
rect 15945 36057 15979 36091
rect 37565 36057 37599 36091
rect 38209 36057 38243 36091
rect 3433 35989 3467 36023
rect 7849 35989 7883 36023
rect 9137 35989 9171 36023
rect 14289 35989 14323 36023
rect 38117 35989 38151 36023
rect 11069 35785 11103 35819
rect 15669 35785 15703 35819
rect 23305 35785 23339 35819
rect 38209 35785 38243 35819
rect 1961 35717 1995 35751
rect 4537 35717 4571 35751
rect 4721 35717 4755 35751
rect 14473 35717 14507 35751
rect 3985 35649 4019 35683
rect 5365 35649 5399 35683
rect 10057 35649 10091 35683
rect 12265 35649 12299 35683
rect 12357 35647 12391 35681
rect 23121 35649 23155 35683
rect 23765 35649 23799 35683
rect 38025 35649 38059 35683
rect 3709 35581 3743 35615
rect 6561 35581 6595 35615
rect 7297 35581 7331 35615
rect 8769 35581 8803 35615
rect 9045 35581 9079 35615
rect 10517 35581 10551 35615
rect 15025 35581 15059 35615
rect 9873 35513 9907 35547
rect 13921 35513 13955 35547
rect 5181 35445 5215 35479
rect 5917 35445 5951 35479
rect 12909 35445 12943 35479
rect 13461 35445 13495 35479
rect 4077 35241 4111 35275
rect 13185 35241 13219 35275
rect 13737 35241 13771 35275
rect 14381 35241 14415 35275
rect 3433 35105 3467 35139
rect 5181 35105 5215 35139
rect 7205 35105 7239 35139
rect 7941 35105 7975 35139
rect 8493 35105 8527 35139
rect 9137 35105 9171 35139
rect 4261 35037 4295 35071
rect 11805 35037 11839 35071
rect 12449 35037 12483 35071
rect 3157 34969 3191 35003
rect 6929 34969 6963 35003
rect 9413 34969 9447 35003
rect 11897 34969 11931 35003
rect 1685 34901 1719 34935
rect 10885 34901 10919 34935
rect 12541 34901 12575 34935
rect 5089 34697 5123 34731
rect 11069 34697 11103 34731
rect 13093 34697 13127 34731
rect 2237 34629 2271 34663
rect 11989 34629 12023 34663
rect 14105 34629 14139 34663
rect 4629 34561 4663 34595
rect 6561 34561 6595 34595
rect 10609 34561 10643 34595
rect 1961 34493 1995 34527
rect 3985 34493 4019 34527
rect 6009 34493 6043 34527
rect 11897 34493 11931 34527
rect 12357 34493 12391 34527
rect 13645 34493 13679 34527
rect 38025 34493 38059 34527
rect 38301 34493 38335 34527
rect 8309 34425 8343 34459
rect 4445 34357 4479 34391
rect 6824 34357 6858 34391
rect 8861 34357 8895 34391
rect 10345 34357 10379 34391
rect 8033 34153 8067 34187
rect 8493 34153 8527 34187
rect 10885 34153 10919 34187
rect 7481 34085 7515 34119
rect 38301 34085 38335 34119
rect 1685 34017 1719 34051
rect 1961 34017 1995 34051
rect 4905 34017 4939 34051
rect 5181 34017 5215 34051
rect 9137 34017 9171 34051
rect 11713 34017 11747 34051
rect 4445 33949 4479 33983
rect 6929 33949 6963 33983
rect 12817 33949 12851 33983
rect 13553 33949 13587 33983
rect 14933 33949 14967 33983
rect 4169 33881 4203 33915
rect 9413 33881 9447 33915
rect 11805 33881 11839 33915
rect 12357 33881 12391 33915
rect 12909 33881 12943 33915
rect 3433 33813 3467 33847
rect 13645 33813 13679 33847
rect 14289 33813 14323 33847
rect 15025 33813 15059 33847
rect 11805 33609 11839 33643
rect 1961 33541 1995 33575
rect 3709 33541 3743 33575
rect 8125 33541 8159 33575
rect 14197 33541 14231 33575
rect 14749 33541 14783 33575
rect 3985 33473 4019 33507
rect 4905 33473 4939 33507
rect 5825 33473 5859 33507
rect 8401 33473 8435 33507
rect 8861 33473 8895 33507
rect 11713 33473 11747 33507
rect 12449 33473 12483 33507
rect 4721 33405 4755 33439
rect 5641 33405 5675 33439
rect 9137 33405 9171 33439
rect 11069 33405 11103 33439
rect 14105 33405 14139 33439
rect 6653 33269 6687 33303
rect 10609 33269 10643 33303
rect 4077 33065 4111 33099
rect 9137 33065 9171 33099
rect 9689 33065 9723 33099
rect 10885 33065 10919 33099
rect 11437 33065 11471 33099
rect 3157 32929 3191 32963
rect 3433 32929 3467 32963
rect 4813 32929 4847 32963
rect 4261 32861 4295 32895
rect 6837 32861 6871 32895
rect 7297 32861 7331 32895
rect 7849 32861 7883 32895
rect 11345 32861 11379 32895
rect 6561 32793 6595 32827
rect 8401 32793 8435 32827
rect 38025 32793 38059 32827
rect 38209 32793 38243 32827
rect 1685 32725 1719 32759
rect 10241 32725 10275 32759
rect 37565 32725 37599 32759
rect 7113 32521 7147 32555
rect 15025 32453 15059 32487
rect 15945 32453 15979 32487
rect 1593 32385 1627 32419
rect 4997 32385 5031 32419
rect 5641 32385 5675 32419
rect 8861 32385 8895 32419
rect 9321 32385 9355 32419
rect 9873 32385 9907 32419
rect 10425 32385 10459 32419
rect 12541 32385 12575 32419
rect 13185 32385 13219 32419
rect 1869 32317 1903 32351
rect 2973 32317 3007 32351
rect 4721 32317 4755 32351
rect 8585 32317 8619 32351
rect 14933 32317 14967 32351
rect 12633 32249 12667 32283
rect 5549 32181 5583 32215
rect 13277 32181 13311 32215
rect 6377 31977 6411 32011
rect 9137 31977 9171 32011
rect 9689 31977 9723 32011
rect 1961 31841 1995 31875
rect 3433 31841 3467 31875
rect 4629 31841 4663 31875
rect 7113 31841 7147 31875
rect 8585 31841 8619 31875
rect 1685 31773 1719 31807
rect 3985 31773 4019 31807
rect 6837 31773 6871 31807
rect 18521 31773 18555 31807
rect 18613 31773 18647 31807
rect 19441 31773 19475 31807
rect 4905 31705 4939 31739
rect 4077 31637 4111 31671
rect 6561 31433 6595 31467
rect 8033 31365 8067 31399
rect 16129 31365 16163 31399
rect 1777 31297 1811 31331
rect 3985 31297 4019 31331
rect 8769 31297 8803 31331
rect 14749 31297 14783 31331
rect 20453 31297 20487 31331
rect 21097 31297 21131 31331
rect 2053 31229 2087 31263
rect 4261 31229 4295 31263
rect 8309 31229 8343 31263
rect 9413 31229 9447 31263
rect 9965 31229 9999 31263
rect 15393 31229 15427 31263
rect 16221 31229 16255 31263
rect 14105 31161 14139 31195
rect 20637 31161 20671 31195
rect 3525 31093 3559 31127
rect 5733 31093 5767 31127
rect 8861 31093 8895 31127
rect 14657 31093 14691 31127
rect 1869 30889 1903 30923
rect 2513 30889 2547 30923
rect 3157 30889 3191 30923
rect 4721 30889 4755 30923
rect 6180 30889 6214 30923
rect 16313 30889 16347 30923
rect 16865 30889 16899 30923
rect 37565 30889 37599 30923
rect 5365 30821 5399 30855
rect 7665 30821 7699 30855
rect 5917 30753 5951 30787
rect 11621 30753 11655 30787
rect 12265 30753 12299 30787
rect 12541 30753 12575 30787
rect 14565 30753 14599 30787
rect 1961 30685 1995 30719
rect 2421 30685 2455 30719
rect 3249 30685 3283 30719
rect 3985 30685 4019 30719
rect 4621 30695 4655 30729
rect 5273 30685 5307 30719
rect 8125 30685 8159 30719
rect 9137 30685 9171 30719
rect 11529 30685 11563 30719
rect 15853 30685 15887 30719
rect 37381 30685 37415 30719
rect 38025 30685 38059 30719
rect 4077 30617 4111 30651
rect 11069 30617 11103 30651
rect 12357 30617 12391 30651
rect 14657 30617 14691 30651
rect 15209 30617 15243 30651
rect 8217 30549 8251 30583
rect 9229 30549 9263 30583
rect 15761 30549 15795 30583
rect 38209 30549 38243 30583
rect 12357 30345 12391 30379
rect 2421 30277 2455 30311
rect 4077 30277 4111 30311
rect 5457 30277 5491 30311
rect 6653 30277 6687 30311
rect 7205 30277 7239 30311
rect 7757 30277 7791 30311
rect 14749 30277 14783 30311
rect 14841 30277 14875 30311
rect 16129 30277 16163 30311
rect 1869 30209 1903 30243
rect 2329 30209 2363 30243
rect 2973 30209 3007 30243
rect 4169 30209 4203 30243
rect 4721 30209 4755 30243
rect 5365 30209 5399 30243
rect 6561 30209 6595 30243
rect 10149 30209 10183 30243
rect 12449 30209 12483 30243
rect 1777 30141 1811 30175
rect 3065 30141 3099 30175
rect 13737 30141 13771 30175
rect 15577 30141 15611 30175
rect 16221 30141 16255 30175
rect 4813 30073 4847 30107
rect 14289 30073 14323 30107
rect 10241 30005 10275 30039
rect 16865 30005 16899 30039
rect 17969 30005 18003 30039
rect 18429 30005 18463 30039
rect 3341 29801 3375 29835
rect 4905 29801 4939 29835
rect 6561 29801 6595 29835
rect 7113 29801 7147 29835
rect 12541 29801 12575 29835
rect 14657 29801 14691 29835
rect 4261 29733 4295 29767
rect 2697 29665 2731 29699
rect 5917 29665 5951 29699
rect 15301 29665 15335 29699
rect 1869 29597 1903 29631
rect 2605 29597 2639 29631
rect 3433 29597 3467 29631
rect 4169 29597 4203 29631
rect 4813 29597 4847 29631
rect 6009 29597 6043 29631
rect 13553 29597 13587 29631
rect 14565 29597 14599 29631
rect 17049 29597 17083 29631
rect 18061 29597 18095 29631
rect 18705 29597 18739 29631
rect 30113 29597 30147 29631
rect 15393 29529 15427 29563
rect 16313 29529 16347 29563
rect 1685 29461 1719 29495
rect 13093 29461 13127 29495
rect 13645 29461 13679 29495
rect 17141 29461 17175 29495
rect 18153 29461 18187 29495
rect 30021 29461 30055 29495
rect 2237 29257 2271 29291
rect 4169 29257 4203 29291
rect 5917 29257 5951 29291
rect 6653 29257 6687 29291
rect 7297 29257 7331 29291
rect 13553 29257 13587 29291
rect 20361 29257 20395 29291
rect 8309 29189 8343 29223
rect 12081 29189 12115 29223
rect 14289 29189 14323 29223
rect 15485 29189 15519 29223
rect 16865 29189 16899 29223
rect 17417 29189 17451 29223
rect 18061 29189 18095 29223
rect 18613 29189 18647 29223
rect 2145 29121 2179 29155
rect 2789 29121 2823 29155
rect 3433 29121 3467 29155
rect 4261 29121 4295 29155
rect 4721 29121 4755 29155
rect 5825 29121 5859 29155
rect 6745 29121 6779 29155
rect 10333 29121 10367 29155
rect 13461 29121 13495 29155
rect 19809 29121 19843 29155
rect 37565 29121 37599 29155
rect 38209 29121 38243 29155
rect 3525 29053 3559 29087
rect 8217 29053 8251 29087
rect 8861 29053 8895 29087
rect 11989 29053 12023 29087
rect 12633 29053 12667 29087
rect 14197 29053 14231 29087
rect 15393 29053 15427 29087
rect 16037 29053 16071 29087
rect 17509 29053 17543 29087
rect 18705 29053 18739 29087
rect 19717 29053 19751 29087
rect 1685 28985 1719 29019
rect 10425 28985 10459 29019
rect 14749 28985 14783 29019
rect 38025 28985 38059 29019
rect 2881 28917 2915 28951
rect 4813 28917 4847 28951
rect 1685 28713 1719 28747
rect 2881 28713 2915 28747
rect 6561 28713 6595 28747
rect 7205 28713 7239 28747
rect 7757 28713 7791 28747
rect 11345 28713 11379 28747
rect 11989 28713 12023 28747
rect 13645 28713 13679 28747
rect 2237 28645 2271 28679
rect 4077 28645 4111 28679
rect 5917 28645 5951 28679
rect 4813 28577 4847 28611
rect 9781 28577 9815 28611
rect 14381 28577 14415 28611
rect 15393 28577 15427 28611
rect 16589 28577 16623 28611
rect 17601 28577 17635 28611
rect 2145 28509 2179 28543
rect 2789 28509 2823 28543
rect 4169 28509 4203 28543
rect 4721 28509 4755 28543
rect 5825 28509 5859 28543
rect 6469 28509 6503 28543
rect 7113 28509 7147 28543
rect 10517 28509 10551 28543
rect 11897 28509 11931 28543
rect 12909 28509 12943 28543
rect 13553 28509 13587 28543
rect 16037 28509 16071 28543
rect 18245 28509 18279 28543
rect 18705 28509 18739 28543
rect 20085 28509 20119 28543
rect 20637 28509 20671 28543
rect 37841 28509 37875 28543
rect 9137 28441 9171 28475
rect 9689 28441 9723 28475
rect 10609 28441 10643 28475
rect 14473 28441 14507 28475
rect 16681 28441 16715 28475
rect 13001 28373 13035 28407
rect 15945 28373 15979 28407
rect 18153 28373 18187 28407
rect 18797 28373 18831 28407
rect 19993 28373 20027 28407
rect 38025 28373 38059 28407
rect 3525 28169 3559 28203
rect 4169 28169 4203 28203
rect 6009 28169 6043 28203
rect 6837 28169 6871 28203
rect 11805 28169 11839 28203
rect 2881 28101 2915 28135
rect 14565 28101 14599 28135
rect 15761 28101 15795 28135
rect 18061 28101 18095 28135
rect 1869 28033 1903 28067
rect 2789 28033 2823 28067
rect 3617 28033 3651 28067
rect 10149 28033 10183 28067
rect 10793 28033 10827 28067
rect 11713 28033 11747 28067
rect 12449 28033 12483 28067
rect 13093 28033 13127 28067
rect 13737 28033 13771 28067
rect 16313 28033 16347 28067
rect 23673 28033 23707 28067
rect 24317 28033 24351 28067
rect 13185 27965 13219 27999
rect 14473 27965 14507 27999
rect 15669 27965 15703 27999
rect 17877 27965 17911 27999
rect 18153 27965 18187 27999
rect 18705 27965 18739 27999
rect 19349 27965 19383 27999
rect 1685 27897 1719 27931
rect 12541 27897 12575 27931
rect 15025 27897 15059 27931
rect 20085 27897 20119 27931
rect 23857 27897 23891 27931
rect 10057 27829 10091 27863
rect 10885 27829 10919 27863
rect 13829 27829 13863 27863
rect 20545 27829 20579 27863
rect 1593 27557 1627 27591
rect 21189 27557 21223 27591
rect 9781 27489 9815 27523
rect 11161 27489 11195 27523
rect 13369 27489 13403 27523
rect 15669 27489 15703 27523
rect 15945 27489 15979 27523
rect 16865 27489 16899 27523
rect 17141 27489 17175 27523
rect 17969 27489 18003 27523
rect 18337 27489 18371 27523
rect 11989 27421 12023 27455
rect 14657 27421 14691 27455
rect 19625 27421 19659 27455
rect 20637 27421 20671 27455
rect 9137 27353 9171 27387
rect 9689 27353 9723 27387
rect 10885 27353 10919 27387
rect 10977 27353 11011 27387
rect 13093 27353 13127 27387
rect 13185 27353 13219 27387
rect 15853 27353 15887 27387
rect 17049 27353 17083 27387
rect 18245 27353 18279 27387
rect 20085 27353 20119 27387
rect 12081 27285 12115 27319
rect 14749 27285 14783 27319
rect 19533 27285 19567 27319
rect 9413 27081 9447 27115
rect 12817 27081 12851 27115
rect 14013 27013 14047 27047
rect 14565 27013 14599 27047
rect 14657 27013 14691 27047
rect 15761 27013 15795 27047
rect 15853 27013 15887 27047
rect 18429 27013 18463 27047
rect 18521 27013 18555 27047
rect 20361 27013 20395 27047
rect 8953 26945 8987 26979
rect 12081 26945 12115 26979
rect 12725 26945 12759 26979
rect 13553 26945 13587 26979
rect 17325 26945 17359 26979
rect 19257 26945 19291 26979
rect 19901 26945 19935 26979
rect 38025 26945 38059 26979
rect 10057 26877 10091 26911
rect 10609 26877 10643 26911
rect 15209 26877 15243 26911
rect 18153 26877 18187 26911
rect 11161 26809 11195 26843
rect 12173 26809 12207 26843
rect 19809 26809 19843 26843
rect 13369 26741 13403 26775
rect 17233 26741 17267 26775
rect 19165 26741 19199 26775
rect 20913 26741 20947 26775
rect 38209 26741 38243 26775
rect 12081 26401 12115 26435
rect 12909 26401 12943 26435
rect 15393 26401 15427 26435
rect 15853 26401 15887 26435
rect 17601 26401 17635 26435
rect 18797 26401 18831 26435
rect 19441 26401 19475 26435
rect 1869 26333 1903 26367
rect 9873 26333 9907 26367
rect 10701 26333 10735 26367
rect 10793 26333 10827 26367
rect 20269 26333 20303 26367
rect 20361 26333 20395 26367
rect 20821 26333 20855 26367
rect 29193 26333 29227 26367
rect 8493 26265 8527 26299
rect 9965 26265 9999 26299
rect 11437 26265 11471 26299
rect 11529 26265 11563 26299
rect 12633 26265 12667 26299
rect 12725 26265 12759 26299
rect 14841 26265 14875 26299
rect 15485 26265 15519 26299
rect 16957 26265 16991 26299
rect 17509 26265 17543 26299
rect 18153 26265 18187 26299
rect 18705 26265 18739 26299
rect 19625 26265 19659 26299
rect 21373 26265 21407 26299
rect 29101 26265 29135 26299
rect 1685 26197 1719 26231
rect 9413 26197 9447 26231
rect 11069 25993 11103 26027
rect 20177 25993 20211 26027
rect 20913 25993 20947 26027
rect 12633 25925 12667 25959
rect 13277 25925 13311 25959
rect 15301 25925 15335 25959
rect 15853 25925 15887 25959
rect 17601 25925 17635 25959
rect 18245 25925 18279 25959
rect 18797 25925 18831 25959
rect 9321 25857 9355 25891
rect 10333 25857 10367 25891
rect 10977 25857 11011 25891
rect 12541 25857 12575 25891
rect 14657 25857 14691 25891
rect 17049 25857 17083 25891
rect 19625 25857 19659 25891
rect 20269 25857 20303 25891
rect 20729 25857 20763 25891
rect 11897 25789 11931 25823
rect 13185 25789 13219 25823
rect 13461 25789 13495 25823
rect 14749 25789 14783 25823
rect 15945 25789 15979 25823
rect 17693 25789 17727 25823
rect 18889 25789 18923 25823
rect 10425 25721 10459 25755
rect 9781 25653 9815 25687
rect 19533 25653 19567 25687
rect 21465 25653 21499 25687
rect 10793 25449 10827 25483
rect 19533 25449 19567 25483
rect 20637 25449 20671 25483
rect 21649 25449 21683 25483
rect 28641 25449 28675 25483
rect 36277 25449 36311 25483
rect 11989 25381 12023 25415
rect 13185 25381 13219 25415
rect 7941 25313 7975 25347
rect 9597 25313 9631 25347
rect 12633 25313 12667 25347
rect 16129 25313 16163 25347
rect 18153 25313 18187 25347
rect 38025 25313 38059 25347
rect 10057 25245 10091 25279
rect 10701 25245 10735 25279
rect 14473 25245 14507 25279
rect 15117 25245 15151 25279
rect 17509 25245 17543 25279
rect 19625 25245 19659 25279
rect 20177 25245 20211 25279
rect 21741 25245 21775 25279
rect 22293 25245 22327 25279
rect 28457 25245 28491 25279
rect 36829 25245 36863 25279
rect 38301 25245 38335 25279
rect 7297 25177 7331 25211
rect 7389 25177 7423 25211
rect 10149 25177 10183 25211
rect 11437 25177 11471 25211
rect 11529 25177 11563 25211
rect 12725 25177 12759 25211
rect 15853 25177 15887 25211
rect 15945 25177 15979 25211
rect 18705 25177 18739 25211
rect 18797 25177 18831 25211
rect 29193 25177 29227 25211
rect 14565 25109 14599 25143
rect 15209 25109 15243 25143
rect 17601 25109 17635 25143
rect 36921 25109 36955 25143
rect 7573 24905 7607 24939
rect 38301 24905 38335 24939
rect 9873 24837 9907 24871
rect 11713 24837 11747 24871
rect 13185 24837 13219 24871
rect 14657 24837 14691 24871
rect 17417 24837 17451 24871
rect 18153 24837 18187 24871
rect 18705 24837 18739 24871
rect 20085 24837 20119 24871
rect 1869 24769 1903 24803
rect 2513 24769 2547 24803
rect 7665 24769 7699 24803
rect 10517 24769 10551 24803
rect 10977 24769 11011 24803
rect 11989 24769 12023 24803
rect 13829 24769 13863 24803
rect 16129 24769 16163 24803
rect 16221 24769 16255 24803
rect 19625 24769 19659 24803
rect 20177 24769 20211 24803
rect 20821 24769 20855 24803
rect 11069 24701 11103 24735
rect 12817 24701 12851 24735
rect 13277 24701 13311 24735
rect 14565 24701 14599 24735
rect 15577 24701 15611 24735
rect 17509 24701 17543 24735
rect 18797 24701 18831 24735
rect 19349 24701 19383 24735
rect 2053 24633 2087 24667
rect 10425 24633 10459 24667
rect 13921 24633 13955 24667
rect 16957 24633 16991 24667
rect 5089 24361 5123 24395
rect 14657 24361 14691 24395
rect 18889 24361 18923 24395
rect 26893 24361 26927 24395
rect 19441 24293 19475 24327
rect 12449 24225 12483 24259
rect 13737 24225 13771 24259
rect 15945 24225 15979 24259
rect 16589 24225 16623 24259
rect 17785 24225 17819 24259
rect 1869 24157 1903 24191
rect 4997 24157 5031 24191
rect 5641 24157 5675 24191
rect 10609 24157 10643 24191
rect 12357 24157 12391 24191
rect 14289 24157 14323 24191
rect 14473 24157 14507 24191
rect 17049 24157 17083 24191
rect 19625 24157 19659 24191
rect 26709 24157 26743 24191
rect 10701 24089 10735 24123
rect 13093 24089 13127 24123
rect 13185 24089 13219 24123
rect 16014 24089 16048 24123
rect 18153 24089 18187 24123
rect 18245 24089 18279 24123
rect 1685 24021 1719 24055
rect 11345 24021 11379 24055
rect 11897 24021 11931 24055
rect 20085 24021 20119 24055
rect 27445 24021 27479 24055
rect 11805 23817 11839 23851
rect 12817 23817 12851 23851
rect 14197 23817 14231 23851
rect 14841 23817 14875 23851
rect 19349 23817 19383 23851
rect 15577 23749 15611 23783
rect 16129 23749 16163 23783
rect 17049 23749 17083 23783
rect 18153 23749 18187 23783
rect 18245 23749 18279 23783
rect 12265 23681 12299 23715
rect 13369 23681 13403 23715
rect 14197 23681 14231 23715
rect 14749 23681 14783 23715
rect 19533 23681 19567 23715
rect 38025 23681 38059 23715
rect 15485 23613 15519 23647
rect 16957 23613 16991 23647
rect 18429 23613 18463 23647
rect 13461 23545 13495 23579
rect 17509 23545 17543 23579
rect 20085 23477 20119 23511
rect 38209 23477 38243 23511
rect 1961 23273 1995 23307
rect 13553 23273 13587 23307
rect 14841 23273 14875 23307
rect 17601 23205 17635 23239
rect 13001 23137 13035 23171
rect 14381 23137 14415 23171
rect 15301 23137 15335 23171
rect 15485 23137 15519 23171
rect 2145 23069 2179 23103
rect 12449 23069 12483 23103
rect 13645 23069 13679 23103
rect 19901 23069 19935 23103
rect 20085 23069 20119 23103
rect 16037 23001 16071 23035
rect 16129 23001 16163 23035
rect 17049 23001 17083 23035
rect 18061 23001 18095 23035
rect 18153 23001 18187 23035
rect 2697 22933 2731 22967
rect 18705 22933 18739 22967
rect 19441 22933 19475 22967
rect 13185 22729 13219 22763
rect 13737 22729 13771 22763
rect 16129 22729 16163 22763
rect 17233 22729 17267 22763
rect 23397 22729 23431 22763
rect 24041 22729 24075 22763
rect 14933 22661 14967 22695
rect 15025 22661 15059 22695
rect 17969 22661 18003 22695
rect 14197 22593 14231 22627
rect 16221 22593 16255 22627
rect 17141 22593 17175 22627
rect 23489 22593 23523 22627
rect 15209 22525 15243 22559
rect 17877 22525 17911 22559
rect 18889 22525 18923 22559
rect 14289 22389 14323 22423
rect 15025 22185 15059 22219
rect 18153 22185 18187 22219
rect 14841 22049 14875 22083
rect 16589 22049 16623 22083
rect 1869 21981 1903 22015
rect 14657 21981 14691 22015
rect 18245 21981 18279 22015
rect 37933 21981 37967 22015
rect 15853 21913 15887 21947
rect 16681 21913 16715 21947
rect 17601 21913 17635 21947
rect 1685 21845 1719 21879
rect 13737 21845 13771 21879
rect 15945 21845 15979 21879
rect 18705 21845 18739 21879
rect 37749 21845 37783 21879
rect 14197 21641 14231 21675
rect 14657 21641 14691 21675
rect 15393 21641 15427 21675
rect 18061 21641 18095 21675
rect 13645 21505 13679 21539
rect 14841 21505 14875 21539
rect 15485 21505 15519 21539
rect 18705 21505 18739 21539
rect 19165 21505 19199 21539
rect 38025 21505 38059 21539
rect 16313 21437 16347 21471
rect 17417 21437 17451 21471
rect 17601 21437 17635 21471
rect 16957 21369 16991 21403
rect 18613 21301 18647 21335
rect 38209 21301 38243 21335
rect 14289 21097 14323 21131
rect 14933 21097 14967 21131
rect 16957 21097 16991 21131
rect 17785 21097 17819 21131
rect 16589 20961 16623 20995
rect 16773 20961 16807 20995
rect 15025 20893 15059 20927
rect 16129 20893 16163 20927
rect 17877 20893 17911 20927
rect 18337 20893 18371 20927
rect 1685 20825 1719 20859
rect 1777 20757 1811 20791
rect 16037 20757 16071 20791
rect 15209 20553 15243 20587
rect 16313 20553 16347 20587
rect 17601 20553 17635 20587
rect 30113 20553 30147 20587
rect 38025 20553 38059 20587
rect 1593 20485 1627 20519
rect 15853 20417 15887 20451
rect 17049 20417 17083 20451
rect 17693 20417 17727 20451
rect 30205 20417 30239 20451
rect 37841 20417 37875 20451
rect 15669 20349 15703 20383
rect 14565 20213 14599 20247
rect 16957 20213 16991 20247
rect 18245 20213 18279 20247
rect 15669 20009 15703 20043
rect 16957 20009 16991 20043
rect 17601 20009 17635 20043
rect 16589 19873 16623 19907
rect 15761 19805 15795 19839
rect 16405 19805 16439 19839
rect 17693 19805 17727 19839
rect 15117 19669 15151 19703
rect 18153 19669 18187 19703
rect 15301 19465 15335 19499
rect 17969 19465 18003 19499
rect 15209 19329 15243 19363
rect 15945 19329 15979 19363
rect 17141 19329 17175 19363
rect 17233 19329 17267 19363
rect 18613 19329 18647 19363
rect 37565 19329 37599 19363
rect 38209 19329 38243 19363
rect 18429 19261 18463 19295
rect 38025 19261 38059 19295
rect 16129 19193 16163 19227
rect 17049 18921 17083 18955
rect 6193 18717 6227 18751
rect 1685 18649 1719 18683
rect 1869 18649 1903 18683
rect 6101 18581 6135 18615
rect 1593 18377 1627 18411
rect 19717 17833 19751 17867
rect 19809 17629 19843 17663
rect 20361 17493 20395 17527
rect 20361 17153 20395 17187
rect 20269 16949 20303 16983
rect 21005 16949 21039 16983
rect 1869 16541 1903 16575
rect 14657 16541 14691 16575
rect 1685 16405 1719 16439
rect 14473 16405 14507 16439
rect 15117 16405 15151 16439
rect 10609 16133 10643 16167
rect 9873 16065 9907 16099
rect 12173 16065 12207 16099
rect 12633 16065 12667 16099
rect 19809 16065 19843 16099
rect 20453 16065 20487 16099
rect 37473 16065 37507 16099
rect 38025 16065 38059 16099
rect 11989 15929 12023 15963
rect 9689 15861 9723 15895
rect 10517 15861 10551 15895
rect 19993 15861 20027 15895
rect 38209 15861 38243 15895
rect 9965 15657 9999 15691
rect 10885 15657 10919 15691
rect 16129 15657 16163 15691
rect 16221 15453 16255 15487
rect 16681 15317 16715 15351
rect 1685 14297 1719 14331
rect 1777 14229 1811 14263
rect 1685 14025 1719 14059
rect 38025 13889 38059 13923
rect 38301 13821 38335 13855
rect 38301 13481 38335 13515
rect 1869 13277 1903 13311
rect 1685 13141 1719 13175
rect 37565 11713 37599 11747
rect 38209 11713 38243 11747
rect 38025 11577 38059 11611
rect 16497 11305 16531 11339
rect 2421 11169 2455 11203
rect 1869 11101 1903 11135
rect 16589 11101 16623 11135
rect 17141 11033 17175 11067
rect 1685 10965 1719 10999
rect 15025 10761 15059 10795
rect 17233 10761 17267 10795
rect 18797 10761 18831 10795
rect 15117 10625 15151 10659
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 37565 10625 37599 10659
rect 38209 10625 38243 10659
rect 38025 10489 38059 10523
rect 15669 10421 15703 10455
rect 18337 10421 18371 10455
rect 15117 10217 15151 10251
rect 14565 10013 14599 10047
rect 14381 9877 14415 9911
rect 17417 9877 17451 9911
rect 16957 9605 16991 9639
rect 17049 9537 17083 9571
rect 17509 9333 17543 9367
rect 1869 8925 1903 8959
rect 24593 8925 24627 8959
rect 25237 8925 25271 8959
rect 1685 8789 1719 8823
rect 24777 8789 24811 8823
rect 38117 8585 38151 8619
rect 37657 8449 37691 8483
rect 38301 8449 38335 8483
rect 23213 7973 23247 8007
rect 23029 7769 23063 7803
rect 1685 7361 1719 7395
rect 1777 7157 1811 7191
rect 1593 6953 1627 6987
rect 38025 6341 38059 6375
rect 37565 6273 37599 6307
rect 38209 6273 38243 6307
rect 1869 5661 1903 5695
rect 2329 5661 2363 5695
rect 1685 5525 1719 5559
rect 38025 4709 38059 4743
rect 37565 4505 37599 4539
rect 38209 4505 38243 4539
rect 2329 3689 2363 3723
rect 1869 3485 1903 3519
rect 38025 3417 38059 3451
rect 38209 3417 38243 3451
rect 1685 3349 1719 3383
rect 37565 3349 37599 3383
rect 5733 3145 5767 3179
rect 37473 3145 37507 3179
rect 1869 3009 1903 3043
rect 13001 3009 13035 3043
rect 14565 3009 14599 3043
rect 15761 3009 15795 3043
rect 16221 3009 16255 3043
rect 17417 3009 17451 3043
rect 19165 3009 19199 3043
rect 19809 3009 19843 3043
rect 23765 3009 23799 3043
rect 24869 3009 24903 3043
rect 25513 3009 25547 3043
rect 27169 3009 27203 3043
rect 27813 3009 27847 3043
rect 38025 3009 38059 3043
rect 13829 2941 13863 2975
rect 14289 2941 14323 2975
rect 12817 2873 12851 2907
rect 15577 2873 15611 2907
rect 18153 2873 18187 2907
rect 27353 2873 27387 2907
rect 36921 2873 36955 2907
rect 1685 2805 1719 2839
rect 2789 2805 2823 2839
rect 17601 2805 17635 2839
rect 19257 2805 19291 2839
rect 23581 2805 23615 2839
rect 24961 2805 24995 2839
rect 29653 2805 29687 2839
rect 38209 2805 38243 2839
rect 10609 2601 10643 2635
rect 13185 2601 13219 2635
rect 28549 2601 28583 2635
rect 29837 2601 29871 2635
rect 32413 2601 32447 2635
rect 33701 2601 33735 2635
rect 36737 2601 36771 2635
rect 2421 2533 2455 2567
rect 38025 2533 38059 2567
rect 4261 2465 4295 2499
rect 9413 2465 9447 2499
rect 16313 2465 16347 2499
rect 16865 2465 16899 2499
rect 24869 2465 24903 2499
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 5549 2397 5583 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 11069 2397 11103 2431
rect 12633 2397 12667 2431
rect 16037 2397 16071 2431
rect 17509 2397 17543 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 22753 2397 22787 2431
rect 24041 2397 24075 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 35541 2397 35575 2431
rect 36921 2397 36955 2431
rect 37473 2397 37507 2431
rect 27997 2329 28031 2363
rect 28641 2329 28675 2363
rect 29929 2329 29963 2363
rect 32505 2329 32539 2363
rect 33149 2329 33183 2363
rect 33793 2329 33827 2363
rect 38209 2329 38243 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 5365 2261 5399 2295
rect 7297 2261 7331 2295
rect 8493 2261 8527 2295
rect 12449 2261 12483 2295
rect 17693 2261 17727 2295
rect 19625 2261 19659 2295
rect 22201 2261 22235 2295
rect 22937 2261 22971 2295
rect 27353 2261 27387 2295
rect 31769 2261 31803 2295
rect 35725 2261 35759 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 7282 37448 7288 37460
rect 3896 37420 7288 37448
rect 3145 37315 3203 37321
rect 3145 37281 3157 37315
rect 3191 37312 3203 37315
rect 3896 37312 3924 37420
rect 7282 37408 7288 37420
rect 7340 37408 7346 37460
rect 8315 37451 8373 37457
rect 8315 37417 8327 37451
rect 8361 37448 8373 37451
rect 10134 37448 10140 37460
rect 8361 37420 10140 37448
rect 8361 37417 8373 37420
rect 8315 37411 8373 37417
rect 10134 37408 10140 37420
rect 10192 37448 10198 37460
rect 10870 37448 10876 37460
rect 10192 37420 10876 37448
rect 10192 37408 10198 37420
rect 10870 37408 10876 37420
rect 10928 37408 10934 37460
rect 16301 37451 16359 37457
rect 16301 37417 16313 37451
rect 16347 37448 16359 37451
rect 16758 37448 16764 37460
rect 16347 37420 16764 37448
rect 16347 37417 16359 37420
rect 16301 37411 16359 37417
rect 16758 37408 16764 37420
rect 16816 37408 16822 37460
rect 17681 37451 17739 37457
rect 17681 37417 17693 37451
rect 17727 37448 17739 37451
rect 18046 37448 18052 37460
rect 17727 37420 18052 37448
rect 17727 37417 17739 37420
rect 17681 37411 17739 37417
rect 18046 37408 18052 37420
rect 18104 37408 18110 37460
rect 20346 37340 20352 37392
rect 20404 37380 20410 37392
rect 38013 37383 38071 37389
rect 38013 37380 38025 37383
rect 20404 37352 38025 37380
rect 20404 37340 20410 37352
rect 38013 37349 38025 37352
rect 38059 37349 38071 37383
rect 38013 37343 38071 37349
rect 3191 37284 3924 37312
rect 3973 37315 4031 37321
rect 3191 37281 3203 37284
rect 3145 37275 3203 37281
rect 3973 37281 3985 37315
rect 4019 37312 4031 37315
rect 4522 37312 4528 37324
rect 4019 37284 4528 37312
rect 4019 37281 4031 37284
rect 3973 37275 4031 37281
rect 4522 37272 4528 37284
rect 4580 37272 4586 37324
rect 5626 37272 5632 37324
rect 5684 37312 5690 37324
rect 5721 37315 5779 37321
rect 5721 37312 5733 37315
rect 5684 37284 5733 37312
rect 5684 37272 5690 37284
rect 5721 37281 5733 37284
rect 5767 37281 5779 37315
rect 10502 37312 10508 37324
rect 5721 37275 5779 37281
rect 7116 37284 10508 37312
rect 3421 37247 3479 37253
rect 3421 37213 3433 37247
rect 3467 37244 3479 37247
rect 3878 37244 3884 37256
rect 3467 37216 3884 37244
rect 3467 37213 3479 37216
rect 3421 37207 3479 37213
rect 3878 37204 3884 37216
rect 3936 37204 3942 37256
rect 5994 37204 6000 37256
rect 6052 37244 6058 37256
rect 7116 37244 7144 37284
rect 10502 37272 10508 37284
rect 10560 37312 10566 37324
rect 10597 37315 10655 37321
rect 10597 37312 10609 37315
rect 10560 37284 10609 37312
rect 10560 37272 10566 37284
rect 10597 37281 10609 37284
rect 10643 37281 10655 37315
rect 10597 37275 10655 37281
rect 11054 37272 11060 37324
rect 11112 37312 11118 37324
rect 11701 37315 11759 37321
rect 11701 37312 11713 37315
rect 11112 37284 11713 37312
rect 11112 37272 11118 37284
rect 11701 37281 11713 37284
rect 11747 37312 11759 37315
rect 12066 37312 12072 37324
rect 11747 37284 12072 37312
rect 11747 37281 11759 37284
rect 11701 37275 11759 37281
rect 12066 37272 12072 37284
rect 12124 37272 12130 37324
rect 14277 37315 14335 37321
rect 14277 37281 14289 37315
rect 14323 37281 14335 37315
rect 15565 37315 15623 37321
rect 15565 37312 15577 37315
rect 14277 37275 14335 37281
rect 15120 37284 15577 37312
rect 6052 37216 6097 37244
rect 6472 37216 7144 37244
rect 6052 37204 6058 37216
rect 2498 37136 2504 37188
rect 2556 37136 2562 37188
rect 3142 37136 3148 37188
rect 3200 37176 3206 37188
rect 3200 37148 4554 37176
rect 3200 37136 3206 37148
rect 5442 37136 5448 37188
rect 5500 37176 5506 37188
rect 6472 37176 6500 37216
rect 7190 37204 7196 37256
rect 7248 37204 7254 37256
rect 8570 37204 8576 37256
rect 8628 37244 8634 37256
rect 8628 37216 8673 37244
rect 8628 37204 8634 37216
rect 8754 37204 8760 37256
rect 8812 37244 8818 37256
rect 10873 37247 10931 37253
rect 8812 37216 9522 37244
rect 8812 37204 8818 37216
rect 10873 37213 10885 37247
rect 10919 37244 10931 37247
rect 11514 37244 11520 37256
rect 10919 37216 11520 37244
rect 10919 37213 10931 37216
rect 10873 37207 10931 37213
rect 11514 37204 11520 37216
rect 11572 37204 11578 37256
rect 11977 37247 12035 37253
rect 11977 37213 11989 37247
rect 12023 37244 12035 37247
rect 12023 37216 12434 37244
rect 12023 37213 12035 37216
rect 11977 37207 12035 37213
rect 5500 37148 6500 37176
rect 6549 37179 6607 37185
rect 5500 37136 5506 37148
rect 6549 37145 6561 37179
rect 6595 37176 6607 37179
rect 7006 37176 7012 37188
rect 6595 37148 7012 37176
rect 6595 37145 6607 37148
rect 6549 37139 6607 37145
rect 7006 37136 7012 37148
rect 7064 37136 7070 37188
rect 8404 37148 9260 37176
rect 1486 37068 1492 37120
rect 1544 37108 1550 37120
rect 1673 37111 1731 37117
rect 1673 37108 1685 37111
rect 1544 37080 1685 37108
rect 1544 37068 1550 37080
rect 1673 37077 1685 37080
rect 1719 37077 1731 37111
rect 1673 37071 1731 37077
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 8404 37108 8432 37148
rect 9122 37108 9128 37120
rect 5868 37080 8432 37108
rect 9083 37080 9128 37108
rect 5868 37068 5874 37080
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 9232 37108 9260 37148
rect 10594 37136 10600 37188
rect 10652 37176 10658 37188
rect 12406 37176 12434 37216
rect 12986 37204 12992 37256
rect 13044 37244 13050 37256
rect 13265 37247 13323 37253
rect 13265 37244 13277 37247
rect 13044 37216 13277 37244
rect 13044 37204 13050 37216
rect 13265 37213 13277 37216
rect 13311 37244 13323 37247
rect 14292 37244 14320 37275
rect 13311 37216 14320 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15120 37253 15148 37284
rect 15565 37281 15577 37284
rect 15611 37281 15623 37315
rect 18138 37312 18144 37324
rect 18099 37284 18144 37312
rect 15565 37275 15623 37281
rect 18138 37272 18144 37284
rect 18196 37272 18202 37324
rect 34333 37315 34391 37321
rect 34333 37281 34345 37315
rect 34379 37312 34391 37315
rect 34379 37284 34836 37312
rect 34379 37281 34391 37284
rect 34333 37275 34391 37281
rect 34808 37256 34836 37284
rect 15105 37247 15163 37253
rect 15105 37244 15117 37247
rect 14884 37216 15117 37244
rect 14884 37204 14890 37216
rect 15105 37213 15117 37216
rect 15151 37213 15163 37247
rect 15105 37207 15163 37213
rect 16758 37204 16764 37256
rect 16816 37244 16822 37256
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 16816 37216 17049 37244
rect 16816 37204 16822 37216
rect 17037 37213 17049 37216
rect 17083 37213 17095 37247
rect 17037 37207 17095 37213
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 18325 37207 18383 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 20898 37204 20904 37256
rect 20956 37244 20962 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 20956 37216 22017 37244
rect 20956 37204 20962 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22005 37207 22063 37213
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25314 37244 25320 37256
rect 25275 37216 25320 37244
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 26878 37204 26884 37256
rect 26936 37244 26942 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26936 37216 27169 37244
rect 26936 37204 26942 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 28626 37204 28632 37256
rect 28684 37244 28690 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 28684 37216 29745 37244
rect 28684 37204 28690 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31205 37247 31263 37253
rect 31205 37244 31217 37247
rect 30984 37216 31217 37244
rect 30984 37204 30990 37216
rect 31205 37213 31217 37216
rect 31251 37244 31263 37247
rect 31665 37247 31723 37253
rect 31665 37244 31677 37247
rect 31251 37216 31677 37244
rect 31251 37213 31263 37216
rect 31205 37207 31263 37213
rect 31665 37213 31677 37216
rect 31711 37213 31723 37247
rect 31665 37207 31723 37213
rect 32490 37204 32496 37256
rect 32548 37244 32554 37256
rect 32585 37247 32643 37253
rect 32585 37244 32597 37247
rect 32548 37216 32597 37244
rect 32548 37204 32554 37216
rect 32585 37213 32597 37216
rect 32631 37213 32643 37247
rect 32585 37207 32643 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34848 37216 34897 37244
rect 34848 37204 34854 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 36449 37247 36507 37253
rect 36449 37213 36461 37247
rect 36495 37213 36507 37247
rect 36449 37207 36507 37213
rect 37553 37247 37611 37253
rect 37553 37213 37565 37247
rect 37599 37244 37611 37247
rect 38010 37244 38016 37256
rect 37599 37216 38016 37244
rect 37599 37213 37611 37216
rect 37553 37207 37611 37213
rect 15194 37176 15200 37188
rect 10652 37148 10916 37176
rect 12406 37148 15200 37176
rect 10652 37136 10658 37148
rect 10778 37108 10784 37120
rect 9232 37080 10784 37108
rect 10778 37068 10784 37080
rect 10836 37068 10842 37120
rect 10888 37108 10916 37148
rect 15194 37136 15200 37148
rect 15252 37136 15258 37188
rect 36464 37176 36492 37207
rect 38010 37204 38016 37216
rect 38068 37244 38074 37256
rect 38197 37247 38255 37253
rect 38197 37244 38209 37247
rect 38068 37216 38209 37244
rect 38068 37204 38074 37216
rect 38197 37213 38209 37216
rect 38243 37213 38255 37247
rect 38197 37207 38255 37213
rect 37734 37176 37740 37188
rect 36464 37148 37740 37176
rect 37734 37136 37740 37148
rect 37792 37136 37798 37188
rect 12802 37108 12808 37120
rect 10888 37080 12808 37108
rect 12802 37068 12808 37080
rect 12860 37068 12866 37120
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13081 37111 13139 37117
rect 13081 37108 13093 37111
rect 12952 37080 13093 37108
rect 12952 37068 12958 37080
rect 13081 37077 13093 37080
rect 13127 37077 13139 37111
rect 14918 37108 14924 37120
rect 14879 37080 14924 37108
rect 13081 37071 13139 37077
rect 14918 37068 14924 37080
rect 14976 37068 14982 37120
rect 16942 37108 16948 37120
rect 16903 37080 16948 37108
rect 16942 37068 16948 37080
rect 17000 37068 17006 37120
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 22152 37080 22201 37108
rect 22152 37068 22158 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 23900 37080 24777 37108
rect 23900 37068 23906 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 25501 37071 25559 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 31018 37108 31024 37120
rect 30979 37080 31024 37108
rect 29917 37071 29975 37077
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32401 37111 32459 37117
rect 32401 37108 32413 37111
rect 32272 37080 32413 37108
rect 32272 37068 32278 37080
rect 32401 37077 32413 37080
rect 32447 37077 32459 37111
rect 32401 37071 32459 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 36136 37080 36277 37108
rect 36136 37068 36142 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 36265 37071 36323 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3878 36864 3884 36916
rect 3936 36904 3942 36916
rect 4890 36904 4896 36916
rect 3936 36876 4896 36904
rect 3936 36864 3942 36876
rect 4890 36864 4896 36876
rect 4948 36904 4954 36916
rect 5994 36904 6000 36916
rect 4948 36876 6000 36904
rect 4948 36864 4954 36876
rect 5994 36864 6000 36876
rect 6052 36864 6058 36916
rect 8570 36864 8576 36916
rect 8628 36904 8634 36916
rect 8628 36876 10732 36904
rect 8628 36864 8634 36876
rect 5810 36836 5816 36848
rect 4186 36808 5672 36836
rect 5771 36808 5816 36836
rect 1578 36768 1584 36780
rect 1539 36740 1584 36768
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 4890 36728 4896 36780
rect 4948 36768 4954 36780
rect 5644 36768 5672 36808
rect 5810 36796 5816 36808
rect 5868 36796 5874 36848
rect 6178 36796 6184 36848
rect 6236 36836 6242 36848
rect 6236 36808 7130 36836
rect 6236 36796 6242 36808
rect 9214 36796 9220 36848
rect 9272 36836 9278 36848
rect 10505 36839 10563 36845
rect 9272 36808 9338 36836
rect 9272 36796 9278 36808
rect 10505 36805 10517 36839
rect 10551 36836 10563 36839
rect 10594 36836 10600 36848
rect 10551 36808 10600 36836
rect 10551 36805 10563 36808
rect 10505 36799 10563 36805
rect 10594 36796 10600 36808
rect 10652 36796 10658 36848
rect 10704 36836 10732 36876
rect 10778 36864 10784 36916
rect 10836 36904 10842 36916
rect 14737 36907 14795 36913
rect 14737 36904 14749 36907
rect 10836 36876 14749 36904
rect 10836 36864 10842 36876
rect 14737 36873 14749 36876
rect 14783 36873 14795 36907
rect 14737 36867 14795 36873
rect 17037 36907 17095 36913
rect 17037 36873 17049 36907
rect 17083 36904 17095 36907
rect 20070 36904 20076 36916
rect 17083 36876 20076 36904
rect 17083 36873 17095 36876
rect 17037 36867 17095 36873
rect 20070 36864 20076 36876
rect 20128 36864 20134 36916
rect 32490 36904 32496 36916
rect 32451 36876 32496 36904
rect 32490 36864 32496 36876
rect 32548 36864 32554 36916
rect 38197 36907 38255 36913
rect 38197 36873 38209 36907
rect 38243 36904 38255 36907
rect 39298 36904 39304 36916
rect 38243 36876 39304 36904
rect 38243 36873 38255 36876
rect 38197 36867 38255 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 10704 36808 10824 36836
rect 5718 36768 5724 36780
rect 4948 36740 4993 36768
rect 5644 36740 5724 36768
rect 4948 36728 4954 36740
rect 5718 36728 5724 36740
rect 5776 36728 5782 36780
rect 10796 36777 10824 36808
rect 11054 36796 11060 36848
rect 11112 36836 11118 36848
rect 11977 36839 12035 36845
rect 11977 36836 11989 36839
rect 11112 36808 11989 36836
rect 11112 36796 11118 36808
rect 11977 36805 11989 36808
rect 12023 36805 12035 36839
rect 11977 36799 12035 36805
rect 10781 36771 10839 36777
rect 10781 36737 10793 36771
rect 10827 36768 10839 36771
rect 11514 36768 11520 36780
rect 10827 36740 11520 36768
rect 10827 36737 10839 36740
rect 10781 36731 10839 36737
rect 11514 36728 11520 36740
rect 11572 36768 11578 36780
rect 11701 36771 11759 36777
rect 11701 36768 11713 36771
rect 11572 36740 11713 36768
rect 11572 36728 11578 36740
rect 11701 36737 11713 36740
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 13078 36728 13084 36780
rect 13136 36728 13142 36780
rect 14277 36771 14335 36777
rect 14277 36737 14289 36771
rect 14323 36768 14335 36771
rect 14918 36768 14924 36780
rect 14323 36740 14924 36768
rect 14323 36737 14335 36740
rect 14277 36731 14335 36737
rect 14918 36728 14924 36740
rect 14976 36728 14982 36780
rect 15194 36728 15200 36780
rect 15252 36768 15258 36780
rect 16482 36768 16488 36780
rect 15252 36740 16488 36768
rect 15252 36728 15258 36740
rect 16482 36728 16488 36740
rect 16540 36768 16546 36780
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 16540 36740 16865 36768
rect 16540 36728 16546 36740
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 28169 36771 28227 36777
rect 28169 36737 28181 36771
rect 28215 36768 28227 36771
rect 31018 36768 31024 36780
rect 28215 36740 31024 36768
rect 28215 36737 28227 36740
rect 28169 36731 28227 36737
rect 31018 36728 31024 36740
rect 31076 36728 31082 36780
rect 32309 36771 32367 36777
rect 32309 36768 32321 36771
rect 31772 36740 32321 36768
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36700 1915 36703
rect 2130 36700 2136 36712
rect 1903 36672 2136 36700
rect 1903 36669 1915 36672
rect 1857 36663 1915 36669
rect 2130 36660 2136 36672
rect 2188 36660 2194 36712
rect 2869 36703 2927 36709
rect 2869 36669 2881 36703
rect 2915 36700 2927 36703
rect 3602 36700 3608 36712
rect 2915 36672 3608 36700
rect 2915 36669 2927 36672
rect 2869 36663 2927 36669
rect 3602 36660 3608 36672
rect 3660 36660 3666 36712
rect 4617 36703 4675 36709
rect 4617 36669 4629 36703
rect 4663 36700 4675 36703
rect 5534 36700 5540 36712
rect 4663 36672 5540 36700
rect 4663 36669 4675 36672
rect 4617 36663 4675 36669
rect 5534 36660 5540 36672
rect 5592 36660 5598 36712
rect 6546 36700 6552 36712
rect 6507 36672 6552 36700
rect 6546 36660 6552 36672
rect 6604 36660 6610 36712
rect 7006 36660 7012 36712
rect 7064 36700 7070 36712
rect 8294 36700 8300 36712
rect 7064 36672 8300 36700
rect 7064 36660 7070 36672
rect 8294 36660 8300 36672
rect 8352 36660 8358 36712
rect 8570 36700 8576 36712
rect 8531 36672 8576 36700
rect 8570 36660 8576 36672
rect 8628 36660 8634 36712
rect 8662 36660 8668 36712
rect 8720 36700 8726 36712
rect 9033 36703 9091 36709
rect 9033 36700 9045 36703
rect 8720 36672 9045 36700
rect 8720 36660 8726 36672
rect 9033 36669 9045 36672
rect 9079 36669 9091 36703
rect 9033 36663 9091 36669
rect 9306 36660 9312 36712
rect 9364 36700 9370 36712
rect 10502 36700 10508 36712
rect 9364 36672 10508 36700
rect 9364 36660 9370 36672
rect 10502 36660 10508 36672
rect 10560 36660 10566 36712
rect 13449 36703 13507 36709
rect 13449 36700 13461 36703
rect 10704 36672 13461 36700
rect 5997 36635 6055 36641
rect 5997 36601 6009 36635
rect 6043 36632 6055 36635
rect 6454 36632 6460 36644
rect 6043 36604 6460 36632
rect 6043 36601 6055 36604
rect 5997 36595 6055 36601
rect 6454 36592 6460 36604
rect 6512 36592 6518 36644
rect 7190 36524 7196 36576
rect 7248 36564 7254 36576
rect 10704 36564 10732 36672
rect 13449 36669 13461 36672
rect 13495 36700 13507 36703
rect 13538 36700 13544 36712
rect 13495 36672 13544 36700
rect 13495 36669 13507 36672
rect 13449 36663 13507 36669
rect 13538 36660 13544 36672
rect 13596 36660 13602 36712
rect 27890 36700 27896 36712
rect 27851 36672 27896 36700
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 16022 36592 16028 36644
rect 16080 36632 16086 36644
rect 31772 36641 31800 36740
rect 32309 36737 32321 36740
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 37553 36771 37611 36777
rect 37553 36737 37565 36771
rect 37599 36768 37611 36771
rect 37918 36768 37924 36780
rect 37599 36740 37924 36768
rect 37599 36737 37611 36740
rect 37553 36731 37611 36737
rect 37918 36728 37924 36740
rect 37976 36768 37982 36780
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 37976 36740 38025 36768
rect 37976 36728 37982 36740
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 31757 36635 31815 36641
rect 31757 36632 31769 36635
rect 16080 36604 31769 36632
rect 16080 36592 16086 36604
rect 31757 36601 31769 36604
rect 31803 36601 31815 36635
rect 31757 36595 31815 36601
rect 7248 36536 10732 36564
rect 7248 36524 7254 36536
rect 10962 36524 10968 36576
rect 11020 36564 11026 36576
rect 13170 36564 13176 36576
rect 11020 36536 13176 36564
rect 11020 36524 11026 36536
rect 13170 36524 13176 36536
rect 13228 36524 13234 36576
rect 14090 36564 14096 36576
rect 14051 36536 14096 36564
rect 14090 36524 14096 36536
rect 14148 36524 14154 36576
rect 15286 36564 15292 36576
rect 15247 36536 15292 36564
rect 15286 36524 15292 36536
rect 15344 36564 15350 36576
rect 15841 36567 15899 36573
rect 15841 36564 15853 36567
rect 15344 36536 15853 36564
rect 15344 36524 15350 36536
rect 15841 36533 15853 36536
rect 15887 36564 15899 36567
rect 15930 36564 15936 36576
rect 15887 36536 15936 36564
rect 15887 36533 15899 36536
rect 15841 36527 15899 36533
rect 15930 36524 15936 36536
rect 15988 36524 15994 36576
rect 25225 36567 25283 36573
rect 25225 36533 25237 36567
rect 25271 36564 25283 36567
rect 25314 36564 25320 36576
rect 25271 36536 25320 36564
rect 25271 36533 25283 36536
rect 25225 36527 25283 36533
rect 25314 36524 25320 36536
rect 25372 36524 25378 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2590 36320 2596 36372
rect 2648 36360 2654 36372
rect 4065 36363 4123 36369
rect 4065 36360 4077 36363
rect 2648 36332 4077 36360
rect 2648 36320 2654 36332
rect 4065 36329 4077 36332
rect 4111 36329 4123 36363
rect 14090 36360 14096 36372
rect 4065 36323 4123 36329
rect 4264 36332 14096 36360
rect 1673 36227 1731 36233
rect 1673 36193 1685 36227
rect 1719 36224 1731 36227
rect 3878 36224 3884 36236
rect 1719 36196 3884 36224
rect 1719 36193 1731 36196
rect 1673 36187 1731 36193
rect 3878 36184 3884 36196
rect 3936 36184 3942 36236
rect 3050 36116 3056 36168
rect 3108 36116 3114 36168
rect 4264 36165 4292 36332
rect 14090 36320 14096 36332
rect 14148 36320 14154 36372
rect 15930 36320 15936 36372
rect 15988 36360 15994 36372
rect 16485 36363 16543 36369
rect 16485 36360 16497 36363
rect 15988 36332 16497 36360
rect 15988 36320 15994 36332
rect 16485 36329 16497 36332
rect 16531 36329 16543 36363
rect 16485 36323 16543 36329
rect 5442 36292 5448 36304
rect 5184 36264 5448 36292
rect 4249 36159 4307 36165
rect 4249 36125 4261 36159
rect 4295 36125 4307 36159
rect 4249 36119 4307 36125
rect 1946 36088 1952 36100
rect 1907 36060 1952 36088
rect 1946 36048 1952 36060
rect 2004 36048 2010 36100
rect 4801 36091 4859 36097
rect 4801 36057 4813 36091
rect 4847 36088 4859 36091
rect 5074 36088 5080 36100
rect 4847 36060 5080 36088
rect 4847 36057 4859 36060
rect 4801 36051 4859 36057
rect 5074 36048 5080 36060
rect 5132 36048 5138 36100
rect 3421 36023 3479 36029
rect 3421 35989 3433 36023
rect 3467 36020 3479 36023
rect 5184 36020 5212 36264
rect 5442 36252 5448 36264
rect 5500 36252 5506 36304
rect 8294 36252 8300 36304
rect 8352 36292 8358 36304
rect 9582 36292 9588 36304
rect 8352 36264 9588 36292
rect 8352 36252 8358 36264
rect 9582 36252 9588 36264
rect 9640 36252 9646 36304
rect 10962 36292 10968 36304
rect 10796 36264 10968 36292
rect 10796 36224 10824 36264
rect 10962 36252 10968 36264
rect 11020 36252 11026 36304
rect 12066 36292 12072 36304
rect 12027 36264 12072 36292
rect 12066 36252 12072 36264
rect 12124 36252 12130 36304
rect 13170 36292 13176 36304
rect 13131 36264 13176 36292
rect 13170 36252 13176 36264
rect 13228 36292 13234 36304
rect 13998 36292 14004 36304
rect 13228 36264 14004 36292
rect 13228 36252 13234 36264
rect 13998 36252 14004 36264
rect 14056 36252 14062 36304
rect 27890 36292 27896 36304
rect 16546 36264 27896 36292
rect 8404 36196 10824 36224
rect 10873 36227 10931 36233
rect 5442 36116 5448 36168
rect 5500 36116 5506 36168
rect 6822 36116 6828 36168
rect 6880 36156 6886 36168
rect 7285 36159 7343 36165
rect 7285 36156 7297 36159
rect 6880 36128 7297 36156
rect 6880 36116 6886 36128
rect 7285 36125 7297 36128
rect 7331 36125 7343 36159
rect 7285 36119 7343 36125
rect 7742 36116 7748 36168
rect 7800 36156 7806 36168
rect 8021 36159 8079 36165
rect 8021 36156 8033 36159
rect 7800 36128 8033 36156
rect 7800 36116 7806 36128
rect 8021 36125 8033 36128
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 6549 36091 6607 36097
rect 6549 36057 6561 36091
rect 6595 36088 6607 36091
rect 6638 36088 6644 36100
rect 6595 36060 6644 36088
rect 6595 36057 6607 36060
rect 6549 36051 6607 36057
rect 6638 36048 6644 36060
rect 6696 36088 6702 36100
rect 8404 36088 8432 36196
rect 10873 36193 10885 36227
rect 10919 36224 10931 36227
rect 11514 36224 11520 36236
rect 10919 36196 11520 36224
rect 10919 36193 10931 36196
rect 10873 36187 10931 36193
rect 11514 36184 11520 36196
rect 11572 36224 11578 36236
rect 12621 36227 12679 36233
rect 12621 36224 12633 36227
rect 11572 36196 12633 36224
rect 11572 36184 11578 36196
rect 12621 36193 12633 36196
rect 12667 36224 12679 36227
rect 14829 36227 14887 36233
rect 14829 36224 14841 36227
rect 12667 36196 14841 36224
rect 12667 36193 12679 36196
rect 12621 36187 12679 36193
rect 14829 36193 14841 36196
rect 14875 36224 14887 36227
rect 15286 36224 15292 36236
rect 14875 36196 15292 36224
rect 14875 36193 14887 36196
rect 14829 36187 14887 36193
rect 15286 36184 15292 36196
rect 15344 36224 15350 36236
rect 15381 36227 15439 36233
rect 15381 36224 15393 36227
rect 15344 36196 15393 36224
rect 15344 36184 15350 36196
rect 15381 36193 15393 36196
rect 15427 36193 15439 36227
rect 15381 36187 15439 36193
rect 8478 36116 8484 36168
rect 8536 36156 8542 36168
rect 9214 36156 9220 36168
rect 8536 36128 9220 36156
rect 8536 36116 8542 36128
rect 9214 36116 9220 36128
rect 9272 36116 9278 36168
rect 9490 36116 9496 36168
rect 9548 36116 9554 36168
rect 10962 36116 10968 36168
rect 11020 36156 11026 36168
rect 16546 36156 16574 36264
rect 27890 36252 27896 36264
rect 27948 36252 27954 36304
rect 11020 36128 16574 36156
rect 11020 36116 11026 36128
rect 6696 36060 8432 36088
rect 8573 36091 8631 36097
rect 6696 36048 6702 36060
rect 8573 36057 8585 36091
rect 8619 36088 8631 36091
rect 10597 36091 10655 36097
rect 8619 36060 9352 36088
rect 8619 36057 8631 36060
rect 8573 36051 8631 36057
rect 3467 35992 5212 36020
rect 3467 35989 3479 35992
rect 3421 35983 3479 35989
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 7837 36023 7895 36029
rect 7837 36020 7849 36023
rect 5592 35992 7849 36020
rect 5592 35980 5598 35992
rect 7837 35989 7849 35992
rect 7883 35989 7895 36023
rect 7837 35983 7895 35989
rect 7926 35980 7932 36032
rect 7984 36020 7990 36032
rect 8588 36020 8616 36051
rect 7984 35992 8616 36020
rect 9125 36023 9183 36029
rect 7984 35980 7990 35992
rect 9125 35989 9137 36023
rect 9171 36020 9183 36023
rect 9214 36020 9220 36032
rect 9171 35992 9220 36020
rect 9171 35989 9183 35992
rect 9125 35983 9183 35989
rect 9214 35980 9220 35992
rect 9272 35980 9278 36032
rect 9324 36020 9352 36060
rect 10597 36057 10609 36091
rect 10643 36088 10655 36091
rect 11698 36088 11704 36100
rect 10643 36060 11704 36088
rect 10643 36057 10655 36060
rect 10597 36051 10655 36057
rect 10704 36020 10732 36060
rect 11698 36048 11704 36060
rect 11756 36048 11762 36100
rect 12802 36048 12808 36100
rect 12860 36088 12866 36100
rect 15933 36091 15991 36097
rect 15933 36088 15945 36091
rect 12860 36060 15945 36088
rect 12860 36048 12866 36060
rect 15933 36057 15945 36060
rect 15979 36088 15991 36091
rect 16850 36088 16856 36100
rect 15979 36060 16856 36088
rect 15979 36057 15991 36060
rect 15933 36051 15991 36057
rect 16850 36048 16856 36060
rect 16908 36048 16914 36100
rect 37553 36091 37611 36097
rect 37553 36057 37565 36091
rect 37599 36088 37611 36091
rect 38194 36088 38200 36100
rect 37599 36060 38200 36088
rect 37599 36057 37611 36060
rect 37553 36051 37611 36057
rect 38194 36048 38200 36060
rect 38252 36048 38258 36100
rect 9324 35992 10732 36020
rect 10870 35980 10876 36032
rect 10928 36020 10934 36032
rect 14277 36023 14335 36029
rect 14277 36020 14289 36023
rect 10928 35992 14289 36020
rect 10928 35980 10934 35992
rect 14277 35989 14289 35992
rect 14323 35989 14335 36023
rect 38102 36020 38108 36032
rect 38063 35992 38108 36020
rect 14277 35983 14335 35989
rect 38102 35980 38108 35992
rect 38160 35980 38166 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 4062 35776 4068 35828
rect 4120 35816 4126 35828
rect 11057 35819 11115 35825
rect 11057 35816 11069 35819
rect 4120 35788 9076 35816
rect 4120 35776 4126 35788
rect 1946 35748 1952 35760
rect 1907 35720 1952 35748
rect 1946 35708 1952 35720
rect 2004 35708 2010 35760
rect 2222 35708 2228 35760
rect 2280 35748 2286 35760
rect 4540 35757 4568 35788
rect 4525 35751 4583 35757
rect 2280 35720 2530 35748
rect 2280 35708 2286 35720
rect 4525 35717 4537 35751
rect 4571 35717 4583 35751
rect 4525 35711 4583 35717
rect 4709 35751 4767 35757
rect 4709 35717 4721 35751
rect 4755 35748 4767 35751
rect 5994 35748 6000 35760
rect 4755 35720 6000 35748
rect 4755 35717 4767 35720
rect 4709 35711 4767 35717
rect 5994 35708 6000 35720
rect 6052 35708 6058 35760
rect 6086 35708 6092 35760
rect 6144 35748 6150 35760
rect 6144 35720 7590 35748
rect 6144 35708 6150 35720
rect 3970 35640 3976 35692
rect 4028 35680 4034 35692
rect 5353 35683 5411 35689
rect 4028 35652 4073 35680
rect 4028 35640 4034 35652
rect 5353 35649 5365 35683
rect 5399 35680 5411 35683
rect 5534 35680 5540 35692
rect 5399 35652 5540 35680
rect 5399 35649 5411 35652
rect 5353 35643 5411 35649
rect 5534 35640 5540 35652
rect 5592 35640 5598 35692
rect 9048 35680 9076 35788
rect 9876 35788 11069 35816
rect 9582 35708 9588 35760
rect 9640 35748 9646 35760
rect 9876 35748 9904 35788
rect 11057 35785 11069 35788
rect 11103 35785 11115 35819
rect 11057 35779 11115 35785
rect 15657 35819 15715 35825
rect 15657 35785 15669 35819
rect 15703 35816 15715 35819
rect 15930 35816 15936 35828
rect 15703 35788 15936 35816
rect 15703 35785 15715 35788
rect 15657 35779 15715 35785
rect 15930 35776 15936 35788
rect 15988 35776 15994 35828
rect 23293 35819 23351 35825
rect 23293 35785 23305 35819
rect 23339 35816 23351 35819
rect 24578 35816 24584 35828
rect 23339 35788 24584 35816
rect 23339 35785 23351 35788
rect 23293 35779 23351 35785
rect 24578 35776 24584 35788
rect 24636 35776 24642 35828
rect 38197 35819 38255 35825
rect 38197 35785 38209 35819
rect 38243 35816 38255 35819
rect 38286 35816 38292 35828
rect 38243 35788 38292 35816
rect 38243 35785 38255 35788
rect 38197 35779 38255 35785
rect 38286 35776 38292 35788
rect 38344 35776 38350 35828
rect 14458 35748 14464 35760
rect 9640 35720 9904 35748
rect 14419 35720 14464 35748
rect 9640 35708 9646 35720
rect 14458 35708 14464 35720
rect 14516 35708 14522 35760
rect 9950 35680 9956 35692
rect 9048 35652 9956 35680
rect 9950 35640 9956 35652
rect 10008 35640 10014 35692
rect 10045 35683 10103 35689
rect 10045 35649 10057 35683
rect 10091 35680 10103 35683
rect 12253 35683 12311 35689
rect 12253 35680 12265 35683
rect 10091 35652 12265 35680
rect 10091 35649 10103 35652
rect 10045 35643 10103 35649
rect 12253 35649 12265 35652
rect 12299 35649 12311 35683
rect 12253 35643 12311 35649
rect 12342 35640 12348 35692
rect 12400 35678 12406 35692
rect 23106 35680 23112 35692
rect 12400 35650 12443 35678
rect 23067 35652 23112 35680
rect 12400 35640 12406 35650
rect 23106 35640 23112 35652
rect 23164 35680 23170 35692
rect 23753 35683 23811 35689
rect 23753 35680 23765 35683
rect 23164 35652 23765 35680
rect 23164 35640 23170 35652
rect 23753 35649 23765 35652
rect 23799 35649 23811 35683
rect 23753 35643 23811 35649
rect 37550 35640 37556 35692
rect 37608 35680 37614 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37608 35652 38025 35680
rect 37608 35640 37614 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 3697 35615 3755 35621
rect 3697 35581 3709 35615
rect 3743 35612 3755 35615
rect 3988 35612 4016 35640
rect 6549 35615 6607 35621
rect 6549 35612 6561 35615
rect 3743 35584 3924 35612
rect 3988 35584 6561 35612
rect 3743 35581 3755 35584
rect 3697 35575 3755 35581
rect 3896 35544 3924 35584
rect 6549 35581 6561 35584
rect 6595 35612 6607 35615
rect 6822 35612 6828 35624
rect 6595 35584 6828 35612
rect 6595 35581 6607 35584
rect 6549 35575 6607 35581
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 7282 35612 7288 35624
rect 7243 35584 7288 35612
rect 7282 35572 7288 35584
rect 7340 35612 7346 35624
rect 8202 35612 8208 35624
rect 7340 35584 8208 35612
rect 7340 35572 7346 35584
rect 8202 35572 8208 35584
rect 8260 35572 8266 35624
rect 8386 35572 8392 35624
rect 8444 35612 8450 35624
rect 8757 35615 8815 35621
rect 8757 35612 8769 35615
rect 8444 35584 8769 35612
rect 8444 35572 8450 35584
rect 8757 35581 8769 35584
rect 8803 35581 8815 35615
rect 9030 35612 9036 35624
rect 8991 35584 9036 35612
rect 8757 35575 8815 35581
rect 9030 35572 9036 35584
rect 9088 35612 9094 35624
rect 10505 35615 10563 35621
rect 10505 35612 10517 35615
rect 9088 35584 10517 35612
rect 9088 35572 9094 35584
rect 10505 35581 10517 35584
rect 10551 35581 10563 35615
rect 15013 35615 15071 35621
rect 15013 35612 15025 35615
rect 10505 35575 10563 35581
rect 10704 35584 15025 35612
rect 4614 35544 4620 35556
rect 3896 35516 4620 35544
rect 4614 35504 4620 35516
rect 4672 35544 4678 35556
rect 4672 35516 6684 35544
rect 4672 35504 4678 35516
rect 4706 35436 4712 35488
rect 4764 35476 4770 35488
rect 5169 35479 5227 35485
rect 5169 35476 5181 35479
rect 4764 35448 5181 35476
rect 4764 35436 4770 35448
rect 5169 35445 5181 35448
rect 5215 35445 5227 35479
rect 5902 35476 5908 35488
rect 5863 35448 5908 35476
rect 5169 35439 5227 35445
rect 5902 35436 5908 35448
rect 5960 35436 5966 35488
rect 6656 35476 6684 35516
rect 9674 35504 9680 35556
rect 9732 35544 9738 35556
rect 9861 35547 9919 35553
rect 9861 35544 9873 35547
rect 9732 35516 9873 35544
rect 9732 35504 9738 35516
rect 9861 35513 9873 35516
rect 9907 35513 9919 35547
rect 9861 35507 9919 35513
rect 10704 35476 10732 35584
rect 15013 35581 15025 35584
rect 15059 35612 15071 35615
rect 16298 35612 16304 35624
rect 15059 35584 16304 35612
rect 15059 35581 15071 35584
rect 15013 35575 15071 35581
rect 16298 35572 16304 35584
rect 16356 35572 16362 35624
rect 10778 35504 10784 35556
rect 10836 35544 10842 35556
rect 13909 35547 13967 35553
rect 13909 35544 13921 35547
rect 10836 35516 13921 35544
rect 10836 35504 10842 35516
rect 13909 35513 13921 35516
rect 13955 35544 13967 35547
rect 14366 35544 14372 35556
rect 13955 35516 14372 35544
rect 13955 35513 13967 35516
rect 13909 35507 13967 35513
rect 14366 35504 14372 35516
rect 14424 35504 14430 35556
rect 6656 35448 10732 35476
rect 12897 35479 12955 35485
rect 12897 35445 12909 35479
rect 12943 35476 12955 35479
rect 13446 35476 13452 35488
rect 12943 35448 13452 35476
rect 12943 35445 12955 35448
rect 12897 35439 12955 35445
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 658 35232 664 35284
rect 716 35272 722 35284
rect 4065 35275 4123 35281
rect 4065 35272 4077 35275
rect 716 35244 4077 35272
rect 716 35232 722 35244
rect 4065 35241 4077 35244
rect 4111 35241 4123 35275
rect 4065 35235 4123 35241
rect 5920 35244 7144 35272
rect 3421 35139 3479 35145
rect 3421 35105 3433 35139
rect 3467 35136 3479 35139
rect 3878 35136 3884 35148
rect 3467 35108 3884 35136
rect 3467 35105 3479 35108
rect 3421 35099 3479 35105
rect 3878 35096 3884 35108
rect 3936 35096 3942 35148
rect 5169 35139 5227 35145
rect 5169 35105 5181 35139
rect 5215 35136 5227 35139
rect 5626 35136 5632 35148
rect 5215 35108 5632 35136
rect 5215 35105 5227 35108
rect 5169 35099 5227 35105
rect 5626 35096 5632 35108
rect 5684 35136 5690 35148
rect 5920 35136 5948 35244
rect 7116 35204 7144 35244
rect 7742 35232 7748 35284
rect 7800 35272 7806 35284
rect 10962 35272 10968 35284
rect 7800 35244 10968 35272
rect 7800 35232 7806 35244
rect 10962 35232 10968 35244
rect 11020 35232 11026 35284
rect 13173 35275 13231 35281
rect 13173 35241 13185 35275
rect 13219 35272 13231 35275
rect 13446 35272 13452 35284
rect 13219 35244 13452 35272
rect 13219 35241 13231 35244
rect 13173 35235 13231 35241
rect 13446 35232 13452 35244
rect 13504 35272 13510 35284
rect 13725 35275 13783 35281
rect 13725 35272 13737 35275
rect 13504 35244 13737 35272
rect 13504 35232 13510 35244
rect 13725 35241 13737 35244
rect 13771 35272 13783 35275
rect 14369 35275 14427 35281
rect 14369 35272 14381 35275
rect 13771 35244 14381 35272
rect 13771 35241 13783 35244
rect 13725 35235 13783 35241
rect 14369 35241 14381 35244
rect 14415 35272 14427 35275
rect 15930 35272 15936 35284
rect 14415 35244 15936 35272
rect 14415 35241 14427 35244
rect 14369 35235 14427 35241
rect 15930 35232 15936 35244
rect 15988 35232 15994 35284
rect 7116 35176 9260 35204
rect 5684 35108 5948 35136
rect 5684 35096 5690 35108
rect 6822 35096 6828 35148
rect 6880 35136 6886 35148
rect 7193 35139 7251 35145
rect 7193 35136 7205 35139
rect 6880 35108 7205 35136
rect 6880 35096 6886 35108
rect 7193 35105 7205 35108
rect 7239 35136 7251 35139
rect 7929 35139 7987 35145
rect 7929 35136 7941 35139
rect 7239 35108 7941 35136
rect 7239 35105 7251 35108
rect 7193 35099 7251 35105
rect 7929 35105 7941 35108
rect 7975 35136 7987 35139
rect 8294 35136 8300 35148
rect 7975 35108 8300 35136
rect 7975 35105 7987 35108
rect 7929 35099 7987 35105
rect 8294 35096 8300 35108
rect 8352 35136 8358 35148
rect 8481 35139 8539 35145
rect 8481 35136 8493 35139
rect 8352 35108 8493 35136
rect 8352 35096 8358 35108
rect 8481 35105 8493 35108
rect 8527 35136 8539 35139
rect 8570 35136 8576 35148
rect 8527 35108 8576 35136
rect 8527 35105 8539 35108
rect 8481 35099 8539 35105
rect 8570 35096 8576 35108
rect 8628 35136 8634 35148
rect 9030 35136 9036 35148
rect 8628 35108 9036 35136
rect 8628 35096 8634 35108
rect 9030 35096 9036 35108
rect 9088 35136 9094 35148
rect 9125 35139 9183 35145
rect 9125 35136 9137 35139
rect 9088 35108 9137 35136
rect 9088 35096 9094 35108
rect 9125 35105 9137 35108
rect 9171 35105 9183 35139
rect 9232 35136 9260 35176
rect 10410 35164 10416 35216
rect 10468 35204 10474 35216
rect 10468 35176 12480 35204
rect 10468 35164 10474 35176
rect 10778 35136 10784 35148
rect 9232 35108 10784 35136
rect 9125 35099 9183 35105
rect 10778 35096 10784 35108
rect 10836 35096 10842 35148
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35068 4307 35071
rect 4706 35068 4712 35080
rect 4295 35040 4712 35068
rect 4295 35037 4307 35040
rect 4249 35031 4307 35037
rect 4706 35028 4712 35040
rect 4764 35028 4770 35080
rect 12452 35077 12480 35176
rect 11793 35071 11851 35077
rect 11793 35068 11805 35071
rect 10704 35040 11805 35068
rect 2682 34960 2688 35012
rect 2740 34960 2746 35012
rect 3145 35003 3203 35009
rect 3145 34969 3157 35003
rect 3191 35000 3203 35003
rect 3191 34972 3372 35000
rect 3191 34969 3203 34972
rect 3145 34963 3203 34969
rect 1673 34935 1731 34941
rect 1673 34901 1685 34935
rect 1719 34932 1731 34935
rect 1854 34932 1860 34944
rect 1719 34904 1860 34932
rect 1719 34901 1731 34904
rect 1673 34895 1731 34901
rect 1854 34892 1860 34904
rect 1912 34892 1918 34944
rect 3344 34932 3372 34972
rect 3418 34960 3424 35012
rect 3476 35000 3482 35012
rect 6917 35003 6975 35009
rect 3476 34972 5750 35000
rect 3476 34960 3482 34972
rect 6917 34969 6929 35003
rect 6963 34969 6975 35003
rect 6917 34963 6975 34969
rect 3694 34932 3700 34944
rect 3344 34904 3700 34932
rect 3694 34892 3700 34904
rect 3752 34892 3758 34944
rect 6932 34932 6960 34963
rect 8570 34960 8576 35012
rect 8628 35000 8634 35012
rect 9122 35000 9128 35012
rect 8628 34972 9128 35000
rect 8628 34960 8634 34972
rect 9122 34960 9128 34972
rect 9180 35000 9186 35012
rect 9180 34972 9352 35000
rect 9180 34960 9186 34972
rect 8846 34932 8852 34944
rect 6932 34904 8852 34932
rect 8846 34892 8852 34904
rect 8904 34892 8910 34944
rect 9324 34932 9352 34972
rect 9398 34960 9404 35012
rect 9456 35000 9462 35012
rect 9456 34972 9501 35000
rect 9456 34960 9462 34972
rect 9858 34960 9864 35012
rect 9916 34960 9922 35012
rect 10704 34932 10732 35040
rect 11793 35037 11805 35040
rect 11839 35037 11851 35071
rect 11793 35031 11851 35037
rect 12437 35071 12495 35077
rect 12437 35037 12449 35071
rect 12483 35037 12495 35071
rect 12437 35031 12495 35037
rect 11885 35003 11943 35009
rect 11885 34969 11897 35003
rect 11931 35000 11943 35003
rect 15010 35000 15016 35012
rect 11931 34972 15016 35000
rect 11931 34969 11943 34972
rect 11885 34963 11943 34969
rect 15010 34960 15016 34972
rect 15068 34960 15074 35012
rect 9324 34904 10732 34932
rect 10778 34892 10784 34944
rect 10836 34932 10842 34944
rect 10873 34935 10931 34941
rect 10873 34932 10885 34935
rect 10836 34904 10885 34932
rect 10836 34892 10842 34904
rect 10873 34901 10885 34904
rect 10919 34901 10931 34935
rect 10873 34895 10931 34901
rect 12529 34935 12587 34941
rect 12529 34901 12541 34935
rect 12575 34932 12587 34935
rect 15102 34932 15108 34944
rect 12575 34904 15108 34932
rect 12575 34901 12587 34904
rect 12529 34895 12587 34901
rect 15102 34892 15108 34904
rect 15160 34892 15166 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2038 34688 2044 34740
rect 2096 34688 2102 34740
rect 2406 34688 2412 34740
rect 2464 34728 2470 34740
rect 2464 34700 3556 34728
rect 2464 34688 2470 34700
rect 2056 34660 2084 34688
rect 2225 34663 2283 34669
rect 2225 34660 2237 34663
rect 2056 34632 2237 34660
rect 2225 34629 2237 34632
rect 2271 34629 2283 34663
rect 2225 34623 2283 34629
rect 3528 34592 3556 34700
rect 3878 34688 3884 34740
rect 3936 34728 3942 34740
rect 5077 34731 5135 34737
rect 5077 34728 5089 34731
rect 3936 34700 5089 34728
rect 3936 34688 3942 34700
rect 5077 34697 5089 34700
rect 5123 34697 5135 34731
rect 5077 34691 5135 34697
rect 4617 34595 4675 34601
rect 4617 34592 4629 34595
rect 1949 34527 2007 34533
rect 1949 34493 1961 34527
rect 1995 34493 2007 34527
rect 3344 34524 3372 34578
rect 3528 34564 4629 34592
rect 4617 34561 4629 34564
rect 4663 34561 4675 34595
rect 5092 34592 5120 34691
rect 5534 34688 5540 34740
rect 5592 34728 5598 34740
rect 5592 34700 8156 34728
rect 5592 34688 5598 34700
rect 5166 34620 5172 34672
rect 5224 34660 5230 34672
rect 8128 34660 8156 34700
rect 9030 34688 9036 34740
rect 9088 34728 9094 34740
rect 9088 34700 10640 34728
rect 9088 34688 9094 34700
rect 5224 34632 7314 34660
rect 8128 34632 9154 34660
rect 5224 34620 5230 34632
rect 10612 34601 10640 34700
rect 10962 34688 10968 34740
rect 11020 34728 11026 34740
rect 11057 34731 11115 34737
rect 11057 34728 11069 34731
rect 11020 34700 11069 34728
rect 11020 34688 11026 34700
rect 11057 34697 11069 34700
rect 11103 34697 11115 34731
rect 11057 34691 11115 34697
rect 11146 34688 11152 34740
rect 11204 34728 11210 34740
rect 11330 34728 11336 34740
rect 11204 34700 11336 34728
rect 11204 34688 11210 34700
rect 11330 34688 11336 34700
rect 11388 34728 11394 34740
rect 13081 34731 13139 34737
rect 11388 34700 12434 34728
rect 11388 34688 11394 34700
rect 11974 34660 11980 34672
rect 11935 34632 11980 34660
rect 11974 34620 11980 34632
rect 12032 34620 12038 34672
rect 12406 34660 12434 34700
rect 13081 34697 13093 34731
rect 13127 34728 13139 34731
rect 13446 34728 13452 34740
rect 13127 34700 13452 34728
rect 13127 34697 13139 34700
rect 13081 34691 13139 34697
rect 13446 34688 13452 34700
rect 13504 34688 13510 34740
rect 14093 34663 14151 34669
rect 14093 34660 14105 34663
rect 12406 34632 14105 34660
rect 14093 34629 14105 34632
rect 14139 34629 14151 34663
rect 14093 34623 14151 34629
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 5092 34564 6561 34592
rect 4617 34555 4675 34561
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 10597 34595 10655 34601
rect 10597 34561 10609 34595
rect 10643 34561 10655 34595
rect 10597 34555 10655 34561
rect 3510 34524 3516 34536
rect 3344 34496 3516 34524
rect 1949 34487 2007 34493
rect 1670 34348 1676 34400
rect 1728 34388 1734 34400
rect 1964 34388 1992 34487
rect 3510 34484 3516 34496
rect 3568 34484 3574 34536
rect 3973 34527 4031 34533
rect 3973 34493 3985 34527
rect 4019 34524 4031 34527
rect 4798 34524 4804 34536
rect 4019 34496 4804 34524
rect 4019 34493 4031 34496
rect 3973 34487 4031 34493
rect 4798 34484 4804 34496
rect 4856 34484 4862 34536
rect 5902 34484 5908 34536
rect 5960 34524 5966 34536
rect 5997 34527 6055 34533
rect 5997 34524 6009 34527
rect 5960 34496 6009 34524
rect 5960 34484 5966 34496
rect 5997 34493 6009 34496
rect 6043 34524 6055 34527
rect 6822 34524 6828 34536
rect 6043 34496 6828 34524
rect 6043 34493 6055 34496
rect 5997 34487 6055 34493
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 9950 34524 9956 34536
rect 9324 34496 9956 34524
rect 8297 34459 8355 34465
rect 8297 34425 8309 34459
rect 8343 34456 8355 34459
rect 8386 34456 8392 34468
rect 8343 34428 8392 34456
rect 8343 34425 8355 34428
rect 8297 34419 8355 34425
rect 8386 34416 8392 34428
rect 8444 34456 8450 34468
rect 9324 34456 9352 34496
rect 9950 34484 9956 34496
rect 10008 34484 10014 34536
rect 11885 34527 11943 34533
rect 11885 34493 11897 34527
rect 11931 34524 11943 34527
rect 12342 34524 12348 34536
rect 11931 34496 12112 34524
rect 12303 34496 12348 34524
rect 11931 34493 11943 34496
rect 11885 34487 11943 34493
rect 8444 34428 9352 34456
rect 12084 34456 12112 34496
rect 12342 34484 12348 34496
rect 12400 34484 12406 34536
rect 13633 34527 13691 34533
rect 13633 34493 13645 34527
rect 13679 34524 13691 34527
rect 13814 34524 13820 34536
rect 13679 34496 13820 34524
rect 13679 34493 13691 34496
rect 13633 34487 13691 34493
rect 13814 34484 13820 34496
rect 13872 34484 13878 34536
rect 37826 34484 37832 34536
rect 37884 34524 37890 34536
rect 38013 34527 38071 34533
rect 38013 34524 38025 34527
rect 37884 34496 38025 34524
rect 37884 34484 37890 34496
rect 38013 34493 38025 34496
rect 38059 34493 38071 34527
rect 38286 34524 38292 34536
rect 38247 34496 38292 34524
rect 38013 34487 38071 34493
rect 38286 34484 38292 34496
rect 38344 34484 38350 34536
rect 12434 34456 12440 34468
rect 12084 34428 12440 34456
rect 8444 34416 8450 34428
rect 12434 34416 12440 34428
rect 12492 34416 12498 34468
rect 3878 34388 3884 34400
rect 1728 34360 3884 34388
rect 1728 34348 1734 34360
rect 3878 34348 3884 34360
rect 3936 34348 3942 34400
rect 4433 34391 4491 34397
rect 4433 34357 4445 34391
rect 4479 34388 4491 34391
rect 4614 34388 4620 34400
rect 4479 34360 4620 34388
rect 4479 34357 4491 34360
rect 4433 34351 4491 34357
rect 4614 34348 4620 34360
rect 4672 34348 4678 34400
rect 6812 34391 6870 34397
rect 6812 34357 6824 34391
rect 6858 34388 6870 34391
rect 6914 34388 6920 34400
rect 6858 34360 6920 34388
rect 6858 34357 6870 34360
rect 6812 34351 6870 34357
rect 6914 34348 6920 34360
rect 6972 34348 6978 34400
rect 8846 34388 8852 34400
rect 8759 34360 8852 34388
rect 8846 34348 8852 34360
rect 8904 34388 8910 34400
rect 9950 34388 9956 34400
rect 8904 34360 9956 34388
rect 8904 34348 8910 34360
rect 9950 34348 9956 34360
rect 10008 34348 10014 34400
rect 10226 34348 10232 34400
rect 10284 34388 10290 34400
rect 10333 34391 10391 34397
rect 10333 34388 10345 34391
rect 10284 34360 10345 34388
rect 10284 34348 10290 34360
rect 10333 34357 10345 34360
rect 10379 34357 10391 34391
rect 10333 34351 10391 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 8021 34187 8079 34193
rect 8021 34153 8033 34187
rect 8067 34184 8079 34187
rect 8294 34184 8300 34196
rect 8067 34156 8300 34184
rect 8067 34153 8079 34156
rect 8021 34147 8079 34153
rect 8294 34144 8300 34156
rect 8352 34184 8358 34196
rect 8481 34187 8539 34193
rect 8481 34184 8493 34187
rect 8352 34156 8493 34184
rect 8352 34144 8358 34156
rect 8481 34153 8493 34156
rect 8527 34153 8539 34187
rect 10873 34187 10931 34193
rect 8481 34147 8539 34153
rect 8588 34156 10456 34184
rect 7469 34119 7527 34125
rect 7469 34085 7481 34119
rect 7515 34116 7527 34119
rect 8588 34116 8616 34156
rect 7515 34088 8616 34116
rect 10428 34116 10456 34156
rect 10873 34153 10885 34187
rect 10919 34184 10931 34187
rect 11054 34184 11060 34196
rect 10919 34156 11060 34184
rect 10919 34153 10931 34156
rect 10873 34147 10931 34153
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 13998 34116 14004 34128
rect 10428 34088 14004 34116
rect 7515 34085 7527 34088
rect 7469 34079 7527 34085
rect 1670 34048 1676 34060
rect 1631 34020 1676 34048
rect 1670 34008 1676 34020
rect 1728 34008 1734 34060
rect 1949 34051 2007 34057
rect 1949 34017 1961 34051
rect 1995 34048 2007 34051
rect 3786 34048 3792 34060
rect 1995 34020 3792 34048
rect 1995 34017 2007 34020
rect 1949 34011 2007 34017
rect 3786 34008 3792 34020
rect 3844 34008 3850 34060
rect 3878 34008 3884 34060
rect 3936 34048 3942 34060
rect 4893 34051 4951 34057
rect 4893 34048 4905 34051
rect 3936 34020 4905 34048
rect 3936 34008 3942 34020
rect 4893 34017 4905 34020
rect 4939 34017 4951 34051
rect 5166 34048 5172 34060
rect 5079 34020 5172 34048
rect 4893 34011 4951 34017
rect 5166 34008 5172 34020
rect 5224 34048 5230 34060
rect 7484 34048 7512 34079
rect 13998 34076 14004 34088
rect 14056 34076 14062 34128
rect 38286 34116 38292 34128
rect 38247 34088 38292 34116
rect 38286 34076 38292 34088
rect 38344 34076 38350 34128
rect 5224 34020 7512 34048
rect 5224 34008 5230 34020
rect 8386 34008 8392 34060
rect 8444 34048 8450 34060
rect 9125 34051 9183 34057
rect 9125 34048 9137 34051
rect 8444 34020 9137 34048
rect 8444 34008 8450 34020
rect 9125 34017 9137 34020
rect 9171 34017 9183 34051
rect 9125 34011 9183 34017
rect 11701 34051 11759 34057
rect 11701 34017 11713 34051
rect 11747 34048 11759 34051
rect 14734 34048 14740 34060
rect 11747 34020 14740 34048
rect 11747 34017 11759 34020
rect 11701 34011 11759 34017
rect 14734 34008 14740 34020
rect 14792 34008 14798 34060
rect 4430 33980 4436 33992
rect 4391 33952 4436 33980
rect 4430 33940 4436 33952
rect 4488 33940 4494 33992
rect 6638 33940 6644 33992
rect 6696 33980 6702 33992
rect 6917 33983 6975 33989
rect 6917 33980 6929 33983
rect 6696 33952 6929 33980
rect 6696 33940 6702 33952
rect 6917 33949 6929 33952
rect 6963 33949 6975 33983
rect 6917 33943 6975 33949
rect 12805 33983 12863 33989
rect 12805 33949 12817 33983
rect 12851 33949 12863 33983
rect 13538 33980 13544 33992
rect 13499 33952 13544 33980
rect 12805 33943 12863 33949
rect 2958 33872 2964 33924
rect 3016 33872 3022 33924
rect 4157 33915 4215 33921
rect 4157 33881 4169 33915
rect 4203 33912 4215 33915
rect 5074 33912 5080 33924
rect 4203 33884 5080 33912
rect 4203 33881 4215 33884
rect 4157 33875 4215 33881
rect 5074 33872 5080 33884
rect 5132 33872 5138 33924
rect 5718 33872 5724 33924
rect 5776 33872 5782 33924
rect 8202 33872 8208 33924
rect 8260 33912 8266 33924
rect 9306 33912 9312 33924
rect 8260 33884 9312 33912
rect 8260 33872 8266 33884
rect 9306 33872 9312 33884
rect 9364 33912 9370 33924
rect 9401 33915 9459 33921
rect 9401 33912 9413 33915
rect 9364 33884 9413 33912
rect 9364 33872 9370 33884
rect 9401 33881 9413 33884
rect 9447 33881 9459 33915
rect 9401 33875 9459 33881
rect 9858 33872 9864 33924
rect 9916 33872 9922 33924
rect 11790 33912 11796 33924
rect 11751 33884 11796 33912
rect 11790 33872 11796 33884
rect 11848 33872 11854 33924
rect 12342 33912 12348 33924
rect 12303 33884 12348 33912
rect 12342 33872 12348 33884
rect 12400 33872 12406 33924
rect 3421 33847 3479 33853
rect 3421 33813 3433 33847
rect 3467 33844 3479 33847
rect 7466 33844 7472 33856
rect 3467 33816 7472 33844
rect 3467 33813 3479 33816
rect 3421 33807 3479 33813
rect 7466 33804 7472 33816
rect 7524 33804 7530 33856
rect 7558 33804 7564 33856
rect 7616 33844 7622 33856
rect 10410 33844 10416 33856
rect 7616 33816 10416 33844
rect 7616 33804 7622 33816
rect 10410 33804 10416 33816
rect 10468 33804 10474 33856
rect 11146 33804 11152 33856
rect 11204 33844 11210 33856
rect 12820 33844 12848 33943
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 14918 33980 14924 33992
rect 14879 33952 14924 33980
rect 14918 33940 14924 33952
rect 14976 33940 14982 33992
rect 12897 33915 12955 33921
rect 12897 33881 12909 33915
rect 12943 33912 12955 33915
rect 14826 33912 14832 33924
rect 12943 33884 14832 33912
rect 12943 33881 12955 33884
rect 12897 33875 12955 33881
rect 14826 33872 14832 33884
rect 14884 33872 14890 33924
rect 11204 33816 12848 33844
rect 13633 33847 13691 33853
rect 11204 33804 11210 33816
rect 13633 33813 13645 33847
rect 13679 33844 13691 33847
rect 14182 33844 14188 33856
rect 13679 33816 14188 33844
rect 13679 33813 13691 33816
rect 13633 33807 13691 33813
rect 14182 33804 14188 33816
rect 14240 33804 14246 33856
rect 14274 33804 14280 33856
rect 14332 33844 14338 33856
rect 14332 33816 14377 33844
rect 14332 33804 14338 33816
rect 14550 33804 14556 33856
rect 14608 33844 14614 33856
rect 15013 33847 15071 33853
rect 15013 33844 15025 33847
rect 14608 33816 15025 33844
rect 14608 33804 14614 33816
rect 15013 33813 15025 33816
rect 15059 33813 15071 33847
rect 15013 33807 15071 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 3786 33600 3792 33652
rect 3844 33640 3850 33652
rect 6546 33640 6552 33652
rect 3844 33612 6552 33640
rect 3844 33600 3850 33612
rect 6546 33600 6552 33612
rect 6604 33640 6610 33652
rect 7742 33640 7748 33652
rect 6604 33612 7748 33640
rect 6604 33600 6610 33612
rect 7742 33600 7748 33612
rect 7800 33600 7806 33652
rect 9122 33640 9128 33652
rect 8680 33612 9128 33640
rect 8680 33584 8708 33612
rect 9122 33600 9128 33612
rect 9180 33600 9186 33652
rect 9306 33600 9312 33652
rect 9364 33640 9370 33652
rect 11793 33643 11851 33649
rect 9364 33612 11744 33640
rect 9364 33600 9370 33612
rect 1949 33575 2007 33581
rect 1949 33541 1961 33575
rect 1995 33572 2007 33575
rect 2038 33572 2044 33584
rect 1995 33544 2044 33572
rect 1995 33541 2007 33544
rect 1949 33535 2007 33541
rect 2038 33532 2044 33544
rect 2096 33532 2102 33584
rect 3602 33532 3608 33584
rect 3660 33572 3666 33584
rect 3697 33575 3755 33581
rect 3697 33572 3709 33575
rect 3660 33544 3709 33572
rect 3660 33532 3666 33544
rect 3697 33541 3709 33544
rect 3743 33541 3755 33575
rect 3697 33535 3755 33541
rect 8113 33575 8171 33581
rect 8113 33541 8125 33575
rect 8159 33572 8171 33575
rect 8662 33572 8668 33584
rect 8159 33544 8668 33572
rect 8159 33541 8171 33544
rect 8113 33535 8171 33541
rect 8662 33532 8668 33544
rect 8720 33532 8726 33584
rect 9030 33532 9036 33584
rect 9088 33572 9094 33584
rect 9088 33544 9614 33572
rect 9088 33532 9094 33544
rect 2590 33464 2596 33516
rect 2648 33464 2654 33516
rect 3970 33464 3976 33516
rect 4028 33504 4034 33516
rect 4028 33476 4073 33504
rect 4028 33464 4034 33476
rect 4430 33464 4436 33516
rect 4488 33504 4494 33516
rect 4893 33507 4951 33513
rect 4893 33504 4905 33507
rect 4488 33476 4905 33504
rect 4488 33464 4494 33476
rect 4893 33473 4905 33476
rect 4939 33504 4951 33507
rect 5813 33507 5871 33513
rect 5813 33504 5825 33507
rect 4939 33476 5825 33504
rect 4939 33473 4951 33476
rect 4893 33467 4951 33473
rect 5813 33473 5825 33476
rect 5859 33504 5871 33507
rect 6822 33504 6828 33516
rect 5859 33476 6828 33504
rect 5859 33473 5871 33476
rect 5813 33467 5871 33473
rect 6822 33464 6828 33476
rect 6880 33464 6886 33516
rect 7006 33464 7012 33516
rect 7064 33464 7070 33516
rect 8386 33464 8392 33516
rect 8444 33504 8450 33516
rect 8846 33504 8852 33516
rect 8444 33476 8852 33504
rect 8444 33464 8450 33476
rect 8846 33464 8852 33476
rect 8904 33464 8910 33516
rect 10410 33464 10416 33516
rect 10468 33504 10474 33516
rect 11716 33513 11744 33612
rect 11793 33609 11805 33643
rect 11839 33640 11851 33643
rect 11974 33640 11980 33652
rect 11839 33612 11980 33640
rect 11839 33609 11851 33612
rect 11793 33603 11851 33609
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 12342 33600 12348 33652
rect 12400 33640 12406 33652
rect 12400 33612 14780 33640
rect 12400 33600 12406 33612
rect 14182 33572 14188 33584
rect 14143 33544 14188 33572
rect 14182 33532 14188 33544
rect 14240 33532 14246 33584
rect 14752 33581 14780 33612
rect 14737 33575 14795 33581
rect 14737 33541 14749 33575
rect 14783 33541 14795 33575
rect 14737 33535 14795 33541
rect 11701 33507 11759 33513
rect 10468 33476 11192 33504
rect 10468 33464 10474 33476
rect 2314 33396 2320 33448
rect 2372 33436 2378 33448
rect 3142 33436 3148 33448
rect 2372 33408 3148 33436
rect 2372 33396 2378 33408
rect 3142 33396 3148 33408
rect 3200 33396 3206 33448
rect 4706 33436 4712 33448
rect 4667 33408 4712 33436
rect 4706 33396 4712 33408
rect 4764 33396 4770 33448
rect 5626 33436 5632 33448
rect 5587 33408 5632 33436
rect 5626 33396 5632 33408
rect 5684 33396 5690 33448
rect 7466 33396 7472 33448
rect 7524 33436 7530 33448
rect 9125 33439 9183 33445
rect 9125 33436 9137 33439
rect 7524 33408 9137 33436
rect 7524 33396 7530 33408
rect 9125 33405 9137 33408
rect 9171 33436 9183 33439
rect 9214 33436 9220 33448
rect 9171 33408 9220 33436
rect 9171 33405 9183 33408
rect 9125 33399 9183 33405
rect 9214 33396 9220 33408
rect 9272 33396 9278 33448
rect 9582 33396 9588 33448
rect 9640 33436 9646 33448
rect 11057 33439 11115 33445
rect 11057 33436 11069 33439
rect 9640 33408 11069 33436
rect 9640 33396 9646 33408
rect 11057 33405 11069 33408
rect 11103 33405 11115 33439
rect 11164 33436 11192 33476
rect 11701 33473 11713 33507
rect 11747 33473 11759 33507
rect 11701 33467 11759 33473
rect 11974 33464 11980 33516
rect 12032 33504 12038 33516
rect 12437 33507 12495 33513
rect 12437 33504 12449 33507
rect 12032 33476 12449 33504
rect 12032 33464 12038 33476
rect 12437 33473 12449 33476
rect 12483 33504 12495 33507
rect 13906 33504 13912 33516
rect 12483 33476 13912 33504
rect 12483 33473 12495 33476
rect 12437 33467 12495 33473
rect 13906 33464 13912 33476
rect 13964 33464 13970 33516
rect 14093 33439 14151 33445
rect 11164 33408 13860 33436
rect 11057 33399 11115 33405
rect 13832 33380 13860 33408
rect 14093 33405 14105 33439
rect 14139 33436 14151 33439
rect 14274 33436 14280 33448
rect 14139 33408 14280 33436
rect 14139 33405 14151 33408
rect 14093 33399 14151 33405
rect 14274 33396 14280 33408
rect 14332 33396 14338 33448
rect 11974 33368 11980 33380
rect 10152 33340 11980 33368
rect 2038 33260 2044 33312
rect 2096 33300 2102 33312
rect 5534 33300 5540 33312
rect 2096 33272 5540 33300
rect 2096 33260 2102 33272
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 6914 33300 6920 33312
rect 6687 33272 6920 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 6914 33260 6920 33272
rect 6972 33300 6978 33312
rect 7650 33300 7656 33312
rect 6972 33272 7656 33300
rect 6972 33260 6978 33272
rect 7650 33260 7656 33272
rect 7708 33260 7714 33312
rect 7742 33260 7748 33312
rect 7800 33300 7806 33312
rect 10152 33300 10180 33340
rect 11974 33328 11980 33340
rect 12032 33328 12038 33380
rect 13814 33328 13820 33380
rect 13872 33368 13878 33380
rect 14918 33368 14924 33380
rect 13872 33340 14924 33368
rect 13872 33328 13878 33340
rect 14918 33328 14924 33340
rect 14976 33328 14982 33380
rect 7800 33272 10180 33300
rect 7800 33260 7806 33272
rect 10226 33260 10232 33312
rect 10284 33300 10290 33312
rect 10597 33303 10655 33309
rect 10597 33300 10609 33303
rect 10284 33272 10609 33300
rect 10284 33260 10290 33272
rect 10597 33269 10609 33272
rect 10643 33269 10655 33303
rect 10597 33263 10655 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 4062 33096 4068 33108
rect 4023 33068 4068 33096
rect 4062 33056 4068 33068
rect 4120 33056 4126 33108
rect 8570 33096 8576 33108
rect 5552 33068 8576 33096
rect 5552 33028 5580 33068
rect 8570 33056 8576 33068
rect 8628 33056 8634 33108
rect 8846 33056 8852 33108
rect 8904 33096 8910 33108
rect 9125 33099 9183 33105
rect 9125 33096 9137 33099
rect 8904 33068 9137 33096
rect 8904 33056 8910 33068
rect 9125 33065 9137 33068
rect 9171 33096 9183 33099
rect 9582 33096 9588 33108
rect 9171 33068 9588 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 9582 33056 9588 33068
rect 9640 33096 9646 33108
rect 9677 33099 9735 33105
rect 9677 33096 9689 33099
rect 9640 33068 9689 33096
rect 9640 33056 9646 33068
rect 9677 33065 9689 33068
rect 9723 33065 9735 33099
rect 10870 33096 10876 33108
rect 10831 33068 10876 33096
rect 9677 33059 9735 33065
rect 10870 33056 10876 33068
rect 10928 33056 10934 33108
rect 11425 33099 11483 33105
rect 11425 33065 11437 33099
rect 11471 33096 11483 33099
rect 11790 33096 11796 33108
rect 11471 33068 11796 33096
rect 11471 33065 11483 33068
rect 11425 33059 11483 33065
rect 11790 33056 11796 33068
rect 11848 33056 11854 33108
rect 3344 33000 5580 33028
rect 3145 32963 3203 32969
rect 3145 32929 3157 32963
rect 3191 32960 3203 32963
rect 3344 32960 3372 33000
rect 6914 32988 6920 33040
rect 6972 33028 6978 33040
rect 7742 33028 7748 33040
rect 6972 33000 7748 33028
rect 6972 32988 6978 33000
rect 7742 32988 7748 33000
rect 7800 33028 7806 33040
rect 10888 33028 10916 33056
rect 7800 33000 10916 33028
rect 7800 32988 7806 33000
rect 3191 32932 3372 32960
rect 3421 32963 3479 32969
rect 3191 32929 3203 32932
rect 3145 32923 3203 32929
rect 3421 32929 3433 32963
rect 3467 32960 3479 32963
rect 3878 32960 3884 32972
rect 3467 32932 3884 32960
rect 3467 32929 3479 32932
rect 3421 32923 3479 32929
rect 3878 32920 3884 32932
rect 3936 32920 3942 32972
rect 4801 32963 4859 32969
rect 4801 32929 4813 32963
rect 4847 32960 4859 32963
rect 5166 32960 5172 32972
rect 4847 32932 5172 32960
rect 4847 32929 4859 32932
rect 4801 32923 4859 32929
rect 5166 32920 5172 32932
rect 5224 32920 5230 32972
rect 10134 32960 10140 32972
rect 5368 32932 10140 32960
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32892 4307 32895
rect 4614 32892 4620 32904
rect 4295 32864 4620 32892
rect 4295 32861 4307 32864
rect 4249 32855 4307 32861
rect 4614 32852 4620 32864
rect 4672 32852 4678 32904
rect 5368 32892 5396 32932
rect 10134 32920 10140 32932
rect 10192 32960 10198 32972
rect 10318 32960 10324 32972
rect 10192 32932 10324 32960
rect 10192 32920 10198 32932
rect 10318 32920 10324 32932
rect 10376 32920 10382 32972
rect 5092 32864 5396 32892
rect 2714 32796 2774 32824
rect 1673 32759 1731 32765
rect 1673 32725 1685 32759
rect 1719 32756 1731 32759
rect 1854 32756 1860 32768
rect 1719 32728 1860 32756
rect 1719 32725 1731 32728
rect 1673 32719 1731 32725
rect 1854 32716 1860 32728
rect 1912 32716 1918 32768
rect 2746 32756 2774 32796
rect 4338 32784 4344 32836
rect 4396 32824 4402 32836
rect 5092 32824 5120 32864
rect 6822 32852 6828 32904
rect 6880 32892 6886 32904
rect 7285 32895 7343 32901
rect 7285 32892 7297 32895
rect 6880 32864 7297 32892
rect 6880 32852 6886 32864
rect 7285 32861 7297 32864
rect 7331 32892 7343 32895
rect 7837 32895 7895 32901
rect 7837 32892 7849 32895
rect 7331 32864 7849 32892
rect 7331 32861 7343 32864
rect 7285 32855 7343 32861
rect 7837 32861 7849 32864
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 11054 32852 11060 32904
rect 11112 32892 11118 32904
rect 11333 32895 11391 32901
rect 11333 32892 11345 32895
rect 11112 32864 11345 32892
rect 11112 32852 11118 32864
rect 11333 32861 11345 32864
rect 11379 32861 11391 32895
rect 11333 32855 11391 32861
rect 4396 32796 5120 32824
rect 4396 32784 4402 32796
rect 5166 32784 5172 32836
rect 5224 32824 5230 32836
rect 6549 32827 6607 32833
rect 5224 32796 5382 32824
rect 5224 32784 5230 32796
rect 6549 32793 6561 32827
rect 6595 32824 6607 32827
rect 8389 32827 8447 32833
rect 8389 32824 8401 32827
rect 6595 32796 8401 32824
rect 6595 32793 6607 32796
rect 6549 32787 6607 32793
rect 8389 32793 8401 32796
rect 8435 32824 8447 32827
rect 8754 32824 8760 32836
rect 8435 32796 8760 32824
rect 8435 32793 8447 32796
rect 8389 32787 8447 32793
rect 8754 32784 8760 32796
rect 8812 32784 8818 32836
rect 38013 32827 38071 32833
rect 38013 32824 38025 32827
rect 10244 32796 12434 32824
rect 3234 32756 3240 32768
rect 2746 32728 3240 32756
rect 3234 32716 3240 32728
rect 3292 32716 3298 32768
rect 3602 32716 3608 32768
rect 3660 32756 3666 32768
rect 10244 32765 10272 32796
rect 10229 32759 10287 32765
rect 10229 32756 10241 32759
rect 3660 32728 10241 32756
rect 3660 32716 3666 32728
rect 10229 32725 10241 32728
rect 10275 32725 10287 32759
rect 12406 32756 12434 32796
rect 26206 32796 38025 32824
rect 12526 32756 12532 32768
rect 12406 32728 12532 32756
rect 10229 32719 10287 32725
rect 12526 32716 12532 32728
rect 12584 32716 12590 32768
rect 23106 32716 23112 32768
rect 23164 32756 23170 32768
rect 26206 32756 26234 32796
rect 38013 32793 38025 32796
rect 38059 32793 38071 32827
rect 38194 32824 38200 32836
rect 38155 32796 38200 32824
rect 38013 32787 38071 32793
rect 38194 32784 38200 32796
rect 38252 32784 38258 32836
rect 23164 32728 26234 32756
rect 37553 32759 37611 32765
rect 23164 32716 23170 32728
rect 37553 32725 37565 32759
rect 37599 32756 37611 32759
rect 38212 32756 38240 32784
rect 37599 32728 38240 32756
rect 37599 32725 37611 32728
rect 37553 32719 37611 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 3878 32512 3884 32564
rect 3936 32552 3942 32564
rect 3936 32524 5028 32552
rect 3936 32512 3942 32524
rect 2866 32444 2872 32496
rect 2924 32484 2930 32496
rect 2924 32456 3542 32484
rect 2924 32444 2930 32456
rect 4614 32444 4620 32496
rect 4672 32484 4678 32496
rect 4798 32484 4804 32496
rect 4672 32456 4804 32484
rect 4672 32444 4678 32456
rect 4798 32444 4804 32456
rect 4856 32444 4862 32496
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 2774 32416 2780 32428
rect 1627 32388 2780 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 2774 32376 2780 32388
rect 2832 32376 2838 32428
rect 5000 32425 5028 32524
rect 5902 32512 5908 32564
rect 5960 32552 5966 32564
rect 7101 32555 7159 32561
rect 7101 32552 7113 32555
rect 5960 32524 7113 32552
rect 5960 32512 5966 32524
rect 7101 32521 7113 32524
rect 7147 32552 7159 32555
rect 7147 32524 12434 32552
rect 7147 32521 7159 32524
rect 7101 32515 7159 32521
rect 6730 32484 6736 32496
rect 5092 32456 6736 32484
rect 4985 32419 5043 32425
rect 4985 32385 4997 32419
rect 5031 32385 5043 32419
rect 4985 32379 5043 32385
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32348 1915 32351
rect 2406 32348 2412 32360
rect 1903 32320 2412 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 2406 32308 2412 32320
rect 2464 32308 2470 32360
rect 2961 32351 3019 32357
rect 2961 32317 2973 32351
rect 3007 32348 3019 32351
rect 4338 32348 4344 32360
rect 3007 32320 4344 32348
rect 3007 32317 3019 32320
rect 2961 32311 3019 32317
rect 4338 32308 4344 32320
rect 4396 32308 4402 32360
rect 4709 32351 4767 32357
rect 4709 32317 4721 32351
rect 4755 32348 4767 32351
rect 5092 32348 5120 32456
rect 6730 32444 6736 32456
rect 6788 32444 6794 32496
rect 7190 32444 7196 32496
rect 7248 32484 7254 32496
rect 12406 32484 12434 32524
rect 14458 32484 14464 32496
rect 7248 32456 7406 32484
rect 12406 32456 14464 32484
rect 7248 32444 7254 32456
rect 14458 32444 14464 32456
rect 14516 32444 14522 32496
rect 15010 32484 15016 32496
rect 14971 32456 15016 32484
rect 15010 32444 15016 32456
rect 15068 32444 15074 32496
rect 15933 32487 15991 32493
rect 15933 32453 15945 32487
rect 15979 32484 15991 32487
rect 16022 32484 16028 32496
rect 15979 32456 16028 32484
rect 15979 32453 15991 32456
rect 15933 32447 15991 32453
rect 16022 32444 16028 32456
rect 16080 32444 16086 32496
rect 5258 32376 5264 32428
rect 5316 32416 5322 32428
rect 5626 32416 5632 32428
rect 5316 32388 5632 32416
rect 5316 32376 5322 32388
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 8846 32376 8852 32428
rect 8904 32416 8910 32428
rect 9309 32419 9367 32425
rect 9309 32416 9321 32419
rect 8904 32388 9321 32416
rect 8904 32376 8910 32388
rect 9309 32385 9321 32388
rect 9355 32416 9367 32419
rect 9861 32419 9919 32425
rect 9861 32416 9873 32419
rect 9355 32388 9873 32416
rect 9355 32385 9367 32388
rect 9309 32379 9367 32385
rect 9861 32385 9873 32388
rect 9907 32416 9919 32419
rect 10413 32419 10471 32425
rect 10413 32416 10425 32419
rect 9907 32388 10425 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 10413 32385 10425 32388
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 12529 32419 12587 32425
rect 12529 32385 12541 32419
rect 12575 32385 12587 32419
rect 13170 32416 13176 32428
rect 13131 32388 13176 32416
rect 12529 32379 12587 32385
rect 8570 32348 8576 32360
rect 4755 32320 5120 32348
rect 8531 32320 8576 32348
rect 4755 32317 4767 32320
rect 4709 32311 4767 32317
rect 8570 32308 8576 32320
rect 8628 32308 8634 32360
rect 5537 32215 5595 32221
rect 5537 32181 5549 32215
rect 5583 32212 5595 32215
rect 5626 32212 5632 32224
rect 5583 32184 5632 32212
rect 5583 32181 5595 32184
rect 5537 32175 5595 32181
rect 5626 32172 5632 32184
rect 5684 32172 5690 32224
rect 6730 32172 6736 32224
rect 6788 32212 6794 32224
rect 12544 32212 12572 32379
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32348 14979 32351
rect 15562 32348 15568 32360
rect 14967 32320 15568 32348
rect 14967 32317 14979 32320
rect 14921 32311 14979 32317
rect 15562 32308 15568 32320
rect 15620 32308 15626 32360
rect 12621 32283 12679 32289
rect 12621 32249 12633 32283
rect 12667 32280 12679 32283
rect 15930 32280 15936 32292
rect 12667 32252 15936 32280
rect 12667 32249 12679 32252
rect 12621 32243 12679 32249
rect 15930 32240 15936 32252
rect 15988 32240 15994 32292
rect 6788 32184 12572 32212
rect 13265 32215 13323 32221
rect 6788 32172 6794 32184
rect 13265 32181 13277 32215
rect 13311 32212 13323 32215
rect 16206 32212 16212 32224
rect 13311 32184 16212 32212
rect 13311 32181 13323 32184
rect 13265 32175 13323 32181
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 6365 32011 6423 32017
rect 6365 31977 6377 32011
rect 6411 32008 6423 32011
rect 8202 32008 8208 32020
rect 6411 31980 8208 32008
rect 6411 31977 6423 31980
rect 6365 31971 6423 31977
rect 8202 31968 8208 31980
rect 8260 31968 8266 32020
rect 8846 31968 8852 32020
rect 8904 32008 8910 32020
rect 9125 32011 9183 32017
rect 9125 32008 9137 32011
rect 8904 31980 9137 32008
rect 8904 31968 8910 31980
rect 9125 31977 9137 31980
rect 9171 32008 9183 32011
rect 9306 32008 9312 32020
rect 9171 31980 9312 32008
rect 9171 31977 9183 31980
rect 9125 31971 9183 31977
rect 9306 31968 9312 31980
rect 9364 32008 9370 32020
rect 9677 32011 9735 32017
rect 9677 32008 9689 32011
rect 9364 31980 9689 32008
rect 9364 31968 9370 31980
rect 9677 31977 9689 31980
rect 9723 31977 9735 32011
rect 9677 31971 9735 31977
rect 6270 31900 6276 31952
rect 6328 31940 6334 31952
rect 6638 31940 6644 31952
rect 6328 31912 6644 31940
rect 6328 31900 6334 31912
rect 6638 31900 6644 31912
rect 6696 31900 6702 31952
rect 1946 31872 1952 31884
rect 1907 31844 1952 31872
rect 1946 31832 1952 31844
rect 2004 31832 2010 31884
rect 3418 31872 3424 31884
rect 3379 31844 3424 31872
rect 3418 31832 3424 31844
rect 3476 31832 3482 31884
rect 4154 31832 4160 31884
rect 4212 31872 4218 31884
rect 4617 31875 4675 31881
rect 4617 31872 4629 31875
rect 4212 31844 4629 31872
rect 4212 31832 4218 31844
rect 4617 31841 4629 31844
rect 4663 31872 4675 31875
rect 4663 31844 6500 31872
rect 4663 31841 4675 31844
rect 4617 31835 4675 31841
rect 1670 31804 1676 31816
rect 1631 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 3973 31807 4031 31813
rect 3973 31773 3985 31807
rect 4019 31804 4031 31807
rect 6270 31804 6276 31816
rect 4019 31776 4292 31804
rect 6026 31776 6276 31804
rect 4019 31773 4031 31776
rect 3973 31767 4031 31773
rect 3602 31736 3608 31748
rect 3174 31708 3608 31736
rect 3602 31696 3608 31708
rect 3660 31696 3666 31748
rect 4065 31671 4123 31677
rect 4065 31637 4077 31671
rect 4111 31668 4123 31671
rect 4154 31668 4160 31680
rect 4111 31640 4160 31668
rect 4111 31637 4123 31640
rect 4065 31631 4123 31637
rect 4154 31628 4160 31640
rect 4212 31628 4218 31680
rect 4264 31668 4292 31776
rect 6270 31764 6276 31776
rect 6328 31764 6334 31816
rect 6472 31804 6500 31844
rect 6546 31832 6552 31884
rect 6604 31872 6610 31884
rect 7101 31875 7159 31881
rect 7101 31872 7113 31875
rect 6604 31844 7113 31872
rect 6604 31832 6610 31844
rect 7101 31841 7113 31844
rect 7147 31872 7159 31875
rect 8570 31872 8576 31884
rect 7147 31844 8340 31872
rect 8483 31844 8576 31872
rect 7147 31841 7159 31844
rect 7101 31835 7159 31841
rect 6822 31804 6828 31816
rect 6472 31776 6828 31804
rect 6822 31764 6828 31776
rect 6880 31764 6886 31816
rect 8312 31804 8340 31844
rect 8570 31832 8576 31844
rect 8628 31872 8634 31884
rect 12250 31872 12256 31884
rect 8628 31844 12256 31872
rect 8628 31832 8634 31844
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 12894 31804 12900 31816
rect 8312 31776 12900 31804
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 15746 31764 15752 31816
rect 15804 31804 15810 31816
rect 18509 31807 18567 31813
rect 18509 31804 18521 31807
rect 15804 31776 18521 31804
rect 15804 31764 15810 31776
rect 18509 31773 18521 31776
rect 18555 31773 18567 31807
rect 18509 31767 18567 31773
rect 18601 31807 18659 31813
rect 18601 31773 18613 31807
rect 18647 31804 18659 31807
rect 19429 31807 19487 31813
rect 19429 31804 19441 31807
rect 18647 31776 19441 31804
rect 18647 31773 18659 31776
rect 18601 31767 18659 31773
rect 19429 31773 19441 31776
rect 19475 31804 19487 31807
rect 23106 31804 23112 31816
rect 19475 31776 23112 31804
rect 19475 31773 19487 31776
rect 19429 31767 19487 31773
rect 23106 31764 23112 31776
rect 23164 31764 23170 31816
rect 4893 31739 4951 31745
rect 4893 31705 4905 31739
rect 4939 31736 4951 31739
rect 4939 31708 5304 31736
rect 4939 31705 4951 31708
rect 4893 31699 4951 31705
rect 5166 31668 5172 31680
rect 4264 31640 5172 31668
rect 5166 31628 5172 31640
rect 5224 31628 5230 31680
rect 5276 31668 5304 31708
rect 6362 31696 6368 31748
rect 6420 31736 6426 31748
rect 6420 31708 7590 31736
rect 6420 31696 6426 31708
rect 5902 31668 5908 31680
rect 5276 31640 5908 31668
rect 5902 31628 5908 31640
rect 5960 31628 5966 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1670 31424 1676 31476
rect 1728 31464 1734 31476
rect 3878 31464 3884 31476
rect 1728 31436 3884 31464
rect 1728 31424 1734 31436
rect 1780 31337 1808 31436
rect 3878 31424 3884 31436
rect 3936 31464 3942 31476
rect 3936 31436 4016 31464
rect 3936 31424 3942 31436
rect 3786 31396 3792 31408
rect 3266 31368 3792 31396
rect 3786 31356 3792 31368
rect 3844 31356 3850 31408
rect 3988 31337 4016 31436
rect 4154 31424 4160 31476
rect 4212 31464 4218 31476
rect 6549 31467 6607 31473
rect 4212 31436 5580 31464
rect 4212 31424 4218 31436
rect 5552 31396 5580 31436
rect 6549 31433 6561 31467
rect 6595 31464 6607 31467
rect 6730 31464 6736 31476
rect 6595 31436 6736 31464
rect 6595 31433 6607 31436
rect 6549 31427 6607 31433
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 7282 31424 7288 31476
rect 7340 31464 7346 31476
rect 7340 31436 12434 31464
rect 7340 31424 7346 31436
rect 8018 31396 8024 31408
rect 5552 31368 6854 31396
rect 7931 31368 8024 31396
rect 8018 31356 8024 31368
rect 8076 31396 8082 31408
rect 11146 31396 11152 31408
rect 8076 31368 11152 31396
rect 8076 31356 8082 31368
rect 11146 31356 11152 31368
rect 11204 31356 11210 31408
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31297 1823 31331
rect 1765 31291 1823 31297
rect 3973 31331 4031 31337
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 5626 31328 5632 31340
rect 5382 31300 5632 31328
rect 3973 31291 4031 31297
rect 5626 31288 5632 31300
rect 5684 31288 5690 31340
rect 5994 31288 6000 31340
rect 6052 31328 6058 31340
rect 6730 31328 6736 31340
rect 6052 31300 6736 31328
rect 6052 31288 6058 31300
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 8754 31328 8760 31340
rect 8715 31300 8760 31328
rect 8754 31288 8760 31300
rect 8812 31288 8818 31340
rect 1486 31220 1492 31272
rect 1544 31260 1550 31272
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1544 31232 2053 31260
rect 1544 31220 1550 31232
rect 2041 31229 2053 31232
rect 2087 31260 2099 31263
rect 4249 31263 4307 31269
rect 2087 31232 4108 31260
rect 2087 31229 2099 31232
rect 2041 31223 2099 31229
rect 3513 31127 3571 31133
rect 3513 31093 3525 31127
rect 3559 31124 3571 31127
rect 3694 31124 3700 31136
rect 3559 31096 3700 31124
rect 3559 31093 3571 31096
rect 3513 31087 3571 31093
rect 3694 31084 3700 31096
rect 3752 31124 3758 31136
rect 3878 31124 3884 31136
rect 3752 31096 3884 31124
rect 3752 31084 3758 31096
rect 3878 31084 3884 31096
rect 3936 31084 3942 31136
rect 4080 31124 4108 31232
rect 4249 31229 4261 31263
rect 4295 31260 4307 31263
rect 4614 31260 4620 31272
rect 4295 31232 4620 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 4614 31220 4620 31232
rect 4672 31220 4678 31272
rect 5258 31220 5264 31272
rect 5316 31260 5322 31272
rect 8297 31263 8355 31269
rect 5316 31232 8248 31260
rect 5316 31220 5322 31232
rect 6914 31192 6920 31204
rect 5276 31164 6920 31192
rect 5276 31124 5304 31164
rect 6914 31152 6920 31164
rect 6972 31152 6978 31204
rect 8220 31192 8248 31232
rect 8297 31229 8309 31263
rect 8343 31260 8355 31263
rect 9306 31260 9312 31272
rect 8343 31232 9312 31260
rect 8343 31229 8355 31232
rect 8297 31223 8355 31229
rect 9306 31220 9312 31232
rect 9364 31260 9370 31272
rect 9401 31263 9459 31269
rect 9401 31260 9413 31263
rect 9364 31232 9413 31260
rect 9364 31220 9370 31232
rect 9401 31229 9413 31232
rect 9447 31260 9459 31263
rect 9953 31263 10011 31269
rect 9953 31260 9965 31263
rect 9447 31232 9965 31260
rect 9447 31229 9459 31232
rect 9401 31223 9459 31229
rect 9953 31229 9965 31232
rect 9999 31229 10011 31263
rect 9953 31223 10011 31229
rect 8938 31192 8944 31204
rect 8220 31164 8944 31192
rect 8938 31152 8944 31164
rect 8996 31152 9002 31204
rect 12406 31192 12434 31436
rect 15102 31356 15108 31408
rect 15160 31396 15166 31408
rect 16117 31399 16175 31405
rect 16117 31396 16129 31399
rect 15160 31368 16129 31396
rect 15160 31356 15166 31368
rect 16117 31365 16129 31368
rect 16163 31365 16175 31399
rect 16117 31359 16175 31365
rect 14737 31331 14795 31337
rect 14737 31297 14749 31331
rect 14783 31297 14795 31331
rect 20438 31328 20444 31340
rect 20399 31300 20444 31328
rect 14737 31291 14795 31297
rect 14093 31195 14151 31201
rect 14093 31192 14105 31195
rect 12406 31164 14105 31192
rect 14093 31161 14105 31164
rect 14139 31192 14151 31195
rect 14752 31192 14780 31291
rect 20438 31288 20444 31300
rect 20496 31328 20502 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 20496 31300 21097 31328
rect 20496 31288 20502 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 15378 31260 15384 31272
rect 15339 31232 15384 31260
rect 15378 31220 15384 31232
rect 15436 31260 15442 31272
rect 16022 31260 16028 31272
rect 15436 31232 16028 31260
rect 15436 31220 15442 31232
rect 16022 31220 16028 31232
rect 16080 31220 16086 31272
rect 16209 31263 16267 31269
rect 16209 31229 16221 31263
rect 16255 31260 16267 31263
rect 18046 31260 18052 31272
rect 16255 31232 18052 31260
rect 16255 31229 16267 31232
rect 16209 31223 16267 31229
rect 18046 31220 18052 31232
rect 18104 31220 18110 31272
rect 17954 31192 17960 31204
rect 14139 31164 17960 31192
rect 14139 31161 14151 31164
rect 14093 31155 14151 31161
rect 17954 31152 17960 31164
rect 18012 31152 18018 31204
rect 20625 31195 20683 31201
rect 20625 31161 20637 31195
rect 20671 31192 20683 31195
rect 20671 31164 26234 31192
rect 20671 31161 20683 31164
rect 20625 31155 20683 31161
rect 5718 31124 5724 31136
rect 4080 31096 5304 31124
rect 5679 31096 5724 31124
rect 5718 31084 5724 31096
rect 5776 31084 5782 31136
rect 6178 31084 6184 31136
rect 6236 31124 6242 31136
rect 8754 31124 8760 31136
rect 6236 31096 8760 31124
rect 6236 31084 6242 31096
rect 8754 31084 8760 31096
rect 8812 31084 8818 31136
rect 8849 31127 8907 31133
rect 8849 31093 8861 31127
rect 8895 31124 8907 31127
rect 9674 31124 9680 31136
rect 8895 31096 9680 31124
rect 8895 31093 8907 31096
rect 8849 31087 8907 31093
rect 9674 31084 9680 31096
rect 9732 31084 9738 31136
rect 14642 31124 14648 31136
rect 14603 31096 14648 31124
rect 14642 31084 14648 31096
rect 14700 31084 14706 31136
rect 26206 31124 26234 31164
rect 38010 31124 38016 31136
rect 26206 31096 38016 31124
rect 38010 31084 38016 31096
rect 38068 31084 38074 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1857 30923 1915 30929
rect 1857 30889 1869 30923
rect 1903 30920 1915 30923
rect 2038 30920 2044 30932
rect 1903 30892 2044 30920
rect 1903 30889 1915 30892
rect 1857 30883 1915 30889
rect 2038 30880 2044 30892
rect 2096 30880 2102 30932
rect 2501 30923 2559 30929
rect 2501 30889 2513 30923
rect 2547 30920 2559 30923
rect 2958 30920 2964 30932
rect 2547 30892 2964 30920
rect 2547 30889 2559 30892
rect 2501 30883 2559 30889
rect 2958 30880 2964 30892
rect 3016 30880 3022 30932
rect 3142 30920 3148 30932
rect 3103 30892 3148 30920
rect 3142 30880 3148 30892
rect 3200 30880 3206 30932
rect 4709 30923 4767 30929
rect 3988 30892 4652 30920
rect 1964 30756 3464 30784
rect 1964 30725 1992 30756
rect 3436 30728 3464 30756
rect 1949 30719 2007 30725
rect 1949 30685 1961 30719
rect 1995 30685 2007 30719
rect 1949 30679 2007 30685
rect 2409 30719 2467 30725
rect 2409 30685 2421 30719
rect 2455 30716 2467 30719
rect 3234 30716 3240 30728
rect 2455 30688 3240 30716
rect 2455 30685 2467 30688
rect 2409 30679 2467 30685
rect 3234 30676 3240 30688
rect 3292 30676 3298 30728
rect 3418 30676 3424 30728
rect 3476 30716 3482 30728
rect 3988 30725 4016 30892
rect 4522 30812 4528 30864
rect 4580 30812 4586 30864
rect 4624 30852 4652 30892
rect 4709 30889 4721 30923
rect 4755 30920 4767 30923
rect 5626 30920 5632 30932
rect 4755 30892 5632 30920
rect 4755 30889 4767 30892
rect 4709 30883 4767 30889
rect 5626 30880 5632 30892
rect 5684 30880 5690 30932
rect 5718 30880 5724 30932
rect 5776 30920 5782 30932
rect 6168 30923 6226 30929
rect 6168 30920 6180 30923
rect 5776 30892 6180 30920
rect 5776 30880 5782 30892
rect 6168 30889 6180 30892
rect 6214 30920 6226 30923
rect 13170 30920 13176 30932
rect 6214 30892 13176 30920
rect 6214 30889 6226 30892
rect 6168 30883 6226 30889
rect 13170 30880 13176 30892
rect 13228 30880 13234 30932
rect 16022 30880 16028 30932
rect 16080 30920 16086 30932
rect 16298 30920 16304 30932
rect 16080 30892 16304 30920
rect 16080 30880 16086 30892
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 16850 30920 16856 30932
rect 16811 30892 16856 30920
rect 16850 30880 16856 30892
rect 16908 30880 16914 30932
rect 37550 30920 37556 30932
rect 37511 30892 37556 30920
rect 37550 30880 37556 30892
rect 37608 30880 37614 30932
rect 5166 30852 5172 30864
rect 4624 30824 5172 30852
rect 5166 30812 5172 30824
rect 5224 30812 5230 30864
rect 5258 30812 5264 30864
rect 5316 30852 5322 30864
rect 5353 30855 5411 30861
rect 5353 30852 5365 30855
rect 5316 30824 5365 30852
rect 5316 30812 5322 30824
rect 5353 30821 5365 30824
rect 5399 30821 5411 30855
rect 5353 30815 5411 30821
rect 7653 30855 7711 30861
rect 7653 30821 7665 30855
rect 7699 30852 7711 30855
rect 8018 30852 8024 30864
rect 7699 30824 8024 30852
rect 7699 30821 7711 30824
rect 7653 30815 7711 30821
rect 8018 30812 8024 30824
rect 8076 30812 8082 30864
rect 20438 30852 20444 30864
rect 11532 30824 20444 30852
rect 4540 30726 4568 30812
rect 5905 30787 5963 30793
rect 5905 30753 5917 30787
rect 5951 30784 5963 30787
rect 6638 30784 6644 30796
rect 5951 30756 6644 30784
rect 5951 30753 5963 30756
rect 5905 30747 5963 30753
rect 6638 30744 6644 30756
rect 6696 30784 6702 30796
rect 6822 30784 6828 30796
rect 6696 30756 6828 30784
rect 6696 30744 6702 30756
rect 6822 30744 6828 30756
rect 6880 30744 6886 30796
rect 6914 30744 6920 30796
rect 6972 30784 6978 30796
rect 6972 30756 9168 30784
rect 6972 30744 6978 30756
rect 4609 30729 4667 30735
rect 4609 30726 4621 30729
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 3476 30688 3985 30716
rect 3476 30676 3482 30688
rect 3973 30685 3985 30688
rect 4019 30685 4031 30719
rect 4540 30698 4621 30726
rect 4609 30695 4621 30698
rect 4655 30695 4667 30729
rect 4609 30689 4667 30695
rect 3973 30679 4031 30685
rect 5166 30676 5172 30728
rect 5224 30716 5230 30728
rect 5261 30719 5319 30725
rect 5261 30716 5273 30719
rect 5224 30688 5273 30716
rect 5224 30676 5230 30688
rect 5261 30685 5273 30688
rect 5307 30716 5319 30719
rect 5718 30716 5724 30728
rect 5307 30688 5724 30716
rect 5307 30685 5319 30688
rect 5261 30679 5319 30685
rect 5718 30676 5724 30688
rect 5776 30676 5782 30728
rect 8110 30716 8116 30728
rect 8071 30688 8116 30716
rect 8110 30676 8116 30688
rect 8168 30676 8174 30728
rect 9140 30725 9168 30756
rect 11532 30725 11560 30824
rect 20438 30812 20444 30824
rect 20496 30812 20502 30864
rect 11609 30787 11667 30793
rect 11609 30753 11621 30787
rect 11655 30784 11667 30787
rect 11974 30784 11980 30796
rect 11655 30756 11980 30784
rect 11655 30753 11667 30756
rect 11609 30747 11667 30753
rect 11974 30744 11980 30756
rect 12032 30784 12038 30796
rect 12253 30787 12311 30793
rect 12253 30784 12265 30787
rect 12032 30756 12265 30784
rect 12032 30744 12038 30756
rect 12253 30753 12265 30756
rect 12299 30753 12311 30787
rect 12253 30747 12311 30753
rect 12434 30744 12440 30796
rect 12492 30784 12498 30796
rect 12529 30787 12587 30793
rect 12529 30784 12541 30787
rect 12492 30756 12541 30784
rect 12492 30744 12498 30756
rect 12529 30753 12541 30756
rect 12575 30753 12587 30787
rect 14550 30784 14556 30796
rect 14511 30756 14556 30784
rect 12529 30747 12587 30753
rect 14550 30744 14556 30756
rect 14608 30744 14614 30796
rect 9125 30719 9183 30725
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 11517 30719 11575 30725
rect 11517 30716 11529 30719
rect 9125 30679 9183 30685
rect 11072 30688 11529 30716
rect 11072 30657 11100 30688
rect 11517 30685 11529 30688
rect 11563 30685 11575 30719
rect 11517 30679 11575 30685
rect 15841 30719 15899 30725
rect 15841 30685 15853 30719
rect 15887 30716 15899 30719
rect 16482 30716 16488 30728
rect 15887 30688 16488 30716
rect 15887 30685 15899 30688
rect 15841 30679 15899 30685
rect 16482 30676 16488 30688
rect 16540 30676 16546 30728
rect 37369 30719 37427 30725
rect 37369 30685 37381 30719
rect 37415 30685 37427 30719
rect 38010 30716 38016 30728
rect 37971 30688 38016 30716
rect 37369 30679 37427 30685
rect 4065 30651 4123 30657
rect 4065 30617 4077 30651
rect 4111 30648 4123 30651
rect 11057 30651 11115 30657
rect 11057 30648 11069 30651
rect 4111 30620 6670 30648
rect 8128 30620 11069 30648
rect 4111 30617 4123 30620
rect 4065 30611 4123 30617
rect 3234 30540 3240 30592
rect 3292 30580 3298 30592
rect 5074 30580 5080 30592
rect 3292 30552 5080 30580
rect 3292 30540 3298 30552
rect 5074 30540 5080 30552
rect 5132 30540 5138 30592
rect 6914 30540 6920 30592
rect 6972 30580 6978 30592
rect 8128 30580 8156 30620
rect 11057 30617 11069 30620
rect 11103 30617 11115 30651
rect 12342 30648 12348 30660
rect 12303 30620 12348 30648
rect 11057 30611 11115 30617
rect 12342 30608 12348 30620
rect 12400 30608 12406 30660
rect 14642 30608 14648 30660
rect 14700 30648 14706 30660
rect 15197 30651 15255 30657
rect 14700 30620 14745 30648
rect 14700 30608 14706 30620
rect 15197 30617 15209 30651
rect 15243 30648 15255 30651
rect 15286 30648 15292 30660
rect 15243 30620 15292 30648
rect 15243 30617 15255 30620
rect 15197 30611 15255 30617
rect 15286 30608 15292 30620
rect 15344 30608 15350 30660
rect 37384 30648 37412 30679
rect 38010 30676 38016 30688
rect 38068 30676 38074 30728
rect 38102 30648 38108 30660
rect 37384 30620 38108 30648
rect 38102 30608 38108 30620
rect 38160 30608 38166 30660
rect 6972 30552 8156 30580
rect 8205 30583 8263 30589
rect 6972 30540 6978 30552
rect 8205 30549 8217 30583
rect 8251 30580 8263 30583
rect 8294 30580 8300 30592
rect 8251 30552 8300 30580
rect 8251 30549 8263 30552
rect 8205 30543 8263 30549
rect 8294 30540 8300 30552
rect 8352 30540 8358 30592
rect 9217 30583 9275 30589
rect 9217 30549 9229 30583
rect 9263 30580 9275 30583
rect 9582 30580 9588 30592
rect 9263 30552 9588 30580
rect 9263 30549 9275 30552
rect 9217 30543 9275 30549
rect 9582 30540 9588 30552
rect 9640 30540 9646 30592
rect 15470 30540 15476 30592
rect 15528 30580 15534 30592
rect 15749 30583 15807 30589
rect 15749 30580 15761 30583
rect 15528 30552 15761 30580
rect 15528 30540 15534 30552
rect 15749 30549 15761 30552
rect 15795 30549 15807 30583
rect 38194 30580 38200 30592
rect 38155 30552 38200 30580
rect 15749 30543 15807 30549
rect 38194 30540 38200 30552
rect 38252 30540 38258 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1946 30336 1952 30388
rect 2004 30376 2010 30388
rect 8110 30376 8116 30388
rect 2004 30348 8116 30376
rect 2004 30336 2010 30348
rect 8110 30336 8116 30348
rect 8168 30336 8174 30388
rect 12342 30376 12348 30388
rect 12303 30348 12348 30376
rect 12342 30336 12348 30348
rect 12400 30336 12406 30388
rect 2409 30311 2467 30317
rect 2409 30277 2421 30311
rect 2455 30308 2467 30311
rect 3142 30308 3148 30320
rect 2455 30280 3148 30308
rect 2455 30277 2467 30280
rect 2409 30271 2467 30277
rect 3142 30268 3148 30280
rect 3200 30268 3206 30320
rect 3786 30268 3792 30320
rect 3844 30308 3850 30320
rect 4065 30311 4123 30317
rect 4065 30308 4077 30311
rect 3844 30280 4077 30308
rect 3844 30268 3850 30280
rect 4065 30277 4077 30280
rect 4111 30277 4123 30311
rect 5442 30308 5448 30320
rect 5403 30280 5448 30308
rect 4065 30271 4123 30277
rect 5442 30268 5448 30280
rect 5500 30268 5506 30320
rect 5810 30268 5816 30320
rect 5868 30308 5874 30320
rect 6641 30311 6699 30317
rect 6641 30308 6653 30311
rect 5868 30280 6653 30308
rect 5868 30268 5874 30280
rect 6641 30277 6653 30280
rect 6687 30277 6699 30311
rect 6641 30271 6699 30277
rect 6730 30268 6736 30320
rect 6788 30308 6794 30320
rect 7193 30311 7251 30317
rect 7193 30308 7205 30311
rect 6788 30280 7205 30308
rect 6788 30268 6794 30280
rect 7193 30277 7205 30280
rect 7239 30308 7251 30311
rect 7745 30311 7803 30317
rect 7745 30308 7757 30311
rect 7239 30280 7757 30308
rect 7239 30277 7251 30280
rect 7193 30271 7251 30277
rect 7745 30277 7757 30280
rect 7791 30277 7803 30311
rect 13078 30308 13084 30320
rect 7745 30271 7803 30277
rect 8772 30280 13084 30308
rect 1857 30243 1915 30249
rect 1857 30209 1869 30243
rect 1903 30240 1915 30243
rect 2317 30243 2375 30249
rect 2317 30240 2329 30243
rect 1903 30212 2329 30240
rect 1903 30209 1915 30212
rect 1857 30203 1915 30209
rect 2317 30209 2329 30212
rect 2363 30240 2375 30243
rect 2961 30243 3019 30249
rect 2961 30240 2973 30243
rect 2363 30212 2973 30240
rect 2363 30209 2375 30212
rect 2317 30203 2375 30209
rect 2961 30209 2973 30212
rect 3007 30240 3019 30243
rect 3234 30240 3240 30252
rect 3007 30212 3240 30240
rect 3007 30209 3019 30212
rect 2961 30203 3019 30209
rect 3234 30200 3240 30212
rect 3292 30200 3298 30252
rect 4157 30243 4215 30249
rect 4157 30209 4169 30243
rect 4203 30240 4215 30243
rect 4522 30240 4528 30252
rect 4203 30212 4528 30240
rect 4203 30209 4215 30212
rect 4157 30203 4215 30209
rect 4522 30200 4528 30212
rect 4580 30240 4586 30252
rect 4706 30240 4712 30252
rect 4580 30212 4712 30240
rect 4580 30200 4586 30212
rect 4706 30200 4712 30212
rect 4764 30240 4770 30252
rect 5353 30243 5411 30249
rect 5353 30240 5365 30243
rect 4764 30212 5365 30240
rect 4764 30200 4770 30212
rect 5353 30209 5365 30212
rect 5399 30209 5411 30243
rect 5353 30203 5411 30209
rect 5718 30200 5724 30252
rect 5776 30240 5782 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 5776 30212 6561 30240
rect 5776 30200 5782 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 8662 30240 8668 30252
rect 6549 30203 6607 30209
rect 6656 30212 8668 30240
rect 1765 30175 1823 30181
rect 1765 30141 1777 30175
rect 1811 30172 1823 30175
rect 2866 30172 2872 30184
rect 1811 30144 2872 30172
rect 1811 30141 1823 30144
rect 1765 30135 1823 30141
rect 2866 30132 2872 30144
rect 2924 30132 2930 30184
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30172 3111 30175
rect 6656 30172 6684 30212
rect 8662 30200 8668 30212
rect 8720 30200 8726 30252
rect 3099 30144 6684 30172
rect 3099 30141 3111 30144
rect 3053 30135 3111 30141
rect 6822 30132 6828 30184
rect 6880 30172 6886 30184
rect 8772 30172 8800 30280
rect 13078 30268 13084 30280
rect 13136 30268 13142 30320
rect 13538 30268 13544 30320
rect 13596 30308 13602 30320
rect 14737 30311 14795 30317
rect 14737 30308 14749 30311
rect 13596 30280 14749 30308
rect 13596 30268 13602 30280
rect 14737 30277 14749 30280
rect 14783 30277 14795 30311
rect 14737 30271 14795 30277
rect 14829 30311 14887 30317
rect 14829 30277 14841 30311
rect 14875 30308 14887 30311
rect 15746 30308 15752 30320
rect 14875 30280 15752 30308
rect 14875 30277 14887 30280
rect 14829 30271 14887 30277
rect 15746 30268 15752 30280
rect 15804 30268 15810 30320
rect 16114 30308 16120 30320
rect 16075 30280 16120 30308
rect 16114 30268 16120 30280
rect 16172 30268 16178 30320
rect 9214 30200 9220 30252
rect 9272 30240 9278 30252
rect 10137 30243 10195 30249
rect 10137 30240 10149 30243
rect 9272 30212 10149 30240
rect 9272 30200 9278 30212
rect 10137 30209 10149 30212
rect 10183 30209 10195 30243
rect 10137 30203 10195 30209
rect 12250 30200 12256 30252
rect 12308 30240 12314 30252
rect 12437 30243 12495 30249
rect 12437 30240 12449 30243
rect 12308 30212 12449 30240
rect 12308 30200 12314 30212
rect 12437 30209 12449 30212
rect 12483 30209 12495 30243
rect 12437 30203 12495 30209
rect 6880 30144 8800 30172
rect 13725 30175 13783 30181
rect 6880 30132 6886 30144
rect 13725 30141 13737 30175
rect 13771 30172 13783 30175
rect 14366 30172 14372 30184
rect 13771 30144 14372 30172
rect 13771 30141 13783 30144
rect 13725 30135 13783 30141
rect 14366 30132 14372 30144
rect 14424 30132 14430 30184
rect 14734 30132 14740 30184
rect 14792 30172 14798 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 14792 30144 15577 30172
rect 14792 30132 14798 30144
rect 15565 30141 15577 30144
rect 15611 30141 15623 30175
rect 15565 30135 15623 30141
rect 16209 30175 16267 30181
rect 16209 30141 16221 30175
rect 16255 30172 16267 30175
rect 17494 30172 17500 30184
rect 16255 30144 17500 30172
rect 16255 30141 16267 30144
rect 16209 30135 16267 30141
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 4801 30107 4859 30113
rect 4801 30073 4813 30107
rect 4847 30104 4859 30107
rect 9490 30104 9496 30116
rect 4847 30076 9496 30104
rect 4847 30073 4859 30076
rect 4801 30067 4859 30073
rect 9490 30064 9496 30076
rect 9548 30064 9554 30116
rect 14277 30107 14335 30113
rect 14277 30104 14289 30107
rect 10152 30076 14289 30104
rect 6454 29996 6460 30048
rect 6512 30036 6518 30048
rect 6730 30036 6736 30048
rect 6512 30008 6736 30036
rect 6512 29996 6518 30008
rect 6730 29996 6736 30008
rect 6788 29996 6794 30048
rect 8202 29996 8208 30048
rect 8260 30036 8266 30048
rect 10152 30036 10180 30076
rect 14277 30073 14289 30076
rect 14323 30073 14335 30107
rect 14277 30067 14335 30073
rect 8260 30008 10180 30036
rect 10229 30039 10287 30045
rect 8260 29996 8266 30008
rect 10229 30005 10241 30039
rect 10275 30036 10287 30039
rect 13446 30036 13452 30048
rect 10275 30008 13452 30036
rect 10275 30005 10287 30008
rect 10229 29999 10287 30005
rect 13446 29996 13452 30008
rect 13504 29996 13510 30048
rect 16666 29996 16672 30048
rect 16724 30036 16730 30048
rect 16853 30039 16911 30045
rect 16853 30036 16865 30039
rect 16724 30008 16865 30036
rect 16724 29996 16730 30008
rect 16853 30005 16865 30008
rect 16899 30005 16911 30039
rect 17954 30036 17960 30048
rect 17915 30008 17960 30036
rect 16853 29999 16911 30005
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 18414 30036 18420 30048
rect 18375 30008 18420 30036
rect 18414 29996 18420 30008
rect 18472 29996 18478 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 2682 29792 2688 29844
rect 2740 29832 2746 29844
rect 3329 29835 3387 29841
rect 3329 29832 3341 29835
rect 2740 29804 3341 29832
rect 2740 29792 2746 29804
rect 3329 29801 3341 29804
rect 3375 29801 3387 29835
rect 4890 29832 4896 29844
rect 4851 29804 4896 29832
rect 3329 29795 3387 29801
rect 4890 29792 4896 29804
rect 4948 29792 4954 29844
rect 6549 29835 6607 29841
rect 6549 29801 6561 29835
rect 6595 29832 6607 29835
rect 7101 29835 7159 29841
rect 7101 29832 7113 29835
rect 6595 29804 7113 29832
rect 6595 29801 6607 29804
rect 6549 29795 6607 29801
rect 7101 29801 7113 29804
rect 7147 29832 7159 29835
rect 7282 29832 7288 29844
rect 7147 29804 7288 29832
rect 7147 29801 7159 29804
rect 7101 29795 7159 29801
rect 4249 29767 4307 29773
rect 4249 29733 4261 29767
rect 4295 29764 4307 29767
rect 6086 29764 6092 29776
rect 4295 29736 6092 29764
rect 4295 29733 4307 29736
rect 4249 29727 4307 29733
rect 6086 29724 6092 29736
rect 6144 29724 6150 29776
rect 2685 29699 2743 29705
rect 2685 29665 2697 29699
rect 2731 29696 2743 29699
rect 3326 29696 3332 29708
rect 2731 29668 3332 29696
rect 2731 29665 2743 29668
rect 2685 29659 2743 29665
rect 3326 29656 3332 29668
rect 3384 29656 3390 29708
rect 3602 29656 3608 29708
rect 3660 29696 3666 29708
rect 5905 29699 5963 29705
rect 5905 29696 5917 29699
rect 3660 29668 5917 29696
rect 3660 29656 3666 29668
rect 5905 29665 5917 29668
rect 5951 29665 5963 29699
rect 5905 29659 5963 29665
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 2038 29628 2044 29640
rect 1903 29600 2044 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 2593 29631 2651 29637
rect 2593 29597 2605 29631
rect 2639 29628 2651 29631
rect 3234 29628 3240 29640
rect 2639 29600 3240 29628
rect 2639 29597 2651 29600
rect 2593 29591 2651 29597
rect 3234 29588 3240 29600
rect 3292 29588 3298 29640
rect 3421 29631 3479 29637
rect 3421 29597 3433 29631
rect 3467 29628 3479 29631
rect 4157 29631 4215 29637
rect 4157 29628 4169 29631
rect 3467 29600 4169 29628
rect 3467 29597 3479 29600
rect 3421 29591 3479 29597
rect 4157 29597 4169 29600
rect 4203 29628 4215 29631
rect 4706 29628 4712 29640
rect 4203 29600 4712 29628
rect 4203 29597 4215 29600
rect 4157 29591 4215 29597
rect 4706 29588 4712 29600
rect 4764 29628 4770 29640
rect 4801 29631 4859 29637
rect 4801 29628 4813 29631
rect 4764 29600 4813 29628
rect 4764 29588 4770 29600
rect 4801 29597 4813 29600
rect 4847 29597 4859 29631
rect 4801 29591 4859 29597
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 6564 29628 6592 29795
rect 7282 29792 7288 29804
rect 7340 29832 7346 29844
rect 7742 29832 7748 29844
rect 7340 29804 7748 29832
rect 7340 29792 7346 29804
rect 7742 29792 7748 29804
rect 7800 29792 7806 29844
rect 12526 29832 12532 29844
rect 12487 29804 12532 29832
rect 12526 29792 12532 29804
rect 12584 29792 12590 29844
rect 14645 29835 14703 29841
rect 14645 29801 14657 29835
rect 14691 29832 14703 29835
rect 16114 29832 16120 29844
rect 14691 29804 16120 29832
rect 14691 29801 14703 29804
rect 14645 29795 14703 29801
rect 16114 29792 16120 29804
rect 16172 29792 16178 29844
rect 15286 29696 15292 29708
rect 15199 29668 15292 29696
rect 15286 29656 15292 29668
rect 15344 29696 15350 29708
rect 16114 29696 16120 29708
rect 15344 29668 16120 29696
rect 15344 29656 15350 29668
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 6043 29600 6592 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 6730 29588 6736 29640
rect 6788 29628 6794 29640
rect 6788 29600 10456 29628
rect 6788 29588 6794 29600
rect 10318 29560 10324 29572
rect 2746 29532 10324 29560
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 2406 29452 2412 29504
rect 2464 29492 2470 29504
rect 2746 29492 2774 29532
rect 10318 29520 10324 29532
rect 10376 29520 10382 29572
rect 10428 29560 10456 29600
rect 12250 29588 12256 29640
rect 12308 29628 12314 29640
rect 13541 29631 13599 29637
rect 13541 29628 13553 29631
rect 12308 29600 13553 29628
rect 12308 29588 12314 29600
rect 13541 29597 13553 29600
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14458 29628 14464 29640
rect 13872 29600 14464 29628
rect 13872 29588 13878 29600
rect 14458 29588 14464 29600
rect 14516 29628 14522 29640
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 14516 29600 14565 29628
rect 14516 29588 14522 29600
rect 14553 29597 14565 29600
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 16850 29588 16856 29640
rect 16908 29628 16914 29640
rect 17037 29631 17095 29637
rect 17037 29628 17049 29631
rect 16908 29600 17049 29628
rect 16908 29588 16914 29600
rect 17037 29597 17049 29600
rect 17083 29628 17095 29631
rect 18049 29631 18107 29637
rect 18049 29628 18061 29631
rect 17083 29600 18061 29628
rect 17083 29597 17095 29600
rect 17037 29591 17095 29597
rect 18049 29597 18061 29600
rect 18095 29628 18107 29631
rect 18414 29628 18420 29640
rect 18095 29600 18420 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 18414 29588 18420 29600
rect 18472 29628 18478 29640
rect 18693 29631 18751 29637
rect 18693 29628 18705 29631
rect 18472 29600 18705 29628
rect 18472 29588 18478 29600
rect 18693 29597 18705 29600
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 30101 29631 30159 29637
rect 30101 29597 30113 29631
rect 30147 29628 30159 29631
rect 37826 29628 37832 29640
rect 30147 29600 37832 29628
rect 30147 29597 30159 29600
rect 30101 29591 30159 29597
rect 37826 29588 37832 29600
rect 37884 29588 37890 29640
rect 15381 29563 15439 29569
rect 10428 29532 13124 29560
rect 13096 29501 13124 29532
rect 15381 29529 15393 29563
rect 15427 29529 15439 29563
rect 15381 29523 15439 29529
rect 16301 29563 16359 29569
rect 16301 29529 16313 29563
rect 16347 29560 16359 29563
rect 17862 29560 17868 29572
rect 16347 29532 17868 29560
rect 16347 29529 16359 29532
rect 16301 29523 16359 29529
rect 2464 29464 2774 29492
rect 13081 29495 13139 29501
rect 2464 29452 2470 29464
rect 13081 29461 13093 29495
rect 13127 29492 13139 29495
rect 13354 29492 13360 29504
rect 13127 29464 13360 29492
rect 13127 29461 13139 29464
rect 13081 29455 13139 29461
rect 13354 29452 13360 29464
rect 13412 29452 13418 29504
rect 13633 29495 13691 29501
rect 13633 29461 13645 29495
rect 13679 29492 13691 29495
rect 14274 29492 14280 29504
rect 13679 29464 14280 29492
rect 13679 29461 13691 29464
rect 13633 29455 13691 29461
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 14826 29452 14832 29504
rect 14884 29492 14890 29504
rect 15396 29492 15424 29523
rect 17862 29520 17868 29532
rect 17920 29520 17926 29572
rect 14884 29464 15424 29492
rect 17129 29495 17187 29501
rect 14884 29452 14890 29464
rect 17129 29461 17141 29495
rect 17175 29492 17187 29495
rect 17402 29492 17408 29504
rect 17175 29464 17408 29492
rect 17175 29461 17187 29464
rect 17129 29455 17187 29461
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 18141 29495 18199 29501
rect 18141 29461 18153 29495
rect 18187 29492 18199 29495
rect 18598 29492 18604 29504
rect 18187 29464 18604 29492
rect 18187 29461 18199 29464
rect 18141 29455 18199 29461
rect 18598 29452 18604 29464
rect 18656 29452 18662 29504
rect 30006 29492 30012 29504
rect 29967 29464 30012 29492
rect 30006 29452 30012 29464
rect 30064 29452 30070 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 2225 29291 2283 29297
rect 2225 29257 2237 29291
rect 2271 29288 2283 29291
rect 2314 29288 2320 29300
rect 2271 29260 2320 29288
rect 2271 29257 2283 29260
rect 2225 29251 2283 29257
rect 2314 29248 2320 29260
rect 2372 29248 2378 29300
rect 2498 29248 2504 29300
rect 2556 29288 2562 29300
rect 4157 29291 4215 29297
rect 4157 29288 4169 29291
rect 2556 29260 4169 29288
rect 2556 29248 2562 29260
rect 4157 29257 4169 29260
rect 4203 29257 4215 29291
rect 4157 29251 4215 29257
rect 5905 29291 5963 29297
rect 5905 29257 5917 29291
rect 5951 29257 5963 29291
rect 5905 29251 5963 29257
rect 2148 29192 2912 29220
rect 2148 29161 2176 29192
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29121 2191 29155
rect 2777 29155 2835 29161
rect 2777 29152 2789 29155
rect 2133 29115 2191 29121
rect 2608 29124 2789 29152
rect 1673 29019 1731 29025
rect 1673 28985 1685 29019
rect 1719 29016 1731 29019
rect 2038 29016 2044 29028
rect 1719 28988 2044 29016
rect 1719 28985 1731 28988
rect 1673 28979 1731 28985
rect 2038 28976 2044 28988
rect 2096 28976 2102 29028
rect 2608 29016 2636 29124
rect 2777 29121 2789 29124
rect 2823 29121 2835 29155
rect 2884 29152 2912 29192
rect 2958 29180 2964 29232
rect 3016 29220 3022 29232
rect 4798 29220 4804 29232
rect 3016 29192 4804 29220
rect 3016 29180 3022 29192
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 5920 29220 5948 29251
rect 6546 29248 6552 29300
rect 6604 29288 6610 29300
rect 6641 29291 6699 29297
rect 6641 29288 6653 29291
rect 6604 29260 6653 29288
rect 6604 29248 6610 29260
rect 6641 29257 6653 29260
rect 6687 29257 6699 29291
rect 7282 29288 7288 29300
rect 7243 29260 7288 29288
rect 6641 29251 6699 29257
rect 7282 29248 7288 29260
rect 7340 29248 7346 29300
rect 13538 29288 13544 29300
rect 13499 29260 13544 29288
rect 13538 29248 13544 29260
rect 13596 29248 13602 29300
rect 20346 29288 20352 29300
rect 20307 29260 20352 29288
rect 20346 29248 20352 29260
rect 20404 29248 20410 29300
rect 6822 29220 6828 29232
rect 5920 29192 6828 29220
rect 6822 29180 6828 29192
rect 6880 29180 6886 29232
rect 3234 29152 3240 29164
rect 2884 29124 3240 29152
rect 2777 29115 2835 29121
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3418 29152 3424 29164
rect 3379 29124 3424 29152
rect 3418 29112 3424 29124
rect 3476 29112 3482 29164
rect 4249 29155 4307 29161
rect 4249 29121 4261 29155
rect 4295 29152 4307 29155
rect 4706 29152 4712 29164
rect 4295 29124 4712 29152
rect 4295 29121 4307 29124
rect 4249 29115 4307 29121
rect 4706 29112 4712 29124
rect 4764 29112 4770 29164
rect 5813 29155 5871 29161
rect 5813 29121 5825 29155
rect 5859 29152 5871 29155
rect 6733 29155 6791 29161
rect 6733 29152 6745 29155
rect 5859 29124 6745 29152
rect 5859 29121 5871 29124
rect 5813 29115 5871 29121
rect 6733 29121 6745 29124
rect 6779 29152 6791 29155
rect 7300 29152 7328 29248
rect 8294 29220 8300 29232
rect 8255 29192 8300 29220
rect 8294 29180 8300 29192
rect 8352 29180 8358 29232
rect 12066 29220 12072 29232
rect 12027 29192 12072 29220
rect 12066 29180 12072 29192
rect 12124 29180 12130 29232
rect 14274 29220 14280 29232
rect 14235 29192 14280 29220
rect 14274 29180 14280 29192
rect 14332 29180 14338 29232
rect 14366 29180 14372 29232
rect 14424 29220 14430 29232
rect 15473 29223 15531 29229
rect 15473 29220 15485 29223
rect 14424 29192 15485 29220
rect 14424 29180 14430 29192
rect 15473 29189 15485 29192
rect 15519 29189 15531 29223
rect 15473 29183 15531 29189
rect 15562 29180 15568 29232
rect 15620 29220 15626 29232
rect 16298 29220 16304 29232
rect 15620 29192 16304 29220
rect 15620 29180 15626 29192
rect 16298 29180 16304 29192
rect 16356 29220 16362 29232
rect 16853 29223 16911 29229
rect 16853 29220 16865 29223
rect 16356 29192 16865 29220
rect 16356 29180 16362 29192
rect 16853 29189 16865 29192
rect 16899 29189 16911 29223
rect 17402 29220 17408 29232
rect 17363 29192 17408 29220
rect 16853 29183 16911 29189
rect 17402 29180 17408 29192
rect 17460 29180 17466 29232
rect 18046 29220 18052 29232
rect 18007 29192 18052 29220
rect 18046 29180 18052 29192
rect 18104 29180 18110 29232
rect 18598 29220 18604 29232
rect 18559 29192 18604 29220
rect 18598 29180 18604 29192
rect 18656 29180 18662 29232
rect 10318 29152 10324 29164
rect 6779 29124 7328 29152
rect 10279 29124 10324 29152
rect 6779 29121 6791 29124
rect 6733 29115 6791 29121
rect 10318 29112 10324 29124
rect 10376 29112 10382 29164
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 13449 29155 13507 29161
rect 13449 29152 13461 29155
rect 12860 29124 13461 29152
rect 12860 29112 12866 29124
rect 13449 29121 13461 29124
rect 13495 29121 13507 29155
rect 13449 29115 13507 29121
rect 19797 29155 19855 29161
rect 19797 29121 19809 29155
rect 19843 29152 19855 29155
rect 20070 29152 20076 29164
rect 19843 29124 20076 29152
rect 19843 29121 19855 29124
rect 19797 29115 19855 29121
rect 20070 29112 20076 29124
rect 20128 29152 20134 29164
rect 20364 29152 20392 29248
rect 20128 29124 20392 29152
rect 37553 29155 37611 29161
rect 20128 29112 20134 29124
rect 37553 29121 37565 29155
rect 37599 29152 37611 29155
rect 38194 29152 38200 29164
rect 37599 29124 38200 29152
rect 37599 29121 37611 29124
rect 37553 29115 37611 29121
rect 38194 29112 38200 29124
rect 38252 29112 38258 29164
rect 3513 29087 3571 29093
rect 3513 29053 3525 29087
rect 3559 29084 3571 29087
rect 7006 29084 7012 29096
rect 3559 29056 7012 29084
rect 3559 29053 3571 29056
rect 3513 29047 3571 29053
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 8202 29084 8208 29096
rect 8163 29056 8208 29084
rect 8202 29044 8208 29056
rect 8260 29044 8266 29096
rect 8849 29087 8907 29093
rect 8849 29053 8861 29087
rect 8895 29084 8907 29087
rect 9122 29084 9128 29096
rect 8895 29056 9128 29084
rect 8895 29053 8907 29056
rect 8849 29047 8907 29053
rect 9122 29044 9128 29056
rect 9180 29044 9186 29096
rect 11974 29084 11980 29096
rect 11935 29056 11980 29084
rect 11974 29044 11980 29056
rect 12032 29044 12038 29096
rect 12618 29084 12624 29096
rect 12579 29056 12624 29084
rect 12618 29044 12624 29056
rect 12676 29044 12682 29096
rect 14182 29084 14188 29096
rect 14143 29056 14188 29084
rect 14182 29044 14188 29056
rect 14240 29044 14246 29096
rect 15381 29087 15439 29093
rect 15381 29053 15393 29087
rect 15427 29084 15439 29087
rect 15470 29084 15476 29096
rect 15427 29056 15476 29084
rect 15427 29053 15439 29056
rect 15381 29047 15439 29053
rect 15470 29044 15476 29056
rect 15528 29044 15534 29096
rect 16025 29087 16083 29093
rect 16025 29053 16037 29087
rect 16071 29084 16083 29087
rect 16114 29084 16120 29096
rect 16071 29056 16120 29084
rect 16071 29053 16083 29056
rect 16025 29047 16083 29053
rect 16114 29044 16120 29056
rect 16172 29044 16178 29096
rect 17494 29084 17500 29096
rect 17407 29056 17500 29084
rect 17494 29044 17500 29056
rect 17552 29084 17558 29096
rect 18693 29087 18751 29093
rect 17552 29056 18644 29084
rect 17552 29044 17558 29056
rect 3418 29016 3424 29028
rect 2608 28988 3424 29016
rect 3418 28976 3424 28988
rect 3476 28976 3482 29028
rect 9766 29016 9772 29028
rect 5184 28988 9772 29016
rect 2869 28951 2927 28957
rect 2869 28917 2881 28951
rect 2915 28948 2927 28951
rect 2958 28948 2964 28960
rect 2915 28920 2964 28948
rect 2915 28917 2927 28920
rect 2869 28911 2927 28917
rect 2958 28908 2964 28920
rect 3016 28908 3022 28960
rect 4801 28951 4859 28957
rect 4801 28917 4813 28951
rect 4847 28948 4859 28951
rect 5184 28948 5212 28988
rect 9766 28976 9772 28988
rect 9824 28976 9830 29028
rect 10413 29019 10471 29025
rect 10413 28985 10425 29019
rect 10459 29016 10471 29019
rect 10870 29016 10876 29028
rect 10459 28988 10876 29016
rect 10459 28985 10471 28988
rect 10413 28979 10471 28985
rect 10870 28976 10876 28988
rect 10928 28976 10934 29028
rect 14734 29016 14740 29028
rect 14695 28988 14740 29016
rect 14734 28976 14740 28988
rect 14792 29016 14798 29028
rect 15194 29016 15200 29028
rect 14792 28988 15200 29016
rect 14792 28976 14798 28988
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 18616 29016 18644 29056
rect 18693 29053 18705 29087
rect 18739 29084 18751 29087
rect 19705 29087 19763 29093
rect 19705 29084 19717 29087
rect 18739 29056 19717 29084
rect 18739 29053 18751 29056
rect 18693 29047 18751 29053
rect 19705 29053 19717 29056
rect 19751 29053 19763 29087
rect 19705 29047 19763 29053
rect 30006 29016 30012 29028
rect 18616 28988 30012 29016
rect 30006 28976 30012 28988
rect 30064 28976 30070 29028
rect 37274 28976 37280 29028
rect 37332 29016 37338 29028
rect 38013 29019 38071 29025
rect 38013 29016 38025 29019
rect 37332 28988 38025 29016
rect 37332 28976 37338 28988
rect 38013 28985 38025 28988
rect 38059 28985 38071 29019
rect 38013 28979 38071 28985
rect 4847 28920 5212 28948
rect 4847 28917 4859 28920
rect 4801 28911 4859 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1673 28747 1731 28753
rect 1673 28713 1685 28747
rect 1719 28744 1731 28747
rect 2774 28744 2780 28756
rect 1719 28716 2780 28744
rect 1719 28713 1731 28716
rect 1673 28707 1731 28713
rect 2774 28704 2780 28716
rect 2832 28704 2838 28756
rect 2869 28747 2927 28753
rect 2869 28713 2881 28747
rect 2915 28744 2927 28747
rect 5350 28744 5356 28756
rect 2915 28716 5356 28744
rect 2915 28713 2927 28716
rect 2869 28707 2927 28713
rect 5350 28704 5356 28716
rect 5408 28704 5414 28756
rect 6270 28704 6276 28756
rect 6328 28744 6334 28756
rect 6549 28747 6607 28753
rect 6549 28744 6561 28747
rect 6328 28716 6561 28744
rect 6328 28704 6334 28716
rect 6549 28713 6561 28716
rect 6595 28713 6607 28747
rect 7190 28744 7196 28756
rect 7151 28716 7196 28744
rect 6549 28707 6607 28713
rect 7190 28704 7196 28716
rect 7248 28704 7254 28756
rect 7282 28704 7288 28756
rect 7340 28744 7346 28756
rect 7745 28747 7803 28753
rect 7745 28744 7757 28747
rect 7340 28716 7757 28744
rect 7340 28704 7346 28716
rect 7745 28713 7757 28716
rect 7791 28713 7803 28747
rect 11330 28744 11336 28756
rect 11291 28716 11336 28744
rect 7745 28707 7803 28713
rect 11330 28704 11336 28716
rect 11388 28704 11394 28756
rect 11977 28747 12035 28753
rect 11977 28713 11989 28747
rect 12023 28744 12035 28747
rect 12066 28744 12072 28756
rect 12023 28716 12072 28744
rect 12023 28713 12035 28716
rect 11977 28707 12035 28713
rect 12066 28704 12072 28716
rect 12124 28704 12130 28756
rect 13633 28747 13691 28753
rect 13633 28713 13645 28747
rect 13679 28744 13691 28747
rect 14366 28744 14372 28756
rect 13679 28716 14372 28744
rect 13679 28713 13691 28716
rect 13633 28707 13691 28713
rect 14366 28704 14372 28716
rect 14424 28704 14430 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 18506 28744 18512 28756
rect 14884 28716 18512 28744
rect 14884 28704 14890 28716
rect 18506 28704 18512 28716
rect 18564 28704 18570 28756
rect 2222 28676 2228 28688
rect 2183 28648 2228 28676
rect 2222 28636 2228 28648
rect 2280 28636 2286 28688
rect 2590 28636 2596 28688
rect 2648 28676 2654 28688
rect 4065 28679 4123 28685
rect 4065 28676 4077 28679
rect 2648 28648 4077 28676
rect 2648 28636 2654 28648
rect 4065 28645 4077 28648
rect 4111 28645 4123 28679
rect 4065 28639 4123 28645
rect 5905 28679 5963 28685
rect 5905 28645 5917 28679
rect 5951 28676 5963 28679
rect 9858 28676 9864 28688
rect 5951 28648 9864 28676
rect 5951 28645 5963 28648
rect 5905 28639 5963 28645
rect 9858 28636 9864 28648
rect 9916 28636 9922 28688
rect 12526 28636 12532 28688
rect 12584 28676 12590 28688
rect 17678 28676 17684 28688
rect 12584 28648 13584 28676
rect 12584 28636 12590 28648
rect 4801 28611 4859 28617
rect 4801 28577 4813 28611
rect 4847 28608 4859 28611
rect 8478 28608 8484 28620
rect 4847 28580 8484 28608
rect 4847 28577 4859 28580
rect 4801 28571 4859 28577
rect 8478 28568 8484 28580
rect 8536 28568 8542 28620
rect 9769 28611 9827 28617
rect 9769 28577 9781 28611
rect 9815 28608 9827 28611
rect 12618 28608 12624 28620
rect 9815 28580 12624 28608
rect 9815 28577 9827 28580
rect 9769 28571 9827 28577
rect 12618 28568 12624 28580
rect 12676 28568 12682 28620
rect 2133 28543 2191 28549
rect 2133 28509 2145 28543
rect 2179 28540 2191 28543
rect 2774 28540 2780 28552
rect 2179 28512 2780 28540
rect 2179 28509 2191 28512
rect 2133 28503 2191 28509
rect 2774 28500 2780 28512
rect 2832 28540 2838 28552
rect 3234 28540 3240 28552
rect 2832 28512 3240 28540
rect 2832 28500 2838 28512
rect 3234 28500 3240 28512
rect 3292 28500 3298 28552
rect 3418 28500 3424 28552
rect 3476 28540 3482 28552
rect 4157 28543 4215 28549
rect 4157 28540 4169 28543
rect 3476 28512 4169 28540
rect 3476 28500 3482 28512
rect 4157 28509 4169 28512
rect 4203 28509 4215 28543
rect 4706 28540 4712 28552
rect 4667 28512 4712 28540
rect 4157 28503 4215 28509
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5813 28543 5871 28549
rect 5813 28509 5825 28543
rect 5859 28540 5871 28543
rect 6457 28543 6515 28549
rect 6457 28540 6469 28543
rect 5859 28512 6469 28540
rect 5859 28509 5871 28512
rect 5813 28503 5871 28509
rect 6457 28509 6469 28512
rect 6503 28540 6515 28543
rect 7101 28543 7159 28549
rect 7101 28540 7113 28543
rect 6503 28512 7113 28540
rect 6503 28509 6515 28512
rect 6457 28503 6515 28509
rect 7101 28509 7113 28512
rect 7147 28540 7159 28543
rect 7282 28540 7288 28552
rect 7147 28512 7288 28540
rect 7147 28509 7159 28512
rect 7101 28503 7159 28509
rect 7282 28500 7288 28512
rect 7340 28500 7346 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10505 28543 10563 28549
rect 10505 28540 10517 28543
rect 10008 28512 10517 28540
rect 10008 28500 10014 28512
rect 10505 28509 10517 28512
rect 10551 28509 10563 28543
rect 11882 28540 11888 28552
rect 11843 28512 11888 28540
rect 10505 28503 10563 28509
rect 11882 28500 11888 28512
rect 11940 28540 11946 28552
rect 12802 28540 12808 28552
rect 11940 28512 12808 28540
rect 11940 28500 11946 28512
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 12894 28500 12900 28552
rect 12952 28540 12958 28552
rect 13556 28549 13584 28648
rect 14200 28648 17684 28676
rect 13541 28543 13599 28549
rect 12952 28512 12997 28540
rect 12952 28500 12958 28512
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 14200 28540 14228 28648
rect 17678 28636 17684 28648
rect 17736 28636 17742 28688
rect 14369 28611 14427 28617
rect 14369 28577 14381 28611
rect 14415 28608 14427 28611
rect 14734 28608 14740 28620
rect 14415 28580 14740 28608
rect 14415 28577 14427 28580
rect 14369 28571 14427 28577
rect 14734 28568 14740 28580
rect 14792 28568 14798 28620
rect 15378 28608 15384 28620
rect 15339 28580 15384 28608
rect 15378 28568 15384 28580
rect 15436 28568 15442 28620
rect 16577 28611 16635 28617
rect 16577 28577 16589 28611
rect 16623 28608 16635 28611
rect 16850 28608 16856 28620
rect 16623 28580 16856 28608
rect 16623 28577 16635 28580
rect 16577 28571 16635 28577
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 17589 28611 17647 28617
rect 17589 28577 17601 28611
rect 17635 28608 17647 28611
rect 17862 28608 17868 28620
rect 17635 28580 17868 28608
rect 17635 28577 17647 28580
rect 17589 28571 17647 28577
rect 17862 28568 17868 28580
rect 17920 28608 17926 28620
rect 17920 28580 26234 28608
rect 17920 28568 17926 28580
rect 16022 28540 16028 28552
rect 13587 28512 14228 28540
rect 15983 28512 16028 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 16022 28500 16028 28512
rect 16080 28500 16086 28552
rect 17954 28500 17960 28552
rect 18012 28540 18018 28552
rect 18233 28543 18291 28549
rect 18233 28540 18245 28543
rect 18012 28512 18245 28540
rect 18012 28500 18018 28512
rect 18233 28509 18245 28512
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 9122 28472 9128 28484
rect 9083 28444 9128 28472
rect 9122 28432 9128 28444
rect 9180 28432 9186 28484
rect 9674 28472 9680 28484
rect 9635 28444 9680 28472
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 10597 28475 10655 28481
rect 10597 28441 10609 28475
rect 10643 28472 10655 28475
rect 13262 28472 13268 28484
rect 10643 28444 13268 28472
rect 10643 28441 10655 28444
rect 10597 28435 10655 28441
rect 13262 28432 13268 28444
rect 13320 28432 13326 28484
rect 14458 28432 14464 28484
rect 14516 28472 14522 28484
rect 16669 28475 16727 28481
rect 14516 28444 14561 28472
rect 14516 28432 14522 28444
rect 16669 28441 16681 28475
rect 16715 28441 16727 28475
rect 18248 28472 18276 28503
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18693 28543 18751 28549
rect 18693 28540 18705 28543
rect 18472 28512 18705 28540
rect 18472 28500 18478 28512
rect 18693 28509 18705 28512
rect 18739 28509 18751 28543
rect 20070 28540 20076 28552
rect 20031 28512 20076 28540
rect 18693 28503 18751 28509
rect 20070 28500 20076 28512
rect 20128 28540 20134 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 20128 28512 20637 28540
rect 20128 28500 20134 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 20625 28503 20683 28509
rect 18506 28472 18512 28484
rect 18248 28444 18512 28472
rect 16669 28435 16727 28441
rect 1854 28364 1860 28416
rect 1912 28404 1918 28416
rect 7374 28404 7380 28416
rect 1912 28376 7380 28404
rect 1912 28364 1918 28376
rect 7374 28364 7380 28376
rect 7432 28364 7438 28416
rect 12989 28407 13047 28413
rect 12989 28373 13001 28407
rect 13035 28404 13047 28407
rect 13170 28404 13176 28416
rect 13035 28376 13176 28404
rect 13035 28373 13047 28376
rect 12989 28367 13047 28373
rect 13170 28364 13176 28376
rect 13228 28364 13234 28416
rect 15746 28364 15752 28416
rect 15804 28404 15810 28416
rect 15933 28407 15991 28413
rect 15933 28404 15945 28407
rect 15804 28376 15945 28404
rect 15804 28364 15810 28376
rect 15933 28373 15945 28376
rect 15979 28373 15991 28407
rect 15933 28367 15991 28373
rect 16206 28364 16212 28416
rect 16264 28404 16270 28416
rect 16684 28404 16712 28435
rect 18506 28432 18512 28444
rect 18564 28432 18570 28484
rect 26206 28472 26234 28580
rect 37826 28540 37832 28552
rect 37787 28512 37832 28540
rect 37826 28500 37832 28512
rect 37884 28500 37890 28552
rect 36262 28472 36268 28484
rect 26206 28444 36268 28472
rect 36262 28432 36268 28444
rect 36320 28432 36326 28484
rect 16264 28376 16712 28404
rect 16264 28364 16270 28376
rect 16758 28364 16764 28416
rect 16816 28404 16822 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 16816 28376 18153 28404
rect 16816 28364 16822 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 18782 28404 18788 28416
rect 18743 28376 18788 28404
rect 18141 28367 18199 28373
rect 18782 28364 18788 28376
rect 18840 28364 18846 28416
rect 19981 28407 20039 28413
rect 19981 28373 19993 28407
rect 20027 28404 20039 28407
rect 20438 28404 20444 28416
rect 20027 28376 20444 28404
rect 20027 28373 20039 28376
rect 19981 28367 20039 28373
rect 20438 28364 20444 28376
rect 20496 28364 20502 28416
rect 38010 28404 38016 28416
rect 37971 28376 38016 28404
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3510 28200 3516 28212
rect 3471 28172 3516 28200
rect 3510 28160 3516 28172
rect 3568 28160 3574 28212
rect 4157 28203 4215 28209
rect 4157 28169 4169 28203
rect 4203 28200 4215 28203
rect 4614 28200 4620 28212
rect 4203 28172 4620 28200
rect 4203 28169 4215 28172
rect 4157 28163 4215 28169
rect 4614 28160 4620 28172
rect 4672 28160 4678 28212
rect 5997 28203 6055 28209
rect 5997 28169 6009 28203
rect 6043 28200 6055 28203
rect 6825 28203 6883 28209
rect 6825 28200 6837 28203
rect 6043 28172 6837 28200
rect 6043 28169 6055 28172
rect 5997 28163 6055 28169
rect 6825 28169 6837 28172
rect 6871 28200 6883 28203
rect 7282 28200 7288 28212
rect 6871 28172 7288 28200
rect 6871 28169 6883 28172
rect 6825 28163 6883 28169
rect 7282 28160 7288 28172
rect 7340 28160 7346 28212
rect 11793 28203 11851 28209
rect 11793 28169 11805 28203
rect 11839 28200 11851 28203
rect 14458 28200 14464 28212
rect 11839 28172 14464 28200
rect 11839 28169 11851 28172
rect 11793 28163 11851 28169
rect 14458 28160 14464 28172
rect 14516 28160 14522 28212
rect 2869 28135 2927 28141
rect 2869 28101 2881 28135
rect 2915 28132 2927 28135
rect 7098 28132 7104 28144
rect 2915 28104 7104 28132
rect 2915 28101 2927 28104
rect 2869 28095 2927 28101
rect 7098 28092 7104 28104
rect 7156 28092 7162 28144
rect 7558 28092 7564 28144
rect 7616 28132 7622 28144
rect 11882 28132 11888 28144
rect 7616 28104 11888 28132
rect 7616 28092 7622 28104
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28033 1915 28067
rect 1857 28027 1915 28033
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 1872 27860 1900 28027
rect 2774 28024 2780 28076
rect 2832 28064 2838 28076
rect 2832 28036 2877 28064
rect 2832 28024 2838 28036
rect 3418 28024 3424 28076
rect 3476 28064 3482 28076
rect 3605 28067 3663 28073
rect 3605 28064 3617 28067
rect 3476 28036 3617 28064
rect 3476 28024 3482 28036
rect 3605 28033 3617 28036
rect 3651 28033 3663 28067
rect 3605 28027 3663 28033
rect 10137 28067 10195 28073
rect 10137 28033 10149 28067
rect 10183 28064 10195 28067
rect 10226 28064 10232 28076
rect 10183 28036 10232 28064
rect 10183 28033 10195 28036
rect 10137 28027 10195 28033
rect 10226 28024 10232 28036
rect 10284 28024 10290 28076
rect 10796 28073 10824 28104
rect 11882 28092 11888 28104
rect 11940 28092 11946 28144
rect 13630 28132 13636 28144
rect 12452 28104 13636 28132
rect 12452 28073 12480 28104
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 13814 28092 13820 28144
rect 13872 28132 13878 28144
rect 14553 28135 14611 28141
rect 14553 28132 14565 28135
rect 13872 28104 14565 28132
rect 13872 28092 13878 28104
rect 14553 28101 14565 28104
rect 14599 28101 14611 28135
rect 15746 28132 15752 28144
rect 15707 28104 15752 28132
rect 14553 28095 14611 28101
rect 15746 28092 15752 28104
rect 15804 28092 15810 28144
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 18049 28135 18107 28141
rect 18049 28132 18061 28135
rect 15988 28104 18061 28132
rect 15988 28092 15994 28104
rect 18049 28101 18061 28104
rect 18095 28101 18107 28135
rect 18049 28095 18107 28101
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10781 28027 10839 28033
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 7374 27956 7380 28008
rect 7432 27996 7438 28008
rect 11716 27996 11744 28027
rect 12894 28024 12900 28076
rect 12952 28064 12958 28076
rect 13081 28067 13139 28073
rect 13081 28064 13093 28067
rect 12952 28036 13093 28064
rect 12952 28024 12958 28036
rect 13081 28033 13093 28036
rect 13127 28033 13139 28067
rect 13081 28027 13139 28033
rect 13354 28024 13360 28076
rect 13412 28064 13418 28076
rect 13722 28064 13728 28076
rect 13412 28036 13728 28064
rect 13412 28024 13418 28036
rect 13722 28024 13728 28036
rect 13780 28024 13786 28076
rect 16298 28024 16304 28076
rect 16356 28064 16362 28076
rect 23658 28064 23664 28076
rect 16356 28036 16401 28064
rect 23619 28036 23664 28064
rect 16356 28024 16362 28036
rect 23658 28024 23664 28036
rect 23716 28064 23722 28076
rect 24305 28067 24363 28073
rect 24305 28064 24317 28067
rect 23716 28036 24317 28064
rect 23716 28024 23722 28036
rect 24305 28033 24317 28036
rect 24351 28033 24363 28067
rect 24305 28027 24363 28033
rect 7432 27968 11744 27996
rect 13173 27999 13231 28005
rect 7432 27956 7438 27968
rect 13173 27965 13185 27999
rect 13219 27996 13231 27999
rect 14274 27996 14280 28008
rect 13219 27968 14280 27996
rect 13219 27965 13231 27968
rect 13173 27959 13231 27965
rect 14274 27956 14280 27968
rect 14332 27956 14338 28008
rect 14461 27999 14519 28005
rect 14461 27965 14473 27999
rect 14507 27996 14519 27999
rect 15470 27996 15476 28008
rect 14507 27968 15476 27996
rect 14507 27965 14519 27968
rect 14461 27959 14519 27965
rect 15470 27956 15476 27968
rect 15528 27956 15534 28008
rect 15657 27999 15715 28005
rect 15657 27965 15669 27999
rect 15703 27965 15715 27999
rect 17862 27996 17868 28008
rect 17823 27968 17868 27996
rect 15657 27959 15715 27965
rect 12434 27928 12440 27940
rect 9646 27900 12440 27928
rect 9646 27860 9674 27900
rect 12434 27888 12440 27900
rect 12492 27888 12498 27940
rect 12529 27931 12587 27937
rect 12529 27897 12541 27931
rect 12575 27928 12587 27931
rect 14550 27928 14556 27940
rect 12575 27900 14556 27928
rect 12575 27897 12587 27900
rect 12529 27891 12587 27897
rect 14550 27888 14556 27900
rect 14608 27888 14614 27940
rect 15013 27931 15071 27937
rect 15013 27897 15025 27931
rect 15059 27928 15071 27931
rect 15378 27928 15384 27940
rect 15059 27900 15384 27928
rect 15059 27897 15071 27900
rect 15013 27891 15071 27897
rect 15378 27888 15384 27900
rect 15436 27888 15442 27940
rect 10042 27860 10048 27872
rect 1872 27832 9674 27860
rect 10003 27832 10048 27860
rect 10042 27820 10048 27832
rect 10100 27820 10106 27872
rect 10873 27863 10931 27869
rect 10873 27829 10885 27863
rect 10919 27860 10931 27863
rect 10962 27860 10968 27872
rect 10919 27832 10968 27860
rect 10919 27829 10931 27832
rect 10873 27823 10931 27829
rect 10962 27820 10968 27832
rect 11020 27820 11026 27872
rect 13817 27863 13875 27869
rect 13817 27829 13829 27863
rect 13863 27860 13875 27863
rect 14182 27860 14188 27872
rect 13863 27832 14188 27860
rect 13863 27829 13875 27832
rect 13817 27823 13875 27829
rect 14182 27820 14188 27832
rect 14240 27860 14246 27872
rect 15672 27860 15700 27959
rect 17862 27956 17868 27968
rect 17920 27956 17926 28008
rect 18138 27996 18144 28008
rect 18099 27968 18144 27996
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 18690 27996 18696 28008
rect 18651 27968 18696 27996
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 19334 27996 19340 28008
rect 19295 27968 19340 27996
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 20073 27931 20131 27937
rect 20073 27897 20085 27931
rect 20119 27928 20131 27931
rect 20346 27928 20352 27940
rect 20119 27900 20352 27928
rect 20119 27897 20131 27900
rect 20073 27891 20131 27897
rect 20346 27888 20352 27900
rect 20404 27928 20410 27940
rect 23845 27931 23903 27937
rect 20404 27900 22094 27928
rect 20404 27888 20410 27900
rect 14240 27832 15700 27860
rect 14240 27820 14246 27832
rect 17310 27820 17316 27872
rect 17368 27860 17374 27872
rect 19978 27860 19984 27872
rect 17368 27832 19984 27860
rect 17368 27820 17374 27832
rect 19978 27820 19984 27832
rect 20036 27860 20042 27872
rect 20533 27863 20591 27869
rect 20533 27860 20545 27863
rect 20036 27832 20545 27860
rect 20036 27820 20042 27832
rect 20533 27829 20545 27832
rect 20579 27829 20591 27863
rect 22066 27860 22094 27900
rect 23845 27897 23857 27931
rect 23891 27928 23903 27931
rect 34790 27928 34796 27940
rect 23891 27900 34796 27928
rect 23891 27897 23903 27900
rect 23845 27891 23903 27897
rect 34790 27888 34796 27900
rect 34848 27888 34854 27940
rect 38286 27860 38292 27872
rect 22066 27832 38292 27860
rect 20533 27823 20591 27829
rect 38286 27820 38292 27832
rect 38344 27820 38350 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 10042 27616 10048 27668
rect 10100 27656 10106 27668
rect 14642 27656 14648 27668
rect 10100 27628 14648 27656
rect 10100 27616 10106 27628
rect 14642 27616 14648 27628
rect 14700 27616 14706 27668
rect 16022 27616 16028 27668
rect 16080 27656 16086 27668
rect 17310 27656 17316 27668
rect 16080 27628 17316 27656
rect 16080 27616 16086 27628
rect 17310 27616 17316 27628
rect 17368 27616 17374 27668
rect 1578 27588 1584 27600
rect 1539 27560 1584 27588
rect 1578 27548 1584 27560
rect 1636 27548 1642 27600
rect 11238 27548 11244 27600
rect 11296 27588 11302 27600
rect 14366 27588 14372 27600
rect 11296 27560 14372 27588
rect 11296 27548 11302 27560
rect 14366 27548 14372 27560
rect 14424 27548 14430 27600
rect 14734 27548 14740 27600
rect 14792 27588 14798 27600
rect 17770 27588 17776 27600
rect 14792 27560 17776 27588
rect 14792 27548 14798 27560
rect 17770 27548 17776 27560
rect 17828 27548 17834 27600
rect 21177 27591 21235 27597
rect 21177 27588 21189 27591
rect 17880 27560 21189 27588
rect 9769 27523 9827 27529
rect 9769 27489 9781 27523
rect 9815 27520 9827 27523
rect 11149 27523 11207 27529
rect 11149 27520 11161 27523
rect 9815 27492 11161 27520
rect 9815 27489 9827 27492
rect 9769 27483 9827 27489
rect 11149 27489 11161 27492
rect 11195 27520 11207 27523
rect 11195 27492 12434 27520
rect 11195 27489 11207 27492
rect 11149 27483 11207 27489
rect 11977 27455 12035 27461
rect 11977 27421 11989 27455
rect 12023 27421 12035 27455
rect 11977 27415 12035 27421
rect 9122 27384 9128 27396
rect 9083 27356 9128 27384
rect 9122 27344 9128 27356
rect 9180 27344 9186 27396
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9640 27356 9689 27384
rect 9640 27344 9646 27356
rect 9677 27353 9689 27356
rect 9723 27353 9735 27387
rect 10870 27384 10876 27396
rect 10831 27356 10876 27384
rect 9677 27347 9735 27353
rect 10870 27344 10876 27356
rect 10928 27344 10934 27396
rect 10962 27344 10968 27396
rect 11020 27384 11026 27396
rect 11020 27356 11065 27384
rect 11020 27344 11026 27356
rect 11330 27344 11336 27396
rect 11388 27384 11394 27396
rect 11992 27384 12020 27415
rect 11388 27356 12020 27384
rect 12406 27384 12434 27492
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 13354 27520 13360 27532
rect 12584 27492 13360 27520
rect 12584 27480 12590 27492
rect 13354 27480 13360 27492
rect 13412 27480 13418 27532
rect 15657 27523 15715 27529
rect 15657 27489 15669 27523
rect 15703 27520 15715 27523
rect 15838 27520 15844 27532
rect 15703 27492 15844 27520
rect 15703 27489 15715 27492
rect 15657 27483 15715 27489
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 15933 27523 15991 27529
rect 15933 27489 15945 27523
rect 15979 27520 15991 27523
rect 16482 27520 16488 27532
rect 15979 27492 16488 27520
rect 15979 27489 15991 27492
rect 15933 27483 15991 27489
rect 16482 27480 16488 27492
rect 16540 27480 16546 27532
rect 16850 27520 16856 27532
rect 16811 27492 16856 27520
rect 16850 27480 16856 27492
rect 16908 27480 16914 27532
rect 17126 27520 17132 27532
rect 17087 27492 17132 27520
rect 17126 27480 17132 27492
rect 17184 27520 17190 27532
rect 17880 27520 17908 27560
rect 21177 27557 21189 27560
rect 21223 27557 21235 27591
rect 21177 27551 21235 27557
rect 17184 27492 17908 27520
rect 17184 27480 17190 27492
rect 17954 27480 17960 27532
rect 18012 27520 18018 27532
rect 18325 27523 18383 27529
rect 18012 27492 18057 27520
rect 18012 27480 18018 27492
rect 18325 27489 18337 27523
rect 18371 27520 18383 27523
rect 19334 27520 19340 27532
rect 18371 27492 19340 27520
rect 18371 27489 18383 27492
rect 18325 27483 18383 27489
rect 19334 27480 19340 27492
rect 19392 27480 19398 27532
rect 14366 27412 14372 27464
rect 14424 27452 14430 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14424 27424 14657 27452
rect 14424 27412 14430 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 18564 27424 19625 27452
rect 18564 27412 18570 27424
rect 19613 27421 19625 27424
rect 19659 27452 19671 27455
rect 20625 27455 20683 27461
rect 20625 27452 20637 27455
rect 19659 27424 20637 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 20625 27421 20637 27424
rect 20671 27421 20683 27455
rect 20625 27415 20683 27421
rect 12802 27384 12808 27396
rect 12406 27356 12808 27384
rect 11388 27344 11394 27356
rect 12802 27344 12808 27356
rect 12860 27344 12866 27396
rect 13078 27384 13084 27396
rect 13039 27356 13084 27384
rect 13078 27344 13084 27356
rect 13136 27344 13142 27396
rect 13170 27344 13176 27396
rect 13228 27384 13234 27396
rect 13228 27356 13273 27384
rect 13228 27344 13234 27356
rect 14274 27344 14280 27396
rect 14332 27384 14338 27396
rect 15654 27384 15660 27396
rect 14332 27356 15660 27384
rect 14332 27344 14338 27356
rect 15654 27344 15660 27356
rect 15712 27344 15718 27396
rect 15841 27387 15899 27393
rect 15841 27353 15853 27387
rect 15887 27353 15899 27387
rect 15841 27347 15899 27353
rect 12069 27319 12127 27325
rect 12069 27285 12081 27319
rect 12115 27316 12127 27319
rect 12710 27316 12716 27328
rect 12115 27288 12716 27316
rect 12115 27285 12127 27288
rect 12069 27279 12127 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 14737 27319 14795 27325
rect 14737 27285 14749 27319
rect 14783 27316 14795 27319
rect 15746 27316 15752 27328
rect 14783 27288 15752 27316
rect 14783 27285 14795 27288
rect 14737 27279 14795 27285
rect 15746 27276 15752 27288
rect 15804 27276 15810 27328
rect 15856 27316 15884 27347
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 16850 27384 16856 27396
rect 15988 27356 16856 27384
rect 15988 27344 15994 27356
rect 16850 27344 16856 27356
rect 16908 27344 16914 27396
rect 17037 27387 17095 27393
rect 17037 27353 17049 27387
rect 17083 27384 17095 27387
rect 18233 27387 18291 27393
rect 17083 27356 18184 27384
rect 17083 27353 17095 27356
rect 17037 27347 17095 27353
rect 16758 27316 16764 27328
rect 15856 27288 16764 27316
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 18156 27316 18184 27356
rect 18233 27353 18245 27387
rect 18279 27384 18291 27387
rect 18782 27384 18788 27396
rect 18279 27356 18788 27384
rect 18279 27353 18291 27356
rect 18233 27347 18291 27353
rect 18782 27344 18788 27356
rect 18840 27344 18846 27396
rect 20070 27384 20076 27396
rect 20031 27356 20076 27384
rect 20070 27344 20076 27356
rect 20128 27344 20134 27396
rect 18322 27316 18328 27328
rect 18156 27288 18328 27316
rect 18322 27276 18328 27288
rect 18380 27276 18386 27328
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 19521 27319 19579 27325
rect 19521 27316 19533 27319
rect 18472 27288 19533 27316
rect 18472 27276 18478 27288
rect 19521 27285 19533 27288
rect 19567 27285 19579 27319
rect 19521 27279 19579 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 9401 27115 9459 27121
rect 9401 27112 9413 27115
rect 8444 27084 9413 27112
rect 8444 27072 8450 27084
rect 9401 27081 9413 27084
rect 9447 27112 9459 27115
rect 12342 27112 12348 27124
rect 9447 27084 12348 27112
rect 9447 27081 9459 27084
rect 9401 27075 9459 27081
rect 12342 27072 12348 27084
rect 12400 27112 12406 27124
rect 12805 27115 12863 27121
rect 12400 27084 12664 27112
rect 12400 27072 12406 27084
rect 8941 26979 8999 26985
rect 8941 26945 8953 26979
rect 8987 26976 8999 26979
rect 12069 26979 12127 26985
rect 12069 26976 12081 26979
rect 8987 26948 12081 26976
rect 8987 26945 8999 26948
rect 8941 26939 8999 26945
rect 12069 26945 12081 26948
rect 12115 26945 12127 26979
rect 12636 26976 12664 27084
rect 12805 27081 12817 27115
rect 12851 27112 12863 27115
rect 13814 27112 13820 27124
rect 12851 27084 13820 27112
rect 12851 27081 12863 27084
rect 12805 27075 12863 27081
rect 13814 27072 13820 27084
rect 13872 27072 13878 27124
rect 14182 27072 14188 27124
rect 14240 27112 14246 27124
rect 17218 27112 17224 27124
rect 14240 27084 17224 27112
rect 14240 27072 14246 27084
rect 13354 27004 13360 27056
rect 13412 27044 13418 27056
rect 14001 27047 14059 27053
rect 14001 27044 14013 27047
rect 13412 27016 14013 27044
rect 13412 27004 13418 27016
rect 14001 27013 14013 27016
rect 14047 27013 14059 27047
rect 14550 27044 14556 27056
rect 14511 27016 14556 27044
rect 14001 27007 14059 27013
rect 14550 27004 14556 27016
rect 14608 27004 14614 27056
rect 14660 27053 14688 27084
rect 17218 27072 17224 27084
rect 17276 27072 17282 27124
rect 17402 27072 17408 27124
rect 17460 27112 17466 27124
rect 37274 27112 37280 27124
rect 17460 27084 37280 27112
rect 17460 27072 17466 27084
rect 37274 27072 37280 27084
rect 37332 27072 37338 27124
rect 14645 27047 14703 27053
rect 14645 27013 14657 27047
rect 14691 27013 14703 27047
rect 14645 27007 14703 27013
rect 15654 27004 15660 27056
rect 15712 27044 15718 27056
rect 15749 27047 15807 27053
rect 15749 27044 15761 27047
rect 15712 27016 15761 27044
rect 15712 27004 15718 27016
rect 15749 27013 15761 27016
rect 15795 27013 15807 27047
rect 15749 27007 15807 27013
rect 15841 27047 15899 27053
rect 15841 27013 15853 27047
rect 15887 27044 15899 27047
rect 16758 27044 16764 27056
rect 15887 27016 16764 27044
rect 15887 27013 15899 27016
rect 15841 27007 15899 27013
rect 16758 27004 16764 27016
rect 16816 27004 16822 27056
rect 18230 27044 18236 27056
rect 16868 27016 18236 27044
rect 12713 26979 12771 26985
rect 12713 26976 12725 26979
rect 12636 26948 12725 26976
rect 12069 26939 12127 26945
rect 12713 26945 12725 26948
rect 12759 26945 12771 26979
rect 13538 26976 13544 26988
rect 13451 26948 13544 26976
rect 12713 26939 12771 26945
rect 10042 26908 10048 26920
rect 10003 26880 10048 26908
rect 10042 26868 10048 26880
rect 10100 26868 10106 26920
rect 10594 26908 10600 26920
rect 10555 26880 10600 26908
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 12084 26908 12112 26939
rect 13538 26936 13544 26948
rect 13596 26976 13602 26988
rect 13596 26948 14044 26976
rect 13596 26936 13602 26948
rect 12250 26908 12256 26920
rect 12084 26880 12256 26908
rect 12250 26868 12256 26880
rect 12308 26908 12314 26920
rect 12308 26880 13492 26908
rect 12308 26868 12314 26880
rect 11149 26843 11207 26849
rect 11149 26809 11161 26843
rect 11195 26840 11207 26843
rect 11238 26840 11244 26852
rect 11195 26812 11244 26840
rect 11195 26809 11207 26812
rect 11149 26803 11207 26809
rect 11238 26800 11244 26812
rect 11296 26800 11302 26852
rect 12161 26843 12219 26849
rect 12161 26809 12173 26843
rect 12207 26840 12219 26843
rect 13078 26840 13084 26852
rect 12207 26812 13084 26840
rect 12207 26809 12219 26812
rect 12161 26803 12219 26809
rect 13078 26800 13084 26812
rect 13136 26800 13142 26852
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 13357 26775 13415 26781
rect 13357 26772 13369 26775
rect 12492 26744 13369 26772
rect 12492 26732 12498 26744
rect 13357 26741 13369 26744
rect 13403 26741 13415 26775
rect 13464 26772 13492 26880
rect 14016 26840 14044 26948
rect 15194 26908 15200 26920
rect 15155 26880 15200 26908
rect 15194 26868 15200 26880
rect 15252 26868 15258 26920
rect 16868 26908 16896 27016
rect 18230 27004 18236 27016
rect 18288 27004 18294 27056
rect 18414 27044 18420 27056
rect 18375 27016 18420 27044
rect 18414 27004 18420 27016
rect 18472 27004 18478 27056
rect 18509 27047 18567 27053
rect 18509 27013 18521 27047
rect 18555 27044 18567 27047
rect 18690 27044 18696 27056
rect 18555 27016 18696 27044
rect 18555 27013 18567 27016
rect 18509 27007 18567 27013
rect 18690 27004 18696 27016
rect 18748 27004 18754 27056
rect 19610 27044 19616 27056
rect 19260 27016 19616 27044
rect 17310 26936 17316 26988
rect 17368 26976 17374 26988
rect 19260 26985 19288 27016
rect 19610 27004 19616 27016
rect 19668 27044 19674 27056
rect 20346 27044 20352 27056
rect 19668 27016 20352 27044
rect 19668 27004 19674 27016
rect 20346 27004 20352 27016
rect 20404 27004 20410 27056
rect 19245 26979 19303 26985
rect 17368 26948 17413 26976
rect 17368 26936 17374 26948
rect 19245 26945 19257 26979
rect 19291 26945 19303 26979
rect 19245 26939 19303 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 38010 26976 38016 26988
rect 19935 26948 20392 26976
rect 37971 26948 38016 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 18138 26908 18144 26920
rect 15304 26880 16896 26908
rect 18099 26880 18144 26908
rect 15304 26840 15332 26880
rect 18138 26868 18144 26880
rect 18196 26868 18202 26920
rect 18230 26868 18236 26920
rect 18288 26908 18294 26920
rect 20162 26908 20168 26920
rect 18288 26880 20168 26908
rect 18288 26868 18294 26880
rect 20162 26868 20168 26880
rect 20220 26868 20226 26920
rect 17402 26840 17408 26852
rect 14016 26812 15332 26840
rect 15396 26812 17408 26840
rect 15396 26772 15424 26812
rect 17402 26800 17408 26812
rect 17460 26800 17466 26852
rect 17494 26800 17500 26852
rect 17552 26840 17558 26852
rect 19797 26843 19855 26849
rect 19797 26840 19809 26843
rect 17552 26812 19809 26840
rect 17552 26800 17558 26812
rect 19797 26809 19809 26812
rect 19843 26809 19855 26843
rect 19797 26803 19855 26809
rect 20364 26784 20392 26948
rect 38010 26936 38016 26948
rect 38068 26936 38074 26988
rect 13464 26744 15424 26772
rect 13357 26735 13415 26741
rect 17034 26732 17040 26784
rect 17092 26772 17098 26784
rect 17221 26775 17279 26781
rect 17221 26772 17233 26775
rect 17092 26744 17233 26772
rect 17092 26732 17098 26744
rect 17221 26741 17233 26744
rect 17267 26741 17279 26775
rect 17221 26735 17279 26741
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 19153 26775 19211 26781
rect 19153 26772 19165 26775
rect 18840 26744 19165 26772
rect 18840 26732 18846 26744
rect 19153 26741 19165 26744
rect 19199 26741 19211 26775
rect 19153 26735 19211 26741
rect 20346 26732 20352 26784
rect 20404 26772 20410 26784
rect 20901 26775 20959 26781
rect 20901 26772 20913 26775
rect 20404 26744 20913 26772
rect 20404 26732 20410 26744
rect 20901 26741 20913 26744
rect 20947 26741 20959 26775
rect 38194 26772 38200 26784
rect 38155 26744 38200 26772
rect 20901 26735 20959 26741
rect 38194 26732 38200 26744
rect 38252 26732 38258 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 11974 26528 11980 26580
rect 12032 26568 12038 26580
rect 16942 26568 16948 26580
rect 12032 26540 16948 26568
rect 12032 26528 12038 26540
rect 16942 26528 16948 26540
rect 17000 26528 17006 26580
rect 17678 26528 17684 26580
rect 17736 26568 17742 26580
rect 20070 26568 20076 26580
rect 17736 26540 20076 26568
rect 17736 26528 17742 26540
rect 20070 26528 20076 26540
rect 20128 26528 20134 26580
rect 14734 26500 14740 26512
rect 12544 26472 14740 26500
rect 9398 26392 9404 26444
rect 9456 26432 9462 26444
rect 12069 26435 12127 26441
rect 9456 26404 10732 26432
rect 9456 26392 9462 26404
rect 1854 26364 1860 26376
rect 1815 26336 1860 26364
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 10704 26373 10732 26404
rect 12069 26401 12081 26435
rect 12115 26432 12127 26435
rect 12544 26432 12572 26472
rect 14734 26460 14740 26472
rect 14792 26460 14798 26512
rect 17604 26472 22094 26500
rect 12115 26404 12572 26432
rect 12115 26401 12127 26404
rect 12069 26395 12127 26401
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 12897 26435 12955 26441
rect 12897 26432 12909 26435
rect 12676 26404 12909 26432
rect 12676 26392 12682 26404
rect 12897 26401 12909 26404
rect 12943 26401 12955 26435
rect 15378 26432 15384 26444
rect 15339 26404 15384 26432
rect 12897 26395 12955 26401
rect 15378 26392 15384 26404
rect 15436 26432 15442 26444
rect 15654 26432 15660 26444
rect 15436 26404 15660 26432
rect 15436 26392 15442 26404
rect 15654 26392 15660 26404
rect 15712 26392 15718 26444
rect 15838 26432 15844 26444
rect 15799 26404 15844 26432
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 16482 26392 16488 26444
rect 16540 26432 16546 26444
rect 17604 26441 17632 26472
rect 17589 26435 17647 26441
rect 17589 26432 17601 26435
rect 16540 26404 17601 26432
rect 16540 26392 16546 26404
rect 17589 26401 17601 26404
rect 17635 26401 17647 26435
rect 18782 26432 18788 26444
rect 18743 26404 18788 26432
rect 17589 26395 17647 26401
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 19426 26432 19432 26444
rect 19387 26404 19432 26432
rect 19426 26392 19432 26404
rect 19484 26392 19490 26444
rect 9861 26367 9919 26373
rect 9861 26364 9873 26367
rect 8496 26336 9873 26364
rect 2130 26256 2136 26308
rect 2188 26296 2194 26308
rect 8496 26305 8524 26336
rect 9861 26333 9873 26336
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 10689 26367 10747 26373
rect 10689 26333 10701 26367
rect 10735 26333 10747 26367
rect 10689 26327 10747 26333
rect 10781 26367 10839 26373
rect 10781 26333 10793 26367
rect 10827 26364 10839 26367
rect 11238 26364 11244 26376
rect 10827 26336 11244 26364
rect 10827 26333 10839 26336
rect 10781 26327 10839 26333
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 20257 26367 20315 26373
rect 20257 26364 20269 26367
rect 19444 26336 20269 26364
rect 8481 26299 8539 26305
rect 8481 26296 8493 26299
rect 2188 26268 8493 26296
rect 2188 26256 2194 26268
rect 8481 26265 8493 26268
rect 8527 26265 8539 26299
rect 8481 26259 8539 26265
rect 9953 26299 10011 26305
rect 9953 26265 9965 26299
rect 9999 26296 10011 26299
rect 11425 26299 11483 26305
rect 11425 26296 11437 26299
rect 9999 26268 11437 26296
rect 9999 26265 10011 26268
rect 9953 26259 10011 26265
rect 11425 26265 11437 26268
rect 11471 26265 11483 26299
rect 11425 26259 11483 26265
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 12618 26296 12624 26308
rect 11572 26268 11617 26296
rect 12579 26268 12624 26296
rect 11572 26256 11578 26268
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 12710 26256 12716 26308
rect 12768 26296 12774 26308
rect 12768 26268 12813 26296
rect 12768 26256 12774 26268
rect 13446 26256 13452 26308
rect 13504 26296 13510 26308
rect 14829 26299 14887 26305
rect 13504 26268 14780 26296
rect 13504 26256 13510 26268
rect 1670 26228 1676 26240
rect 1631 26200 1676 26228
rect 1670 26188 1676 26200
rect 1728 26188 1734 26240
rect 9398 26228 9404 26240
rect 9359 26200 9404 26228
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 14752 26228 14780 26268
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 15194 26296 15200 26308
rect 14875 26268 15200 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 15473 26299 15531 26305
rect 15473 26296 15485 26299
rect 15304 26268 15485 26296
rect 15304 26228 15332 26268
rect 15473 26265 15485 26268
rect 15519 26265 15531 26299
rect 15473 26259 15531 26265
rect 15654 26256 15660 26308
rect 15712 26296 15718 26308
rect 16482 26296 16488 26308
rect 15712 26268 16488 26296
rect 15712 26256 15718 26268
rect 16482 26256 16488 26268
rect 16540 26296 16546 26308
rect 16945 26299 17003 26305
rect 16945 26296 16957 26299
rect 16540 26268 16957 26296
rect 16540 26256 16546 26268
rect 16945 26265 16957 26268
rect 16991 26265 17003 26299
rect 17494 26296 17500 26308
rect 17455 26268 17500 26296
rect 16945 26259 17003 26265
rect 17494 26256 17500 26268
rect 17552 26256 17558 26308
rect 17770 26256 17776 26308
rect 17828 26296 17834 26308
rect 18141 26299 18199 26305
rect 18141 26296 18153 26299
rect 17828 26268 18153 26296
rect 17828 26256 17834 26268
rect 18141 26265 18153 26268
rect 18187 26265 18199 26299
rect 18141 26259 18199 26265
rect 18693 26299 18751 26305
rect 18693 26265 18705 26299
rect 18739 26296 18751 26299
rect 19444 26296 19472 26336
rect 20257 26333 20269 26336
rect 20303 26333 20315 26367
rect 20257 26327 20315 26333
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 20404 26336 20821 26364
rect 20404 26324 20410 26336
rect 20809 26333 20821 26336
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 19610 26296 19616 26308
rect 18739 26268 19472 26296
rect 19571 26268 19616 26296
rect 18739 26265 18751 26268
rect 18693 26259 18751 26265
rect 19610 26256 19616 26268
rect 19668 26256 19674 26308
rect 21361 26299 21419 26305
rect 21361 26296 21373 26299
rect 19720 26268 21373 26296
rect 14752 26200 15332 26228
rect 17678 26188 17684 26240
rect 17736 26228 17742 26240
rect 19720 26228 19748 26268
rect 21361 26265 21373 26268
rect 21407 26265 21419 26299
rect 22066 26296 22094 26472
rect 29181 26367 29239 26373
rect 29181 26333 29193 26367
rect 29227 26364 29239 26367
rect 38102 26364 38108 26376
rect 29227 26336 38108 26364
rect 29227 26333 29239 26336
rect 29181 26327 29239 26333
rect 38102 26324 38108 26336
rect 38160 26324 38166 26376
rect 29089 26299 29147 26305
rect 29089 26296 29101 26299
rect 22066 26268 29101 26296
rect 21361 26259 21419 26265
rect 29089 26265 29101 26268
rect 29135 26265 29147 26299
rect 29089 26259 29147 26265
rect 17736 26200 19748 26228
rect 17736 26188 17742 26200
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 11057 26027 11115 26033
rect 11057 25993 11069 26027
rect 11103 26024 11115 26027
rect 16298 26024 16304 26036
rect 11103 25996 13308 26024
rect 11103 25993 11115 25996
rect 11057 25987 11115 25993
rect 11330 25956 11336 25968
rect 10980 25928 11336 25956
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25888 9367 25891
rect 9398 25888 9404 25900
rect 9355 25860 9404 25888
rect 9355 25857 9367 25860
rect 9309 25851 9367 25857
rect 9398 25848 9404 25860
rect 9456 25888 9462 25900
rect 10980 25897 11008 25928
rect 11330 25916 11336 25928
rect 11388 25916 11394 25968
rect 12618 25956 12624 25968
rect 12579 25928 12624 25956
rect 12618 25916 12624 25928
rect 12676 25916 12682 25968
rect 13280 25965 13308 25996
rect 15304 25996 16304 26024
rect 15304 25965 15332 25996
rect 16298 25984 16304 25996
rect 16356 25984 16362 26036
rect 18322 25984 18328 26036
rect 18380 26024 18386 26036
rect 20165 26027 20223 26033
rect 20165 26024 20177 26027
rect 18380 25996 20177 26024
rect 18380 25984 18386 25996
rect 20165 25993 20177 25996
rect 20211 25993 20223 26027
rect 20898 26024 20904 26036
rect 20859 25996 20904 26024
rect 20165 25987 20223 25993
rect 20898 25984 20904 25996
rect 20956 25984 20962 26036
rect 13265 25959 13323 25965
rect 13265 25925 13277 25959
rect 13311 25925 13323 25959
rect 13265 25919 13323 25925
rect 15289 25959 15347 25965
rect 15289 25925 15301 25959
rect 15335 25925 15347 25959
rect 15289 25919 15347 25925
rect 15746 25916 15752 25968
rect 15804 25956 15810 25968
rect 15841 25959 15899 25965
rect 15841 25956 15853 25959
rect 15804 25928 15853 25956
rect 15804 25916 15810 25928
rect 15841 25925 15853 25928
rect 15887 25925 15899 25959
rect 15841 25919 15899 25925
rect 16574 25916 16580 25968
rect 16632 25956 16638 25968
rect 17589 25959 17647 25965
rect 17589 25956 17601 25959
rect 16632 25928 17601 25956
rect 16632 25916 16638 25928
rect 17589 25925 17601 25928
rect 17635 25925 17647 25959
rect 17589 25919 17647 25925
rect 17954 25916 17960 25968
rect 18012 25956 18018 25968
rect 18233 25959 18291 25965
rect 18233 25956 18245 25959
rect 18012 25928 18245 25956
rect 18012 25916 18018 25928
rect 18233 25925 18245 25928
rect 18279 25925 18291 25959
rect 18233 25919 18291 25925
rect 18785 25959 18843 25965
rect 18785 25925 18797 25959
rect 18831 25956 18843 25959
rect 19518 25956 19524 25968
rect 18831 25928 19524 25956
rect 18831 25925 18843 25928
rect 18785 25919 18843 25925
rect 19518 25916 19524 25928
rect 19576 25916 19582 25968
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 9456 25860 10333 25888
rect 9456 25848 9462 25860
rect 10321 25857 10333 25860
rect 10367 25888 10379 25891
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10367 25860 10977 25888
rect 10367 25857 10379 25860
rect 10321 25851 10379 25857
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 12529 25891 12587 25897
rect 12529 25888 12541 25891
rect 10965 25851 11023 25857
rect 11072 25860 12541 25888
rect 11072 25820 11100 25860
rect 12529 25857 12541 25860
rect 12575 25888 12587 25891
rect 12894 25888 12900 25900
rect 12575 25860 12900 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12894 25848 12900 25860
rect 12952 25848 12958 25900
rect 14458 25848 14464 25900
rect 14516 25888 14522 25900
rect 14645 25891 14703 25897
rect 14645 25888 14657 25891
rect 14516 25860 14657 25888
rect 14516 25848 14522 25860
rect 14645 25857 14657 25860
rect 14691 25857 14703 25891
rect 14645 25851 14703 25857
rect 16850 25848 16856 25900
rect 16908 25888 16914 25900
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16908 25860 17049 25888
rect 16908 25848 16914 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25888 19671 25891
rect 20070 25888 20076 25900
rect 19659 25860 20076 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 20070 25848 20076 25860
rect 20128 25888 20134 25900
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 20128 25860 20269 25888
rect 20128 25848 20134 25860
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25888 20775 25891
rect 21450 25888 21456 25900
rect 20763 25860 21456 25888
rect 20763 25857 20775 25860
rect 20717 25851 20775 25857
rect 21450 25848 21456 25860
rect 21508 25848 21514 25900
rect 9784 25792 11100 25820
rect 11885 25823 11943 25829
rect 9784 25696 9812 25792
rect 11885 25789 11897 25823
rect 11931 25820 11943 25823
rect 13173 25823 13231 25829
rect 13173 25820 13185 25823
rect 11931 25792 13185 25820
rect 11931 25789 11943 25792
rect 11885 25783 11943 25789
rect 13173 25789 13185 25792
rect 13219 25789 13231 25823
rect 13173 25783 13231 25789
rect 13449 25823 13507 25829
rect 13449 25789 13461 25823
rect 13495 25789 13507 25823
rect 13449 25783 13507 25789
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25820 14795 25823
rect 15930 25820 15936 25832
rect 14783 25792 15792 25820
rect 15891 25792 15936 25820
rect 14783 25789 14795 25792
rect 14737 25783 14795 25789
rect 10413 25755 10471 25761
rect 10413 25721 10425 25755
rect 10459 25752 10471 25755
rect 10459 25724 11468 25752
rect 10459 25721 10471 25724
rect 10413 25715 10471 25721
rect 9766 25684 9772 25696
rect 9727 25656 9772 25684
rect 9766 25644 9772 25656
rect 9824 25644 9830 25696
rect 11440 25684 11468 25724
rect 11606 25712 11612 25764
rect 11664 25752 11670 25764
rect 13464 25752 13492 25783
rect 15764 25752 15792 25792
rect 15930 25780 15936 25792
rect 15988 25780 15994 25832
rect 16758 25780 16764 25832
rect 16816 25820 16822 25832
rect 17678 25820 17684 25832
rect 16816 25792 17684 25820
rect 16816 25780 16822 25792
rect 17678 25780 17684 25792
rect 17736 25780 17742 25832
rect 18877 25823 18935 25829
rect 18877 25789 18889 25823
rect 18923 25820 18935 25823
rect 21634 25820 21640 25832
rect 18923 25792 21640 25820
rect 18923 25789 18935 25792
rect 18877 25783 18935 25789
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 17586 25752 17592 25764
rect 11664 25724 13492 25752
rect 13556 25724 14872 25752
rect 15764 25724 17592 25752
rect 11664 25712 11670 25724
rect 12710 25684 12716 25696
rect 11440 25656 12716 25684
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 12894 25644 12900 25696
rect 12952 25684 12958 25696
rect 13556 25684 13584 25724
rect 12952 25656 13584 25684
rect 14844 25684 14872 25724
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 23658 25752 23664 25764
rect 18432 25724 23664 25752
rect 18432 25684 18460 25724
rect 23658 25712 23664 25724
rect 23716 25712 23722 25764
rect 14844 25656 18460 25684
rect 12952 25644 12958 25656
rect 18690 25644 18696 25696
rect 18748 25684 18754 25696
rect 19521 25687 19579 25693
rect 19521 25684 19533 25687
rect 18748 25656 19533 25684
rect 18748 25644 18754 25656
rect 19521 25653 19533 25656
rect 19567 25653 19579 25687
rect 21450 25684 21456 25696
rect 21411 25656 21456 25684
rect 19521 25647 19579 25653
rect 21450 25644 21456 25656
rect 21508 25644 21514 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25480 10839 25483
rect 11514 25480 11520 25492
rect 10827 25452 11520 25480
rect 10827 25449 10839 25452
rect 10781 25443 10839 25449
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 13262 25440 13268 25492
rect 13320 25480 13326 25492
rect 16022 25480 16028 25492
rect 13320 25452 16028 25480
rect 13320 25440 13326 25452
rect 16022 25440 16028 25452
rect 16080 25440 16086 25492
rect 19518 25480 19524 25492
rect 19479 25452 19524 25480
rect 19518 25440 19524 25452
rect 19576 25440 19582 25492
rect 20070 25440 20076 25492
rect 20128 25480 20134 25492
rect 20625 25483 20683 25489
rect 20625 25480 20637 25483
rect 20128 25452 20637 25480
rect 20128 25440 20134 25452
rect 20625 25449 20637 25452
rect 20671 25449 20683 25483
rect 21634 25480 21640 25492
rect 21595 25452 21640 25480
rect 20625 25443 20683 25449
rect 21634 25440 21640 25452
rect 21692 25440 21698 25492
rect 28626 25480 28632 25492
rect 28587 25452 28632 25480
rect 28626 25440 28632 25452
rect 28684 25440 28690 25492
rect 36262 25480 36268 25492
rect 36223 25452 36268 25480
rect 36262 25440 36268 25452
rect 36320 25440 36326 25492
rect 11606 25412 11612 25424
rect 8220 25384 11612 25412
rect 8220 25356 8248 25384
rect 11606 25372 11612 25384
rect 11664 25372 11670 25424
rect 11977 25415 12035 25421
rect 11977 25381 11989 25415
rect 12023 25412 12035 25415
rect 12526 25412 12532 25424
rect 12023 25384 12532 25412
rect 12023 25381 12035 25384
rect 11977 25375 12035 25381
rect 12526 25372 12532 25384
rect 12584 25372 12590 25424
rect 12802 25372 12808 25424
rect 12860 25412 12866 25424
rect 13173 25415 13231 25421
rect 13173 25412 13185 25415
rect 12860 25384 13185 25412
rect 12860 25372 12866 25384
rect 13173 25381 13185 25384
rect 13219 25381 13231 25415
rect 13173 25375 13231 25381
rect 15838 25372 15844 25424
rect 15896 25412 15902 25424
rect 15896 25384 16160 25412
rect 15896 25372 15902 25384
rect 7929 25347 7987 25353
rect 7929 25313 7941 25347
rect 7975 25344 7987 25347
rect 8202 25344 8208 25356
rect 7975 25316 8208 25344
rect 7975 25313 7987 25316
rect 7929 25307 7987 25313
rect 8202 25304 8208 25316
rect 8260 25304 8266 25356
rect 9585 25347 9643 25353
rect 9585 25313 9597 25347
rect 9631 25344 9643 25347
rect 12621 25347 12679 25353
rect 9631 25316 10732 25344
rect 9631 25313 9643 25316
rect 9585 25307 9643 25313
rect 9950 25236 9956 25288
rect 10008 25276 10014 25288
rect 10704 25285 10732 25316
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 13078 25344 13084 25356
rect 12667 25316 13084 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 16132 25353 16160 25384
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25313 16175 25347
rect 18138 25344 18144 25356
rect 18099 25316 18144 25344
rect 16117 25307 16175 25313
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 38010 25344 38016 25356
rect 37971 25316 38016 25344
rect 38010 25304 38016 25316
rect 38068 25304 38074 25356
rect 10045 25279 10103 25285
rect 10045 25276 10057 25279
rect 10008 25248 10057 25276
rect 10008 25236 10014 25248
rect 10045 25245 10057 25248
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10689 25279 10747 25285
rect 10689 25245 10701 25279
rect 10735 25276 10747 25279
rect 11146 25276 11152 25288
rect 10735 25248 11152 25276
rect 10735 25245 10747 25248
rect 10689 25239 10747 25245
rect 5534 25168 5540 25220
rect 5592 25208 5598 25220
rect 7285 25211 7343 25217
rect 7285 25208 7297 25211
rect 5592 25180 7297 25208
rect 5592 25168 5598 25180
rect 7285 25177 7297 25180
rect 7331 25177 7343 25211
rect 7285 25171 7343 25177
rect 7374 25168 7380 25220
rect 7432 25208 7438 25220
rect 7432 25180 7477 25208
rect 7432 25168 7438 25180
rect 10060 25140 10088 25239
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 13964 25248 14473 25276
rect 13964 25236 13970 25248
rect 14461 25245 14473 25248
rect 14507 25245 14519 25279
rect 14461 25239 14519 25245
rect 14918 25236 14924 25288
rect 14976 25276 14982 25288
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 14976 25248 15117 25276
rect 14976 25236 14982 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 17497 25279 17555 25285
rect 17497 25245 17509 25279
rect 17543 25245 17555 25279
rect 17497 25239 17555 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 19886 25276 19892 25288
rect 19659 25248 19892 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 10137 25211 10195 25217
rect 10137 25177 10149 25211
rect 10183 25208 10195 25211
rect 11422 25208 11428 25220
rect 10183 25180 11100 25208
rect 11383 25180 11428 25208
rect 10183 25177 10195 25180
rect 10137 25171 10195 25177
rect 10962 25140 10968 25152
rect 10060 25112 10968 25140
rect 10962 25100 10968 25112
rect 11020 25100 11026 25152
rect 11072 25140 11100 25180
rect 11422 25168 11428 25180
rect 11480 25168 11486 25220
rect 11517 25211 11575 25217
rect 11517 25177 11529 25211
rect 11563 25177 11575 25211
rect 11517 25171 11575 25177
rect 11532 25140 11560 25171
rect 12710 25168 12716 25220
rect 12768 25208 12774 25220
rect 15841 25211 15899 25217
rect 12768 25180 12813 25208
rect 12768 25168 12774 25180
rect 15841 25177 15853 25211
rect 15887 25177 15899 25211
rect 15841 25171 15899 25177
rect 15933 25211 15991 25217
rect 15933 25177 15945 25211
rect 15979 25208 15991 25211
rect 16022 25208 16028 25220
rect 15979 25180 16028 25208
rect 15979 25177 15991 25180
rect 15933 25171 15991 25177
rect 11072 25112 11560 25140
rect 14553 25143 14611 25149
rect 14553 25109 14565 25143
rect 14599 25140 14611 25143
rect 15010 25140 15016 25152
rect 14599 25112 15016 25140
rect 14599 25109 14611 25112
rect 14553 25103 14611 25109
rect 15010 25100 15016 25112
rect 15068 25100 15074 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 15562 25140 15568 25152
rect 15243 25112 15568 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 15856 25140 15884 25171
rect 16022 25168 16028 25180
rect 16080 25168 16086 25220
rect 16666 25168 16672 25220
rect 16724 25208 16730 25220
rect 17512 25208 17540 25239
rect 19886 25236 19892 25248
rect 19944 25236 19950 25288
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20165 25279 20223 25285
rect 20165 25276 20177 25279
rect 20036 25248 20177 25276
rect 20036 25236 20042 25248
rect 20165 25245 20177 25248
rect 20211 25276 20223 25279
rect 21450 25276 21456 25288
rect 20211 25248 21456 25276
rect 20211 25245 20223 25248
rect 20165 25239 20223 25245
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25276 21787 25279
rect 22281 25279 22339 25285
rect 22281 25276 22293 25279
rect 21775 25248 22293 25276
rect 21775 25245 21787 25248
rect 21729 25239 21787 25245
rect 22281 25245 22293 25248
rect 22327 25276 22339 25279
rect 28445 25279 28503 25285
rect 28445 25276 28457 25279
rect 22327 25248 28457 25276
rect 22327 25245 22339 25248
rect 22281 25239 22339 25245
rect 28445 25245 28457 25248
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 18690 25208 18696 25220
rect 16724 25180 17540 25208
rect 18651 25180 18696 25208
rect 16724 25168 16730 25180
rect 18690 25168 18696 25180
rect 18748 25168 18754 25220
rect 18785 25211 18843 25217
rect 18785 25177 18797 25211
rect 18831 25208 18843 25211
rect 19334 25208 19340 25220
rect 18831 25180 19340 25208
rect 18831 25177 18843 25180
rect 18785 25171 18843 25177
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 28460 25208 28488 25239
rect 36262 25236 36268 25288
rect 36320 25276 36326 25288
rect 36817 25279 36875 25285
rect 36817 25276 36829 25279
rect 36320 25248 36829 25276
rect 36320 25236 36326 25248
rect 36817 25245 36829 25248
rect 36863 25245 36875 25279
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 36817 25239 36875 25245
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 29181 25211 29239 25217
rect 29181 25208 29193 25211
rect 28460 25180 29193 25208
rect 29181 25177 29193 25180
rect 29227 25208 29239 25211
rect 37642 25208 37648 25220
rect 29227 25180 37648 25208
rect 29227 25177 29239 25180
rect 29181 25171 29239 25177
rect 37642 25168 37648 25180
rect 37700 25168 37706 25220
rect 16206 25140 16212 25152
rect 15856 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25140 17647 25143
rect 18598 25140 18604 25152
rect 17635 25112 18604 25140
rect 17635 25109 17647 25112
rect 17589 25103 17647 25109
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 36909 25143 36967 25149
rect 36909 25109 36921 25143
rect 36955 25140 36967 25143
rect 38010 25140 38016 25152
rect 36955 25112 38016 25140
rect 36955 25109 36967 25112
rect 36909 25103 36967 25109
rect 38010 25100 38016 25112
rect 38068 25100 38074 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7374 24896 7380 24948
rect 7432 24936 7438 24948
rect 7561 24939 7619 24945
rect 7561 24936 7573 24939
rect 7432 24908 7573 24936
rect 7432 24896 7438 24908
rect 7561 24905 7573 24908
rect 7607 24905 7619 24939
rect 7561 24899 7619 24905
rect 13814 24896 13820 24948
rect 13872 24936 13878 24948
rect 14918 24936 14924 24948
rect 13872 24908 14924 24936
rect 13872 24896 13878 24908
rect 14918 24896 14924 24908
rect 14976 24936 14982 24948
rect 38286 24936 38292 24948
rect 14976 24908 16160 24936
rect 38247 24908 38292 24936
rect 14976 24896 14982 24908
rect 9858 24868 9864 24880
rect 9771 24840 9864 24868
rect 9858 24828 9864 24840
rect 9916 24868 9922 24880
rect 9916 24840 11376 24868
rect 9916 24828 9922 24840
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2130 24800 2136 24812
rect 1903 24772 2136 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2130 24760 2136 24772
rect 2188 24800 2194 24812
rect 2501 24803 2559 24809
rect 2501 24800 2513 24803
rect 2188 24772 2513 24800
rect 2188 24760 2194 24772
rect 2501 24769 2513 24772
rect 2547 24769 2559 24803
rect 2501 24763 2559 24769
rect 7653 24803 7711 24809
rect 7653 24769 7665 24803
rect 7699 24800 7711 24803
rect 9950 24800 9956 24812
rect 7699 24772 9956 24800
rect 7699 24769 7711 24772
rect 7653 24763 7711 24769
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10778 24800 10784 24812
rect 10551 24772 10784 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 11348 24800 11376 24840
rect 11422 24828 11428 24880
rect 11480 24868 11486 24880
rect 11701 24871 11759 24877
rect 11701 24868 11713 24871
rect 11480 24840 11713 24868
rect 11480 24828 11486 24840
rect 11701 24837 11713 24840
rect 11747 24837 11759 24871
rect 13173 24871 13231 24877
rect 13173 24868 13185 24871
rect 11701 24831 11759 24837
rect 12636 24840 13185 24868
rect 11974 24800 11980 24812
rect 11020 24772 11065 24800
rect 11348 24772 11980 24800
rect 11020 24760 11026 24772
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 12636 24800 12664 24840
rect 13173 24837 13185 24840
rect 13219 24837 13231 24871
rect 14642 24868 14648 24880
rect 14603 24840 14648 24868
rect 13173 24831 13231 24837
rect 14642 24828 14648 24840
rect 14700 24828 14706 24880
rect 12406 24772 12664 24800
rect 13817 24803 13875 24809
rect 11057 24735 11115 24741
rect 11057 24701 11069 24735
rect 11103 24732 11115 24735
rect 12406 24732 12434 24772
rect 13817 24769 13829 24803
rect 13863 24800 13875 24803
rect 13906 24800 13912 24812
rect 13863 24772 13912 24800
rect 13863 24769 13875 24772
rect 13817 24763 13875 24769
rect 13906 24760 13912 24772
rect 13964 24760 13970 24812
rect 16132 24809 16160 24908
rect 38286 24896 38292 24908
rect 38344 24896 38350 24948
rect 17405 24871 17463 24877
rect 17405 24868 17417 24871
rect 16868 24840 17417 24868
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16117 24763 16175 24769
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16574 24800 16580 24812
rect 16255 24772 16580 24800
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 12802 24732 12808 24744
rect 11103 24704 12434 24732
rect 12763 24704 12808 24732
rect 11103 24701 11115 24704
rect 11057 24695 11115 24701
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 14274 24732 14280 24744
rect 13311 24704 14280 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 14274 24692 14280 24704
rect 14332 24692 14338 24744
rect 14550 24732 14556 24744
rect 14511 24704 14556 24732
rect 14550 24692 14556 24704
rect 14608 24692 14614 24744
rect 15565 24735 15623 24741
rect 15565 24701 15577 24735
rect 15611 24732 15623 24735
rect 15838 24732 15844 24744
rect 15611 24704 15844 24732
rect 15611 24701 15623 24704
rect 15565 24695 15623 24701
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 16132 24732 16160 24763
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 16666 24732 16672 24744
rect 16132 24704 16672 24732
rect 16666 24692 16672 24704
rect 16724 24692 16730 24744
rect 2041 24667 2099 24673
rect 2041 24633 2053 24667
rect 2087 24664 2099 24667
rect 2314 24664 2320 24676
rect 2087 24636 2320 24664
rect 2087 24633 2099 24636
rect 2041 24627 2099 24633
rect 2314 24624 2320 24636
rect 2372 24624 2378 24676
rect 10413 24667 10471 24673
rect 10413 24633 10425 24667
rect 10459 24664 10471 24667
rect 10459 24636 12434 24664
rect 10459 24633 10471 24636
rect 10413 24627 10471 24633
rect 12406 24596 12434 24636
rect 12710 24624 12716 24676
rect 12768 24664 12774 24676
rect 13814 24664 13820 24676
rect 12768 24636 13820 24664
rect 12768 24624 12774 24636
rect 13814 24624 13820 24636
rect 13872 24624 13878 24676
rect 13909 24667 13967 24673
rect 13909 24633 13921 24667
rect 13955 24664 13967 24667
rect 16868 24664 16896 24840
rect 17405 24837 17417 24840
rect 17451 24837 17463 24871
rect 18138 24868 18144 24880
rect 18099 24840 18144 24868
rect 17405 24831 17463 24837
rect 18138 24828 18144 24840
rect 18196 24828 18202 24880
rect 18598 24828 18604 24880
rect 18656 24868 18662 24880
rect 18693 24871 18751 24877
rect 18693 24868 18705 24871
rect 18656 24840 18705 24868
rect 18656 24828 18662 24840
rect 18693 24837 18705 24840
rect 18739 24837 18751 24871
rect 18693 24831 18751 24837
rect 19334 24828 19340 24880
rect 19392 24868 19398 24880
rect 20073 24871 20131 24877
rect 20073 24868 20085 24871
rect 19392 24840 20085 24868
rect 19392 24828 19398 24840
rect 20073 24837 20085 24840
rect 20119 24837 20131 24871
rect 20073 24831 20131 24837
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24800 19671 24803
rect 19978 24800 19984 24812
rect 19659 24772 19984 24800
rect 19659 24769 19671 24772
rect 19613 24763 19671 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20162 24800 20168 24812
rect 20123 24772 20168 24800
rect 20162 24760 20168 24772
rect 20220 24800 20226 24812
rect 20809 24803 20867 24809
rect 20809 24800 20821 24803
rect 20220 24772 20821 24800
rect 20220 24760 20226 24772
rect 20809 24769 20821 24772
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 17497 24735 17555 24741
rect 17497 24701 17509 24735
rect 17543 24732 17555 24735
rect 17862 24732 17868 24744
rect 17543 24704 17868 24732
rect 17543 24701 17555 24704
rect 17497 24695 17555 24701
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 18785 24735 18843 24741
rect 18785 24701 18797 24735
rect 18831 24732 18843 24735
rect 19337 24735 19395 24741
rect 19337 24732 19349 24735
rect 18831 24704 19349 24732
rect 18831 24701 18843 24704
rect 18785 24695 18843 24701
rect 19337 24701 19349 24704
rect 19383 24701 19395 24735
rect 19337 24695 19395 24701
rect 13955 24636 16896 24664
rect 16945 24667 17003 24673
rect 13955 24633 13967 24636
rect 13909 24627 13967 24633
rect 16945 24633 16957 24667
rect 16991 24633 17003 24667
rect 16945 24627 17003 24633
rect 15102 24596 15108 24608
rect 12406 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 16960 24596 16988 24627
rect 16540 24568 16988 24596
rect 20824 24596 20852 24763
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 32398 24732 32404 24744
rect 21508 24704 32404 24732
rect 21508 24692 21514 24704
rect 32398 24692 32404 24704
rect 32456 24692 32462 24744
rect 28534 24596 28540 24608
rect 20824 24568 28540 24596
rect 16540 24556 16546 24568
rect 28534 24556 28540 24568
rect 28592 24556 28598 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 5077 24395 5135 24401
rect 5077 24361 5089 24395
rect 5123 24392 5135 24395
rect 5534 24392 5540 24404
rect 5123 24364 5540 24392
rect 5123 24361 5135 24364
rect 5077 24355 5135 24361
rect 5534 24352 5540 24364
rect 5592 24352 5598 24404
rect 10870 24352 10876 24404
rect 10928 24392 10934 24404
rect 13078 24392 13084 24404
rect 10928 24364 13084 24392
rect 10928 24352 10934 24364
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 14550 24352 14556 24404
rect 14608 24392 14614 24404
rect 14645 24395 14703 24401
rect 14645 24392 14657 24395
rect 14608 24364 14657 24392
rect 14608 24352 14614 24364
rect 14645 24361 14657 24364
rect 14691 24361 14703 24395
rect 14645 24355 14703 24361
rect 15102 24352 15108 24404
rect 15160 24392 15166 24404
rect 17954 24392 17960 24404
rect 15160 24364 17960 24392
rect 15160 24352 15166 24364
rect 17954 24352 17960 24364
rect 18012 24352 18018 24404
rect 18877 24395 18935 24401
rect 18877 24361 18889 24395
rect 18923 24392 18935 24395
rect 20070 24392 20076 24404
rect 18923 24364 20076 24392
rect 18923 24361 18935 24364
rect 18877 24355 18935 24361
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 26878 24392 26884 24404
rect 26839 24364 26884 24392
rect 26878 24352 26884 24364
rect 26936 24352 26942 24404
rect 19429 24327 19487 24333
rect 19429 24324 19441 24327
rect 2746 24296 19441 24324
rect 2038 24216 2044 24268
rect 2096 24256 2102 24268
rect 2746 24256 2774 24296
rect 19429 24293 19441 24296
rect 19475 24293 19487 24327
rect 19429 24287 19487 24293
rect 2096 24228 2774 24256
rect 12437 24259 12495 24265
rect 2096 24216 2102 24228
rect 12437 24225 12449 24259
rect 12483 24256 12495 24259
rect 13725 24259 13783 24265
rect 12483 24228 12940 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 1854 24188 1860 24200
rect 1815 24160 1860 24188
rect 1854 24148 1860 24160
rect 1912 24148 1918 24200
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4672 24160 4997 24188
rect 4672 24148 4678 24160
rect 4985 24157 4997 24160
rect 5031 24188 5043 24191
rect 5629 24191 5687 24197
rect 5629 24188 5641 24191
rect 5031 24160 5641 24188
rect 5031 24157 5043 24160
rect 4985 24151 5043 24157
rect 5629 24157 5641 24160
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 10597 24191 10655 24197
rect 10597 24188 10609 24191
rect 9088 24160 10609 24188
rect 9088 24148 9094 24160
rect 10597 24157 10609 24160
rect 10643 24157 10655 24191
rect 12342 24188 12348 24200
rect 12303 24160 12348 24188
rect 10597 24151 10655 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 10689 24123 10747 24129
rect 10689 24089 10701 24123
rect 10735 24120 10747 24123
rect 12802 24120 12808 24132
rect 10735 24092 12808 24120
rect 10735 24089 10747 24092
rect 10689 24083 10747 24089
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 1670 24052 1676 24064
rect 1631 24024 1676 24052
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 11330 24052 11336 24064
rect 11291 24024 11336 24052
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11885 24055 11943 24061
rect 11885 24021 11897 24055
rect 11931 24052 11943 24055
rect 12710 24052 12716 24064
rect 11931 24024 12716 24052
rect 11931 24021 11943 24024
rect 11885 24015 11943 24021
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 12912 24052 12940 24228
rect 13725 24225 13737 24259
rect 13771 24256 13783 24259
rect 15102 24256 15108 24268
rect 13771 24228 15108 24256
rect 13771 24225 13783 24228
rect 13725 24219 13783 24225
rect 15102 24216 15108 24228
rect 15160 24216 15166 24268
rect 15194 24216 15200 24268
rect 15252 24256 15258 24268
rect 15933 24259 15991 24265
rect 15933 24256 15945 24259
rect 15252 24228 15945 24256
rect 15252 24216 15258 24228
rect 15933 24225 15945 24228
rect 15979 24225 15991 24259
rect 15933 24219 15991 24225
rect 16206 24216 16212 24268
rect 16264 24256 16270 24268
rect 16577 24259 16635 24265
rect 16577 24256 16589 24259
rect 16264 24228 16589 24256
rect 16264 24216 16270 24228
rect 16577 24225 16589 24228
rect 16623 24256 16635 24259
rect 17770 24256 17776 24268
rect 16623 24228 17776 24256
rect 16623 24225 16635 24228
rect 16577 24219 16635 24225
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 14182 24148 14188 24200
rect 14240 24190 14246 24200
rect 14277 24191 14335 24197
rect 14277 24190 14289 24191
rect 14240 24162 14289 24190
rect 14240 24148 14246 24162
rect 14277 24157 14289 24162
rect 14323 24157 14335 24191
rect 14458 24188 14464 24200
rect 14419 24160 14464 24188
rect 14277 24151 14335 24157
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 15010 24148 15016 24200
rect 15068 24188 15074 24200
rect 15068 24160 15792 24188
rect 15068 24148 15074 24160
rect 13078 24120 13084 24132
rect 13039 24092 13084 24120
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 13170 24080 13176 24132
rect 13228 24120 13234 24132
rect 15764 24120 15792 24160
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16724 24160 17049 24188
rect 16724 24148 16730 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 26697 24191 26755 24197
rect 19659 24160 20116 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 16002 24123 16060 24129
rect 16002 24120 16014 24123
rect 13228 24092 13273 24120
rect 15764 24092 16014 24120
rect 13228 24080 13234 24092
rect 16002 24089 16014 24092
rect 16048 24089 16060 24123
rect 16002 24083 16060 24089
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 18141 24123 18199 24129
rect 18141 24120 18153 24123
rect 17828 24092 18153 24120
rect 17828 24080 17834 24092
rect 18141 24089 18153 24092
rect 18187 24089 18199 24123
rect 18141 24083 18199 24089
rect 18233 24123 18291 24129
rect 18233 24089 18245 24123
rect 18279 24120 18291 24123
rect 19334 24120 19340 24132
rect 18279 24092 19340 24120
rect 18279 24089 18291 24092
rect 18233 24083 18291 24089
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 20088 24064 20116 24160
rect 26697 24157 26709 24191
rect 26743 24188 26755 24191
rect 26743 24160 27476 24188
rect 26743 24157 26755 24160
rect 26697 24151 26755 24157
rect 14458 24052 14464 24064
rect 12912 24024 14464 24052
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 20070 24052 20076 24064
rect 20031 24024 20076 24052
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 27448 24061 27476 24160
rect 27433 24055 27491 24061
rect 27433 24021 27445 24055
rect 27479 24052 27491 24055
rect 27522 24052 27528 24064
rect 27479 24024 27528 24052
rect 27479 24021 27491 24024
rect 27433 24015 27491 24021
rect 27522 24012 27528 24024
rect 27580 24012 27586 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 11793 23851 11851 23857
rect 11793 23817 11805 23851
rect 11839 23848 11851 23851
rect 12342 23848 12348 23860
rect 11839 23820 12348 23848
rect 11839 23817 11851 23820
rect 11793 23811 11851 23817
rect 12342 23808 12348 23820
rect 12400 23848 12406 23860
rect 12805 23851 12863 23857
rect 12805 23848 12817 23851
rect 12400 23820 12817 23848
rect 12400 23808 12406 23820
rect 12805 23817 12817 23820
rect 12851 23817 12863 23851
rect 14182 23848 14188 23860
rect 14143 23820 14188 23848
rect 12805 23811 12863 23817
rect 12820 23780 12848 23811
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14829 23851 14887 23857
rect 14829 23817 14841 23851
rect 14875 23848 14887 23851
rect 17770 23848 17776 23860
rect 14875 23820 17776 23848
rect 14875 23817 14887 23820
rect 14829 23811 14887 23817
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 19334 23848 19340 23860
rect 17880 23820 18276 23848
rect 19295 23820 19340 23848
rect 15562 23780 15568 23792
rect 12820 23752 14780 23780
rect 15523 23752 15568 23780
rect 10410 23672 10416 23724
rect 10468 23712 10474 23724
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 10468 23684 12265 23712
rect 10468 23672 10474 23684
rect 12253 23681 12265 23684
rect 12299 23712 12311 23715
rect 13357 23715 13415 23721
rect 13357 23712 13369 23715
rect 12299 23684 13369 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 13357 23681 13369 23684
rect 13403 23712 13415 23715
rect 13403 23684 14136 23712
rect 13403 23681 13415 23684
rect 13357 23675 13415 23681
rect 14108 23644 14136 23684
rect 14182 23672 14188 23724
rect 14240 23712 14246 23724
rect 14642 23712 14648 23724
rect 14240 23684 14648 23712
rect 14240 23672 14246 23684
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 14752 23721 14780 23752
rect 15562 23740 15568 23752
rect 15620 23740 15626 23792
rect 16114 23780 16120 23792
rect 16075 23752 16120 23780
rect 16114 23740 16120 23752
rect 16172 23740 16178 23792
rect 17034 23780 17040 23792
rect 16995 23752 17040 23780
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 17586 23740 17592 23792
rect 17644 23780 17650 23792
rect 17880 23780 17908 23820
rect 18248 23789 18276 23820
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 18141 23783 18199 23789
rect 18141 23780 18153 23783
rect 17644 23752 17908 23780
rect 17972 23752 18153 23780
rect 17644 23740 17650 23752
rect 14737 23715 14795 23721
rect 14737 23681 14749 23715
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 17862 23672 17868 23724
rect 17920 23712 17926 23724
rect 17972 23712 18000 23752
rect 18141 23749 18153 23752
rect 18187 23749 18199 23783
rect 18141 23743 18199 23749
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23749 18291 23783
rect 18233 23743 18291 23749
rect 17920 23684 18000 23712
rect 19521 23715 19579 23721
rect 17920 23672 17926 23684
rect 19521 23681 19533 23715
rect 19567 23712 19579 23715
rect 20070 23712 20076 23724
rect 19567 23684 20076 23712
rect 19567 23681 19579 23684
rect 19521 23675 19579 23681
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 38010 23712 38016 23724
rect 37971 23684 38016 23712
rect 38010 23672 38016 23684
rect 38068 23672 38074 23724
rect 15473 23647 15531 23653
rect 14108 23616 15424 23644
rect 13449 23579 13507 23585
rect 13449 23545 13461 23579
rect 13495 23576 13507 23579
rect 15286 23576 15292 23588
rect 13495 23548 15292 23576
rect 13495 23545 13507 23548
rect 13449 23539 13507 23545
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 15396 23576 15424 23616
rect 15473 23613 15485 23647
rect 15519 23644 15531 23647
rect 15562 23644 15568 23656
rect 15519 23616 15568 23644
rect 15519 23613 15531 23616
rect 15473 23607 15531 23613
rect 15562 23604 15568 23616
rect 15620 23604 15626 23656
rect 16942 23644 16948 23656
rect 16903 23616 16948 23644
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 18064 23616 18429 23644
rect 18064 23588 18092 23616
rect 18417 23613 18429 23616
rect 18463 23613 18475 23647
rect 18417 23607 18475 23613
rect 17497 23579 17555 23585
rect 15396 23548 16804 23576
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 16666 23508 16672 23520
rect 12860 23480 16672 23508
rect 12860 23468 12866 23480
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 16776 23508 16804 23548
rect 17497 23545 17509 23579
rect 17543 23576 17555 23579
rect 18046 23576 18052 23588
rect 17543 23548 18052 23576
rect 17543 23545 17555 23548
rect 17497 23539 17555 23545
rect 18046 23536 18052 23548
rect 18104 23536 18110 23588
rect 20346 23576 20352 23588
rect 19904 23548 20352 23576
rect 19904 23508 19932 23548
rect 20346 23536 20352 23548
rect 20404 23536 20410 23588
rect 20070 23508 20076 23520
rect 16776 23480 19932 23508
rect 20031 23480 20076 23508
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 27522 23468 27528 23520
rect 27580 23508 27586 23520
rect 29822 23508 29828 23520
rect 27580 23480 29828 23508
rect 27580 23468 27586 23480
rect 29822 23468 29828 23480
rect 29880 23468 29886 23520
rect 38194 23508 38200 23520
rect 38155 23480 38200 23508
rect 38194 23468 38200 23480
rect 38252 23468 38258 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 1949 23307 2007 23313
rect 1949 23304 1961 23307
rect 1912 23276 1961 23304
rect 1912 23264 1918 23276
rect 1949 23273 1961 23276
rect 1995 23273 2007 23307
rect 1949 23267 2007 23273
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13541 23307 13599 23313
rect 13541 23304 13553 23307
rect 13228 23276 13553 23304
rect 13228 23264 13234 23276
rect 13541 23273 13553 23276
rect 13587 23273 13599 23307
rect 13541 23267 13599 23273
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 14829 23307 14887 23313
rect 14829 23304 14841 23307
rect 14608 23276 14841 23304
rect 14608 23264 14614 23276
rect 14829 23273 14841 23276
rect 14875 23273 14887 23307
rect 14829 23267 14887 23273
rect 11238 23196 11244 23248
rect 11296 23236 11302 23248
rect 11296 23208 14964 23236
rect 11296 23196 11302 23208
rect 12894 23128 12900 23180
rect 12952 23168 12958 23180
rect 12989 23171 13047 23177
rect 12989 23168 13001 23171
rect 12952 23140 13001 23168
rect 12952 23128 12958 23140
rect 12989 23137 13001 23140
rect 13035 23168 13047 23171
rect 14182 23168 14188 23180
rect 13035 23140 14188 23168
rect 13035 23137 13047 23140
rect 12989 23131 13047 23137
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23168 14427 23171
rect 14826 23168 14832 23180
rect 14415 23140 14832 23168
rect 14415 23137 14427 23140
rect 14369 23131 14427 23137
rect 14826 23128 14832 23140
rect 14884 23128 14890 23180
rect 2133 23103 2191 23109
rect 2133 23069 2145 23103
rect 2179 23100 2191 23103
rect 12437 23103 12495 23109
rect 2179 23072 2728 23100
rect 2179 23069 2191 23072
rect 2133 23063 2191 23069
rect 2700 22973 2728 23072
rect 12437 23069 12449 23103
rect 12483 23100 12495 23103
rect 13633 23103 13691 23109
rect 13633 23100 13645 23103
rect 12483 23072 13645 23100
rect 12483 23069 12495 23072
rect 12437 23063 12495 23069
rect 13633 23069 13645 23072
rect 13679 23100 13691 23103
rect 13998 23100 14004 23112
rect 13679 23072 14004 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 2685 22967 2743 22973
rect 2685 22933 2697 22967
rect 2731 22964 2743 22967
rect 4614 22964 4620 22976
rect 2731 22936 4620 22964
rect 2731 22933 2743 22936
rect 2685 22927 2743 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 14936 22964 14964 23208
rect 16022 23196 16028 23248
rect 16080 23236 16086 23248
rect 17589 23239 17647 23245
rect 17589 23236 17601 23239
rect 16080 23208 17601 23236
rect 16080 23196 16086 23208
rect 17589 23205 17601 23208
rect 17635 23205 17647 23239
rect 17589 23199 17647 23205
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23168 15531 23171
rect 16390 23168 16396 23180
rect 15519 23140 16396 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 16390 23128 16396 23140
rect 16448 23168 16454 23180
rect 16942 23168 16948 23180
rect 16448 23140 16948 23168
rect 16448 23128 16454 23140
rect 16942 23128 16948 23140
rect 17000 23128 17006 23180
rect 18322 23060 18328 23112
rect 18380 23100 18386 23112
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 18380 23072 19901 23100
rect 18380 23060 18386 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23100 20131 23103
rect 23382 23100 23388 23112
rect 20119 23072 23388 23100
rect 20119 23069 20131 23072
rect 20073 23063 20131 23069
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 16022 23032 16028 23044
rect 15252 23004 16028 23032
rect 15252 22992 15258 23004
rect 16022 22992 16028 23004
rect 16080 22992 16086 23044
rect 16117 23035 16175 23041
rect 16117 23001 16129 23035
rect 16163 23001 16175 23035
rect 17034 23032 17040 23044
rect 16995 23004 17040 23032
rect 16117 22995 16175 23001
rect 16132 22964 16160 22995
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 18046 23032 18052 23044
rect 18007 23004 18052 23032
rect 18046 22992 18052 23004
rect 18104 22992 18110 23044
rect 18141 23035 18199 23041
rect 18141 23001 18153 23035
rect 18187 23032 18199 23035
rect 28902 23032 28908 23044
rect 18187 23004 28908 23032
rect 18187 23001 18199 23004
rect 18141 22995 18199 23001
rect 28902 22992 28908 23004
rect 28960 22992 28966 23044
rect 14936 22936 16160 22964
rect 17678 22924 17684 22976
rect 17736 22964 17742 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 17736 22936 18705 22964
rect 17736 22924 17742 22936
rect 18693 22933 18705 22936
rect 18739 22933 18751 22967
rect 18693 22927 18751 22933
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 18840 22936 19441 22964
rect 18840 22924 18846 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 13173 22763 13231 22769
rect 13173 22760 13185 22763
rect 11388 22732 13185 22760
rect 11388 22720 11394 22732
rect 13173 22729 13185 22732
rect 13219 22760 13231 22763
rect 13725 22763 13783 22769
rect 13725 22760 13737 22763
rect 13219 22732 13737 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13725 22729 13737 22732
rect 13771 22760 13783 22763
rect 13906 22760 13912 22772
rect 13771 22732 13912 22760
rect 13771 22729 13783 22732
rect 13725 22723 13783 22729
rect 13906 22720 13912 22732
rect 13964 22720 13970 22772
rect 15930 22720 15936 22772
rect 15988 22760 15994 22772
rect 16117 22763 16175 22769
rect 16117 22760 16129 22763
rect 15988 22732 16129 22760
rect 15988 22720 15994 22732
rect 16117 22729 16129 22732
rect 16163 22729 16175 22763
rect 16117 22723 16175 22729
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 18322 22760 18328 22772
rect 17267 22732 18328 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 23382 22760 23388 22772
rect 23343 22732 23388 22760
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 24029 22763 24087 22769
rect 24029 22729 24041 22763
rect 24075 22760 24087 22763
rect 27522 22760 27528 22772
rect 24075 22732 27528 22760
rect 24075 22729 24087 22732
rect 24029 22723 24087 22729
rect 13924 22624 13952 22720
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 14918 22692 14924 22704
rect 14332 22664 14924 22692
rect 14332 22652 14338 22664
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 15013 22695 15071 22701
rect 15013 22661 15025 22695
rect 15059 22692 15071 22695
rect 15378 22692 15384 22704
rect 15059 22664 15384 22692
rect 15059 22661 15071 22664
rect 15013 22655 15071 22661
rect 15378 22652 15384 22664
rect 15436 22652 15442 22704
rect 17954 22692 17960 22704
rect 17915 22664 17960 22692
rect 17954 22652 17960 22664
rect 18012 22652 18018 22704
rect 14185 22627 14243 22633
rect 14185 22624 14197 22627
rect 13924 22596 14197 22624
rect 14185 22593 14197 22596
rect 14231 22593 14243 22627
rect 16206 22624 16212 22636
rect 16167 22596 16212 22624
rect 14185 22587 14243 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 16316 22596 17141 22624
rect 15194 22556 15200 22568
rect 15155 22528 15200 22556
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 13998 22448 14004 22500
rect 14056 22488 14062 22500
rect 16316 22488 16344 22596
rect 17129 22593 17141 22596
rect 17175 22624 17187 22627
rect 17678 22624 17684 22636
rect 17175 22596 17684 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17678 22584 17684 22596
rect 17736 22584 17742 22636
rect 23477 22627 23535 22633
rect 23477 22593 23489 22627
rect 23523 22624 23535 22627
rect 24044 22624 24072 22723
rect 27522 22720 27528 22732
rect 27580 22720 27586 22772
rect 23523 22596 24072 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22556 17923 22559
rect 17954 22556 17960 22568
rect 17911 22528 17960 22556
rect 17911 22525 17923 22528
rect 17865 22519 17923 22525
rect 17954 22516 17960 22528
rect 18012 22556 18018 22568
rect 18782 22556 18788 22568
rect 18012 22528 18788 22556
rect 18012 22516 18018 22528
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22525 18935 22559
rect 18877 22519 18935 22525
rect 14056 22460 16344 22488
rect 14056 22448 14062 22460
rect 17034 22448 17040 22500
rect 17092 22488 17098 22500
rect 17678 22488 17684 22500
rect 17092 22460 17684 22488
rect 17092 22448 17098 22460
rect 17678 22448 17684 22460
rect 17736 22488 17742 22500
rect 18892 22488 18920 22519
rect 17736 22460 18920 22488
rect 17736 22448 17742 22460
rect 14274 22420 14280 22432
rect 14235 22392 14280 22420
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 14550 22176 14556 22228
rect 14608 22216 14614 22228
rect 15013 22219 15071 22225
rect 15013 22216 15025 22219
rect 14608 22188 15025 22216
rect 14608 22176 14614 22188
rect 15013 22185 15025 22188
rect 15059 22185 15071 22219
rect 15013 22179 15071 22185
rect 18046 22176 18052 22228
rect 18104 22216 18110 22228
rect 18141 22219 18199 22225
rect 18141 22216 18153 22219
rect 18104 22188 18153 22216
rect 18104 22176 18110 22188
rect 18141 22185 18153 22188
rect 18187 22185 18199 22219
rect 18141 22179 18199 22185
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 14829 22083 14887 22089
rect 14829 22080 14841 22083
rect 14332 22052 14841 22080
rect 14332 22040 14338 22052
rect 14829 22049 14841 22052
rect 14875 22049 14887 22083
rect 14829 22043 14887 22049
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 16942 22080 16948 22092
rect 16623 22052 16948 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 25314 22080 25320 22092
rect 18156 22052 25320 22080
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 14550 22012 14556 22024
rect 1903 21984 14556 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 22012 14703 22015
rect 14918 22012 14924 22024
rect 14691 21984 14924 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15841 21947 15899 21953
rect 15841 21913 15853 21947
rect 15887 21913 15899 21947
rect 15841 21907 15899 21913
rect 1670 21876 1676 21888
rect 1631 21848 1676 21876
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 13725 21879 13783 21885
rect 13725 21845 13737 21879
rect 13771 21876 13783 21879
rect 14458 21876 14464 21888
rect 13771 21848 14464 21876
rect 13771 21845 13783 21848
rect 13725 21839 13783 21845
rect 14458 21836 14464 21848
rect 14516 21876 14522 21888
rect 15856 21876 15884 21907
rect 16666 21904 16672 21956
rect 16724 21944 16730 21956
rect 17589 21947 17647 21953
rect 16724 21916 16769 21944
rect 16724 21904 16730 21916
rect 17589 21913 17601 21947
rect 17635 21944 17647 21947
rect 17678 21944 17684 21956
rect 17635 21916 17684 21944
rect 17635 21913 17647 21916
rect 17589 21907 17647 21913
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 14516 21848 15884 21876
rect 15933 21879 15991 21885
rect 14516 21836 14522 21848
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 18156 21876 18184 22052
rect 25314 22040 25320 22052
rect 25372 22040 25378 22092
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 22012 18291 22015
rect 37921 22015 37979 22021
rect 18279 21984 18736 22012
rect 18279 21981 18291 21984
rect 18233 21975 18291 21981
rect 18708 21888 18736 21984
rect 37921 21981 37933 22015
rect 37967 22012 37979 22015
rect 38286 22012 38292 22024
rect 37967 21984 38292 22012
rect 37967 21981 37979 21984
rect 37921 21975 37979 21981
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 18690 21876 18696 21888
rect 15979 21848 18184 21876
rect 18651 21848 18696 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 37734 21876 37740 21888
rect 37695 21848 37740 21876
rect 37734 21836 37740 21848
rect 37792 21836 37798 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 14185 21675 14243 21681
rect 14185 21641 14197 21675
rect 14231 21672 14243 21675
rect 14366 21672 14372 21684
rect 14231 21644 14372 21672
rect 14231 21641 14243 21644
rect 14185 21635 14243 21641
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 14550 21632 14556 21684
rect 14608 21672 14614 21684
rect 14645 21675 14703 21681
rect 14645 21672 14657 21675
rect 14608 21644 14657 21672
rect 14608 21632 14614 21644
rect 14645 21641 14657 21644
rect 14691 21641 14703 21675
rect 15378 21672 15384 21684
rect 15339 21644 15384 21672
rect 14645 21635 14703 21641
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18049 21675 18107 21681
rect 18049 21672 18061 21675
rect 18012 21644 18061 21672
rect 18012 21632 18018 21644
rect 18049 21641 18061 21644
rect 18095 21641 18107 21675
rect 18049 21635 18107 21641
rect 14384 21604 14412 21632
rect 15102 21604 15108 21616
rect 14384 21576 15108 21604
rect 15102 21564 15108 21576
rect 15160 21604 15166 21616
rect 15160 21576 15516 21604
rect 15160 21564 15166 21576
rect 15488 21545 15516 21576
rect 13633 21539 13691 21545
rect 13633 21505 13645 21539
rect 13679 21536 13691 21539
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 13679 21508 14841 21536
rect 13679 21505 13691 21508
rect 13633 21499 13691 21505
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 18690 21536 18696 21548
rect 18651 21508 18696 21536
rect 15473 21499 15531 21505
rect 14844 21400 14872 21499
rect 18690 21496 18696 21508
rect 18748 21536 18754 21548
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 18748 21508 19165 21536
rect 18748 21496 18754 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 19153 21499 19211 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 16301 21471 16359 21477
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16574 21468 16580 21480
rect 16347 21440 16580 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 17402 21468 17408 21480
rect 17363 21440 17408 21468
rect 17402 21428 17408 21440
rect 17460 21428 17466 21480
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21468 17647 21471
rect 17770 21468 17776 21480
rect 17635 21440 17776 21468
rect 17635 21437 17647 21440
rect 17589 21431 17647 21437
rect 17770 21428 17776 21440
rect 17828 21428 17834 21480
rect 16206 21400 16212 21412
rect 14844 21372 16212 21400
rect 16206 21360 16212 21372
rect 16264 21400 16270 21412
rect 16945 21403 17003 21409
rect 16945 21400 16957 21403
rect 16264 21372 16957 21400
rect 16264 21360 16270 21372
rect 16945 21369 16957 21372
rect 16991 21400 17003 21403
rect 37918 21400 37924 21412
rect 16991 21372 37924 21400
rect 16991 21369 17003 21372
rect 16945 21363 17003 21369
rect 37918 21360 37924 21372
rect 37976 21360 37982 21412
rect 18598 21332 18604 21344
rect 18559 21304 18604 21332
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 13906 21088 13912 21140
rect 13964 21128 13970 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 13964 21100 14289 21128
rect 13964 21088 13970 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 14918 21128 14924 21140
rect 14879 21100 14924 21128
rect 14277 21091 14335 21097
rect 14292 20992 14320 21091
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 16942 21128 16948 21140
rect 16903 21100 16948 21128
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17770 21128 17776 21140
rect 17731 21100 17776 21128
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 14292 20964 16160 20992
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 16132 20933 16160 20964
rect 16574 20952 16580 21004
rect 16632 20992 16638 21004
rect 16761 20995 16819 21001
rect 16632 20964 16677 20992
rect 16632 20952 16638 20964
rect 16761 20961 16773 20995
rect 16807 20992 16819 20995
rect 18598 20992 18604 21004
rect 16807 20964 18604 20992
rect 16807 20961 16819 20964
rect 16761 20955 16819 20961
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 15013 20927 15071 20933
rect 15013 20924 15025 20927
rect 14516 20896 15025 20924
rect 14516 20884 14522 20896
rect 15013 20893 15025 20896
rect 15059 20893 15071 20927
rect 15013 20887 15071 20893
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 17865 20927 17923 20933
rect 17865 20924 17877 20927
rect 16117 20887 16175 20893
rect 16546 20896 17877 20924
rect 1578 20816 1584 20868
rect 1636 20856 1642 20868
rect 1673 20859 1731 20865
rect 1673 20856 1685 20859
rect 1636 20828 1685 20856
rect 1636 20816 1642 20828
rect 1673 20825 1685 20828
rect 1719 20825 1731 20859
rect 1673 20819 1731 20825
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 16546 20856 16574 20896
rect 17865 20893 17877 20896
rect 17911 20924 17923 20927
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 17911 20896 18337 20924
rect 17911 20893 17923 20896
rect 17865 20887 17923 20893
rect 18325 20893 18337 20896
rect 18371 20924 18383 20927
rect 18690 20924 18696 20936
rect 18371 20896 18696 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 12032 20828 16574 20856
rect 12032 20816 12038 20828
rect 1765 20791 1823 20797
rect 1765 20757 1777 20791
rect 1811 20788 1823 20791
rect 11698 20788 11704 20800
rect 1811 20760 11704 20788
rect 1811 20757 1823 20760
rect 1765 20751 1823 20757
rect 11698 20748 11704 20760
rect 11756 20748 11762 20800
rect 16022 20788 16028 20800
rect 15983 20760 16028 20788
rect 16022 20748 16028 20760
rect 16080 20748 16086 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 15102 20544 15108 20596
rect 15160 20584 15166 20596
rect 15197 20587 15255 20593
rect 15197 20584 15209 20587
rect 15160 20556 15209 20584
rect 15160 20544 15166 20556
rect 15197 20553 15209 20556
rect 15243 20553 15255 20587
rect 15197 20547 15255 20553
rect 16301 20587 16359 20593
rect 16301 20553 16313 20587
rect 16347 20584 16359 20587
rect 16942 20584 16948 20596
rect 16347 20556 16948 20584
rect 16347 20553 16359 20556
rect 16301 20547 16359 20553
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17402 20544 17408 20596
rect 17460 20584 17466 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17460 20556 17601 20584
rect 17460 20544 17466 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 28902 20544 28908 20596
rect 28960 20584 28966 20596
rect 30101 20587 30159 20593
rect 30101 20584 30113 20587
rect 28960 20556 30113 20584
rect 28960 20544 28966 20556
rect 30101 20553 30113 20556
rect 30147 20553 30159 20587
rect 38010 20584 38016 20596
rect 37971 20556 38016 20584
rect 30101 20547 30159 20553
rect 38010 20544 38016 20556
rect 38068 20544 38074 20596
rect 1578 20516 1584 20528
rect 1539 20488 1584 20516
rect 1578 20476 1584 20488
rect 1636 20476 1642 20528
rect 11698 20476 11704 20528
rect 11756 20516 11762 20528
rect 11756 20488 17724 20516
rect 11756 20476 11762 20488
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15841 20451 15899 20457
rect 15160 20420 15792 20448
rect 15160 20408 15166 20420
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15344 20352 15669 20380
rect 15344 20340 15350 20352
rect 15657 20349 15669 20352
rect 15703 20349 15715 20383
rect 15764 20380 15792 20420
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16022 20448 16028 20460
rect 15887 20420 16028 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16546 20420 17049 20448
rect 16546 20380 16574 20420
rect 17037 20417 17049 20420
rect 17083 20448 17095 20451
rect 17126 20448 17132 20460
rect 17083 20420 17132 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17696 20457 17724 20488
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 30193 20451 30251 20457
rect 17727 20420 18276 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 15764 20352 16574 20380
rect 15657 20343 15715 20349
rect 14458 20204 14464 20256
rect 14516 20244 14522 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14516 20216 14565 20244
rect 14516 20204 14522 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 18248 20253 18276 20420
rect 30193 20417 30205 20451
rect 30239 20448 30251 20451
rect 37826 20448 37832 20460
rect 30239 20420 37832 20448
rect 30239 20417 30251 20420
rect 30193 20411 30251 20417
rect 37826 20408 37832 20420
rect 37884 20408 37890 20460
rect 16945 20247 17003 20253
rect 16945 20244 16957 20247
rect 16632 20216 16957 20244
rect 16632 20204 16638 20216
rect 16945 20213 16957 20216
rect 16991 20213 17003 20247
rect 16945 20207 17003 20213
rect 18233 20247 18291 20253
rect 18233 20213 18245 20247
rect 18279 20244 18291 20247
rect 18782 20244 18788 20256
rect 18279 20216 18788 20244
rect 18279 20213 18291 20216
rect 18233 20207 18291 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 15470 20000 15476 20052
rect 15528 20040 15534 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15528 20012 15669 20040
rect 15528 20000 15534 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 15657 20003 15715 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17589 20043 17647 20049
rect 17589 20009 17601 20043
rect 17635 20040 17647 20043
rect 17862 20040 17868 20052
rect 17635 20012 17868 20040
rect 17635 20009 17647 20012
rect 17589 20003 17647 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 16632 19876 16677 19904
rect 16632 19864 16638 19876
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15212 19808 15761 19836
rect 15212 19712 15240 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 16393 19839 16451 19845
rect 16393 19805 16405 19839
rect 16439 19836 16451 19839
rect 16482 19836 16488 19848
rect 16439 19808 16488 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 17681 19799 17739 19805
rect 17696 19712 17724 19799
rect 15105 19703 15163 19709
rect 15105 19669 15117 19703
rect 15151 19700 15163 19703
rect 15194 19700 15200 19712
rect 15151 19672 15200 19700
rect 15151 19669 15163 19672
rect 15105 19663 15163 19669
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17736 19672 18153 19700
rect 17736 19660 17742 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 15286 19496 15292 19508
rect 15247 19468 15292 19496
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 17954 19496 17960 19508
rect 17915 19468 17960 19496
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 17678 19388 17684 19440
rect 17736 19428 17742 19440
rect 24578 19428 24584 19440
rect 17736 19400 24584 19428
rect 17736 19388 17742 19400
rect 24578 19388 24584 19400
rect 24636 19388 24642 19440
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 14608 19332 15209 19360
rect 14608 19320 14614 19332
rect 15197 19329 15209 19332
rect 15243 19360 15255 19363
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15243 19332 15945 19360
rect 15243 19329 15255 19332
rect 15197 19323 15255 19329
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 17126 19360 17132 19372
rect 17087 19332 17132 19360
rect 15933 19323 15991 19329
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 18601 19363 18659 19369
rect 17267 19332 18460 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 18432 19301 18460 19332
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 19426 19360 19432 19372
rect 18647 19332 19432 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 37553 19363 37611 19369
rect 37553 19329 37565 19363
rect 37599 19360 37611 19363
rect 38194 19360 38200 19372
rect 37599 19332 38200 19360
rect 37599 19329 37611 19332
rect 37553 19323 37611 19329
rect 38194 19320 38200 19332
rect 38252 19320 38258 19372
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 37918 19252 37924 19304
rect 37976 19292 37982 19304
rect 38013 19295 38071 19301
rect 38013 19292 38025 19295
rect 37976 19264 38025 19292
rect 37976 19252 37982 19264
rect 38013 19261 38025 19264
rect 38059 19261 38071 19295
rect 38013 19255 38071 19261
rect 16117 19227 16175 19233
rect 16117 19193 16129 19227
rect 16163 19224 16175 19227
rect 16163 19196 26234 19224
rect 16163 19193 16175 19196
rect 16117 19187 16175 19193
rect 26206 19156 26234 19196
rect 37734 19156 37740 19168
rect 26206 19128 37740 19156
rect 37734 19116 37740 19128
rect 37792 19116 37798 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 17037 18955 17095 18961
rect 17037 18921 17049 18955
rect 17083 18952 17095 18955
rect 17126 18952 17132 18964
rect 17083 18924 17132 18952
rect 17083 18921 17095 18924
rect 17037 18915 17095 18921
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 6181 18751 6239 18757
rect 6181 18717 6193 18751
rect 6227 18748 6239 18751
rect 9122 18748 9128 18760
rect 6227 18720 9128 18748
rect 6227 18717 6239 18720
rect 6181 18711 6239 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 1578 18640 1584 18692
rect 1636 18680 1642 18692
rect 1673 18683 1731 18689
rect 1673 18680 1685 18683
rect 1636 18652 1685 18680
rect 1636 18640 1642 18652
rect 1673 18649 1685 18652
rect 1719 18649 1731 18683
rect 1673 18643 1731 18649
rect 1857 18683 1915 18689
rect 1857 18649 1869 18683
rect 1903 18680 1915 18683
rect 9766 18680 9772 18692
rect 1903 18652 9772 18680
rect 1903 18649 1915 18652
rect 1857 18643 1915 18649
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 6089 18615 6147 18621
rect 6089 18612 6101 18615
rect 2832 18584 6101 18612
rect 2832 18572 2838 18584
rect 6089 18581 6101 18584
rect 6135 18581 6147 18615
rect 6089 18575 6147 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19484 17836 19717 17864
rect 19484 17824 19490 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 19843 17632 20392 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 20364 17536 20392 17632
rect 20346 17524 20352 17536
rect 20307 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 20346 17184 20352 17196
rect 20259 17156 20352 17184
rect 20346 17144 20352 17156
rect 20404 17184 20410 17196
rect 20404 17156 21036 17184
rect 20404 17144 20410 17156
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 21008 16989 21036 17156
rect 20257 16983 20315 16989
rect 20257 16980 20269 16983
rect 13044 16952 20269 16980
rect 13044 16940 13050 16952
rect 20257 16949 20269 16952
rect 20303 16949 20315 16983
rect 20257 16943 20315 16949
rect 20993 16983 21051 16989
rect 20993 16949 21005 16983
rect 21039 16980 21051 16983
rect 38010 16980 38016 16992
rect 21039 16952 38016 16980
rect 21039 16949 21051 16952
rect 20993 16943 21051 16949
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 14645 16575 14703 16581
rect 1903 16544 14504 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 14476 16445 14504 16544
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 14691 16544 15148 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 15120 16445 15148 16544
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16405 14519 16439
rect 14461 16399 14519 16405
rect 15105 16439 15163 16445
rect 15105 16405 15117 16439
rect 15151 16436 15163 16439
rect 15194 16436 15200 16448
rect 15151 16408 15200 16436
rect 15151 16405 15163 16408
rect 15105 16399 15163 16405
rect 15194 16396 15200 16408
rect 15252 16436 15258 16448
rect 15378 16436 15384 16448
rect 15252 16408 15384 16436
rect 15252 16396 15258 16408
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 10870 16164 10876 16176
rect 10643 16136 10876 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 10870 16124 10876 16136
rect 10928 16164 10934 16176
rect 12894 16164 12900 16176
rect 10928 16136 12900 16164
rect 10928 16124 10934 16136
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 9858 16096 9864 16108
rect 9819 16068 9864 16096
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12250 16096 12256 16108
rect 12207 16068 12256 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12250 16056 12256 16068
rect 12308 16096 12314 16108
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12308 16068 12633 16096
rect 12308 16056 12314 16068
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 13722 16056 13728 16108
rect 13780 16096 13786 16108
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 13780 16068 19809 16096
rect 13780 16056 13786 16068
rect 19797 16065 19809 16068
rect 19843 16096 19855 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19843 16068 20453 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 23198 16056 23204 16108
rect 23256 16096 23262 16108
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 23256 16068 37473 16096
rect 23256 16056 23262 16068
rect 37461 16065 37473 16068
rect 37507 16096 37519 16099
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 37507 16068 38025 16096
rect 37507 16065 37519 16068
rect 37461 16059 37519 16065
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 9456 15932 11989 15960
rect 9456 15920 9462 15932
rect 11977 15929 11989 15932
rect 12023 15929 12035 15963
rect 11977 15923 12035 15929
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 33686 15960 33692 15972
rect 15436 15932 33692 15960
rect 15436 15920 15442 15932
rect 33686 15920 33692 15932
rect 33744 15920 33750 15972
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 7524 15864 9689 15892
rect 7524 15852 7530 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 10502 15892 10508 15904
rect 10463 15864 10508 15892
rect 9677 15855 9735 15861
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 19978 15892 19984 15904
rect 19939 15864 19984 15892
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 9398 15688 9404 15700
rect 1912 15660 9404 15688
rect 1912 15648 1918 15660
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9916 15660 9965 15688
rect 9916 15648 9922 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 9953 15651 10011 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 16117 15691 16175 15697
rect 16117 15657 16129 15691
rect 16163 15688 16175 15691
rect 16390 15688 16396 15700
rect 16163 15660 16396 15688
rect 16163 15657 16175 15660
rect 16117 15651 16175 15657
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15484 16267 15487
rect 16390 15484 16396 15496
rect 16255 15456 16396 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16390 15444 16396 15456
rect 16448 15484 16454 15496
rect 16448 15456 16574 15484
rect 16448 15444 16454 15456
rect 16546 15348 16574 15456
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16546 15320 16681 15348
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1670 14328 1676 14340
rect 1631 14300 1676 14328
rect 1670 14288 1676 14300
rect 1728 14288 1734 14340
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14260 1823 14263
rect 17678 14260 17684 14272
rect 1811 14232 17684 14260
rect 1811 14229 1823 14232
rect 1765 14223 1823 14229
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 37826 13880 37832 13932
rect 37884 13920 37890 13932
rect 38013 13923 38071 13929
rect 38013 13920 38025 13923
rect 37884 13892 38025 13920
rect 37884 13880 37890 13892
rect 38013 13889 38025 13892
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 38286 13852 38292 13864
rect 38247 13824 38292 13852
rect 38286 13812 38292 13824
rect 38344 13812 38350 13864
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 38286 13512 38292 13524
rect 38247 13484 38292 13512
rect 38286 13472 38292 13484
rect 38344 13472 38350 13524
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 2774 13308 2780 13320
rect 1903 13280 2780 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 38194 11744 38200 11756
rect 37599 11716 38200 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 38013 11611 38071 11617
rect 38013 11608 38025 11611
rect 26206 11580 38025 11608
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 26206 11540 26234 11580
rect 38013 11577 38025 11580
rect 38059 11577 38071 11611
rect 38013 11571 38071 11577
rect 20128 11512 26234 11540
rect 20128 11500 20134 11512
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 16482 11336 16488 11348
rect 16443 11308 16488 11336
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 20438 11200 20444 11212
rect 2455 11172 20444 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2424 11132 2452 11163
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 1903 11104 2452 11132
rect 16577 11135 16635 11141
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 16577 11101 16589 11135
rect 16623 11132 16635 11135
rect 16623 11104 17172 11132
rect 16623 11101 16635 11104
rect 16577 11095 16635 11101
rect 17144 11076 17172 11104
rect 17126 11064 17132 11076
rect 17087 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 15010 10792 15016 10804
rect 14971 10764 15016 10792
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 17218 10792 17224 10804
rect 17179 10764 17224 10792
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 18782 10792 18788 10804
rect 18743 10764 18788 10792
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15654 10656 15660 10668
rect 15151 10628 15660 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 17313 10659 17371 10665
rect 17313 10625 17325 10659
rect 17359 10656 17371 10659
rect 17402 10656 17408 10668
rect 17359 10628 17408 10656
rect 17359 10625 17371 10628
rect 17313 10619 17371 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18800 10656 18828 10752
rect 18187 10628 18828 10656
rect 37553 10659 37611 10665
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 37553 10625 37565 10659
rect 37599 10656 37611 10659
rect 38194 10656 38200 10668
rect 37599 10628 38200 10656
rect 37599 10625 37611 10628
rect 37553 10619 37611 10625
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 38013 10523 38071 10529
rect 38013 10520 38025 10523
rect 16448 10492 38025 10520
rect 16448 10480 16454 10492
rect 38013 10489 38025 10492
rect 38059 10489 38071 10523
rect 38013 10483 38071 10489
rect 15654 10452 15660 10464
rect 15615 10424 15660 10452
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 16390 10248 16396 10260
rect 15151 10220 16396 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10044 14611 10047
rect 15120 10044 15148 10211
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 14599 10016 15148 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 14366 9908 14372 9920
rect 14327 9880 14372 9908
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 17402 9908 17408 9920
rect 17363 9880 17408 9908
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16816 9608 16957 9636
rect 16816 9596 16822 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17494 9568 17500 9580
rect 17083 9540 17500 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 14366 8956 14372 8968
rect 1903 8928 14372 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 24578 8956 24584 8968
rect 24539 8928 24584 8956
rect 24578 8916 24584 8928
rect 24636 8956 24642 8968
rect 25225 8959 25283 8965
rect 25225 8956 25237 8959
rect 24636 8928 25237 8956
rect 24636 8916 24642 8928
rect 25225 8925 25237 8928
rect 25271 8925 25283 8959
rect 25225 8919 25283 8925
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 24762 8820 24768 8832
rect 24723 8792 24768 8820
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 38102 8616 38108 8628
rect 38063 8588 38108 8616
rect 38102 8576 38108 8588
rect 38160 8576 38166 8628
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8480 37703 8483
rect 38286 8480 38292 8492
rect 37691 8452 38292 8480
rect 37691 8449 37703 8452
rect 37645 8443 37703 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 23198 8004 23204 8016
rect 23159 7976 23204 8004
rect 23198 7964 23204 7976
rect 23256 7964 23262 8016
rect 10594 7760 10600 7812
rect 10652 7800 10658 7812
rect 23017 7803 23075 7809
rect 23017 7800 23029 7803
rect 10652 7772 23029 7800
rect 10652 7760 10658 7772
rect 23017 7769 23029 7772
rect 23063 7769 23075 7803
rect 23017 7763 23075 7769
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 14458 7188 14464 7200
rect 1811 7160 14464 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 38010 6372 38016 6384
rect 37971 6344 38016 6372
rect 38010 6332 38016 6344
rect 38068 6332 38074 6384
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6304 37611 6307
rect 38194 6304 38200 6316
rect 37599 6276 38200 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 38194 6264 38200 6276
rect 38252 6264 38258 6316
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5692 1918 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 1912 5664 2329 5692
rect 1912 5652 1918 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 37642 4700 37648 4752
rect 37700 4740 37706 4752
rect 38013 4743 38071 4749
rect 38013 4740 38025 4743
rect 37700 4712 38025 4740
rect 37700 4700 37706 4712
rect 38013 4709 38025 4712
rect 38059 4709 38071 4743
rect 38013 4703 38071 4709
rect 37553 4539 37611 4545
rect 37553 4505 37565 4539
rect 37599 4536 37611 4539
rect 38194 4536 38200 4548
rect 37599 4508 38200 4536
rect 37599 4505 37611 4508
rect 37553 4499 37611 4505
rect 38194 4496 38200 4508
rect 38252 4496 38258 4548
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 12802 3516 12808 3528
rect 1903 3488 12808 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 36722 3516 36728 3528
rect 26206 3488 36728 3516
rect 15654 3408 15660 3460
rect 15712 3448 15718 3460
rect 16022 3448 16028 3460
rect 15712 3420 16028 3448
rect 15712 3408 15718 3420
rect 16022 3408 16028 3420
rect 16080 3448 16086 3460
rect 21358 3448 21364 3460
rect 16080 3420 21364 3448
rect 16080 3408 16086 3420
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 23750 3408 23756 3460
rect 23808 3448 23814 3460
rect 26206 3448 26234 3488
rect 36722 3476 36728 3488
rect 36780 3476 36786 3528
rect 38013 3451 38071 3457
rect 38013 3448 38025 3451
rect 23808 3420 26234 3448
rect 35866 3420 38025 3448
rect 23808 3408 23814 3420
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17494 3380 17500 3392
rect 17276 3352 17500 3380
rect 17276 3340 17282 3352
rect 17494 3340 17500 3352
rect 17552 3380 17558 3392
rect 35866 3380 35894 3420
rect 38013 3417 38025 3420
rect 38059 3417 38071 3451
rect 38013 3411 38071 3417
rect 38197 3451 38255 3457
rect 38197 3417 38209 3451
rect 38243 3448 38255 3451
rect 38654 3448 38660 3460
rect 38243 3420 38660 3448
rect 38243 3417 38255 3420
rect 38197 3411 38255 3417
rect 17552 3352 35894 3380
rect 37553 3383 37611 3389
rect 17552 3340 17558 3352
rect 37553 3349 37565 3383
rect 37599 3380 37611 3383
rect 38212 3380 38240 3411
rect 38654 3408 38660 3420
rect 38712 3408 38718 3460
rect 37599 3352 38240 3380
rect 37599 3349 37611 3352
rect 37553 3343 37611 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5592 3148 5733 3176
rect 5592 3136 5598 3148
rect 5721 3145 5733 3148
rect 5767 3176 5779 3179
rect 19426 3176 19432 3188
rect 5767 3148 19432 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 37461 3179 37519 3185
rect 37461 3176 37473 3179
rect 24820 3148 37473 3176
rect 24820 3136 24826 3148
rect 37461 3145 37473 3148
rect 37507 3145 37519 3179
rect 37461 3139 37519 3145
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16356 3080 19196 3108
rect 16356 3068 16362 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 1903 3012 12940 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 12802 2904 12808 2916
rect 12763 2876 12808 2904
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 12912 2904 12940 3012
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 14550 3040 14556 3052
rect 13044 3012 13089 3040
rect 14511 3012 14556 3040
rect 13044 3000 13050 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15795 3012 16221 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 16209 3009 16221 3012
rect 16255 3040 16267 3043
rect 17402 3040 17408 3052
rect 16255 3012 16574 3040
rect 17315 3012 17408 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 14182 2972 14188 2984
rect 13863 2944 14188 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 14182 2932 14188 2944
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 16546 2972 16574 3012
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 19168 3049 19196 3080
rect 21358 3068 21364 3120
rect 21416 3108 21422 3120
rect 21416 3080 26234 3108
rect 21416 3068 21422 3080
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19199 3012 19809 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 23750 3040 23756 3052
rect 23711 3012 23756 3040
rect 19797 3003 19855 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24857 3043 24915 3049
rect 24857 3009 24869 3043
rect 24903 3040 24915 3043
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 24903 3012 25513 3040
rect 24903 3009 24915 3012
rect 24857 3003 24915 3009
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 26206 3040 26234 3080
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26206 3012 27169 3040
rect 25501 3003 25559 3009
rect 27157 3009 27169 3012
rect 27203 3040 27215 3043
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 27203 3012 27813 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 37476 3040 37504 3139
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37476 3012 38025 3040
rect 27801 3003 27859 3009
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 17218 2972 17224 2984
rect 16546 2944 17224 2972
rect 14277 2935 14335 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 12912 2876 15577 2904
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 17420 2904 17448 3000
rect 17862 2932 17868 2984
rect 17920 2972 17926 2984
rect 24872 2972 24900 3003
rect 31018 2972 31024 2984
rect 17920 2944 24900 2972
rect 24964 2944 31024 2972
rect 17920 2932 17926 2944
rect 18141 2907 18199 2913
rect 18141 2904 18153 2907
rect 17420 2876 18153 2904
rect 15565 2867 15623 2873
rect 18141 2873 18153 2876
rect 18187 2904 18199 2907
rect 24964 2904 24992 2944
rect 31018 2932 31024 2944
rect 31076 2932 31082 2984
rect 18187 2876 24992 2904
rect 27341 2907 27399 2913
rect 18187 2873 18199 2876
rect 18141 2867 18199 2873
rect 27341 2873 27353 2907
rect 27387 2904 27399 2907
rect 34422 2904 34428 2916
rect 27387 2876 34428 2904
rect 27387 2873 27399 2876
rect 27341 2867 27399 2873
rect 34422 2864 34428 2876
rect 34480 2864 34486 2916
rect 36909 2907 36967 2913
rect 36909 2873 36921 2907
rect 36955 2904 36967 2907
rect 38102 2904 38108 2916
rect 36955 2876 38108 2904
rect 36955 2873 36967 2876
rect 36909 2867 36967 2873
rect 38102 2864 38108 2876
rect 38160 2864 38166 2916
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 2774 2836 2780 2848
rect 2687 2808 2780 2836
rect 2774 2796 2780 2808
rect 2832 2836 2838 2848
rect 10502 2836 10508 2848
rect 2832 2808 10508 2836
rect 2832 2796 2838 2808
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17552 2808 17601 2836
rect 17552 2796 17558 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 17589 2799 17647 2805
rect 19245 2839 19303 2845
rect 19245 2805 19257 2839
rect 19291 2836 19303 2839
rect 19702 2836 19708 2848
rect 19291 2808 19708 2836
rect 19291 2805 19303 2808
rect 19245 2799 19303 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 23566 2836 23572 2848
rect 23527 2808 23572 2836
rect 23566 2796 23572 2808
rect 23624 2796 23630 2848
rect 24949 2839 25007 2845
rect 24949 2805 24961 2839
rect 24995 2836 25007 2839
rect 27154 2836 27160 2848
rect 24995 2808 27160 2836
rect 24995 2805 25007 2808
rect 24949 2799 25007 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 29638 2836 29644 2848
rect 29599 2808 29644 2836
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 10594 2632 10600 2644
rect 10555 2604 10600 2632
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 13173 2635 13231 2641
rect 13173 2632 13185 2635
rect 13044 2604 13185 2632
rect 13044 2592 13050 2604
rect 13173 2601 13185 2604
rect 13219 2632 13231 2635
rect 17126 2632 17132 2644
rect 13219 2604 17132 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 17126 2592 17132 2604
rect 17184 2632 17190 2644
rect 28534 2632 28540 2644
rect 17184 2604 24900 2632
rect 28495 2604 28540 2632
rect 17184 2592 17190 2604
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 23566 2564 23572 2576
rect 2409 2527 2467 2533
rect 12636 2536 23572 2564
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 8904 2468 9413 2496
rect 8904 2456 8910 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2314 2428 2320 2440
rect 1903 2400 2320 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2774 2428 2780 2440
rect 2639 2400 2780 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3344 2400 3985 2428
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 3973 2391 4031 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8496 2400 9137 2428
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5224 2264 5365 2292
rect 5224 2252 5230 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8496 2301 8524 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 12636 2437 12664 2536
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 15528 2468 16313 2496
rect 15528 2456 15534 2468
rect 16301 2465 16313 2468
rect 16347 2496 16359 2499
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 16347 2468 16865 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 24872 2505 24900 2604
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 29822 2632 29828 2644
rect 29783 2604 29828 2632
rect 29822 2592 29828 2604
rect 29880 2592 29886 2644
rect 32398 2632 32404 2644
rect 32359 2604 32404 2632
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33686 2632 33692 2644
rect 33647 2604 33692 2632
rect 33686 2592 33692 2604
rect 33744 2592 33750 2644
rect 36722 2632 36728 2644
rect 36683 2604 36728 2632
rect 36722 2592 36728 2604
rect 36780 2592 36786 2644
rect 31018 2524 31024 2576
rect 31076 2564 31082 2576
rect 38013 2567 38071 2573
rect 38013 2564 38025 2567
rect 31076 2536 38025 2564
rect 31076 2524 31082 2536
rect 38013 2533 38025 2536
rect 38059 2533 38071 2567
rect 38013 2527 38071 2533
rect 24857 2499 24915 2505
rect 20036 2468 22784 2496
rect 20036 2456 20042 2468
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10376 2400 10425 2428
rect 10376 2388 10382 2400
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 10459 2400 11069 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 12621 2391 12679 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18322 2388 18328 2440
rect 18380 2428 18386 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18380 2400 19441 2428
rect 18380 2388 18386 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 22756 2437 22784 2468
rect 24857 2465 24869 2499
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 19760 2400 22017 2428
rect 19760 2388 19766 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22741 2431 22799 2437
rect 22741 2397 22753 2431
rect 22787 2397 22799 2431
rect 22741 2391 22799 2397
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2428 24087 2431
rect 24486 2428 24492 2440
rect 24075 2400 24492 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 24486 2388 24492 2400
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 27154 2428 27160 2440
rect 27115 2400 27160 2428
rect 24581 2391 24639 2397
rect 27154 2388 27160 2400
rect 27212 2388 27218 2440
rect 34422 2388 34428 2440
rect 34480 2428 34486 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 34480 2400 35541 2428
rect 34480 2388 34486 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 36909 2431 36967 2437
rect 36909 2428 36921 2431
rect 36780 2400 36921 2428
rect 36780 2388 36786 2400
rect 36909 2397 36921 2400
rect 36955 2428 36967 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36955 2400 37473 2428
rect 36955 2397 36967 2400
rect 36909 2391 36967 2397
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 27985 2363 28043 2369
rect 27985 2329 27997 2363
rect 28031 2360 28043 2363
rect 28350 2360 28356 2372
rect 28031 2332 28356 2360
rect 28031 2329 28043 2332
rect 27985 2323 28043 2329
rect 28350 2320 28356 2332
rect 28408 2360 28414 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28408 2332 28641 2360
rect 28408 2320 28414 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 29638 2320 29644 2372
rect 29696 2360 29702 2372
rect 29917 2363 29975 2369
rect 29917 2360 29929 2363
rect 29696 2332 29929 2360
rect 29696 2320 29702 2332
rect 29917 2329 29929 2332
rect 29963 2329 29975 2363
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 29917 2323 29975 2329
rect 31772 2332 32505 2360
rect 31772 2304 31800 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 33137 2363 33195 2369
rect 33137 2329 33149 2363
rect 33183 2360 33195 2363
rect 33502 2360 33508 2372
rect 33183 2332 33508 2360
rect 33183 2329 33195 2332
rect 33137 2323 33195 2329
rect 33502 2320 33508 2332
rect 33560 2360 33566 2372
rect 33781 2363 33839 2369
rect 33781 2360 33793 2363
rect 33560 2332 33793 2360
rect 33560 2320 33566 2332
rect 33781 2329 33793 2332
rect 33827 2329 33839 2363
rect 38194 2360 38200 2372
rect 38155 2332 38200 2360
rect 33781 2323 33839 2329
rect 38194 2320 38200 2332
rect 38252 2320 38258 2372
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12308 2264 12449 2292
rect 12308 2252 12314 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21324 2264 22201 2292
rect 21324 2252 21330 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 22612 2264 22937 2292
rect 22612 2252 22618 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 26476 2264 27353 2292
rect 26476 2252 26482 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 31754 2292 31760 2304
rect 31715 2264 31760 2292
rect 27341 2255 27399 2261
rect 31754 2252 31760 2264
rect 31812 2252 31818 2304
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35713 2295 35771 2301
rect 35713 2292 35725 2295
rect 35492 2264 35725 2292
rect 35492 2252 35498 2264
rect 35713 2261 35725 2264
rect 35759 2261 35771 2295
rect 35713 2255 35771 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7288 37408 7340 37460
rect 10140 37408 10192 37460
rect 10876 37408 10928 37460
rect 16764 37408 16816 37460
rect 18052 37408 18104 37460
rect 20352 37340 20404 37392
rect 4528 37272 4580 37324
rect 5632 37272 5684 37324
rect 3884 37204 3936 37256
rect 6000 37247 6052 37256
rect 6000 37213 6009 37247
rect 6009 37213 6043 37247
rect 6043 37213 6052 37247
rect 10508 37272 10560 37324
rect 11060 37272 11112 37324
rect 12072 37272 12124 37324
rect 6000 37204 6052 37213
rect 2504 37136 2556 37188
rect 3148 37136 3200 37188
rect 5448 37136 5500 37188
rect 7196 37204 7248 37256
rect 8576 37247 8628 37256
rect 8576 37213 8585 37247
rect 8585 37213 8619 37247
rect 8619 37213 8628 37247
rect 8576 37204 8628 37213
rect 8760 37204 8812 37256
rect 11520 37204 11572 37256
rect 7012 37136 7064 37188
rect 1492 37068 1544 37120
rect 5816 37068 5868 37120
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 10600 37136 10652 37188
rect 12992 37204 13044 37256
rect 14832 37204 14884 37256
rect 18144 37315 18196 37324
rect 18144 37281 18153 37315
rect 18153 37281 18187 37315
rect 18187 37281 18196 37315
rect 18144 37272 18196 37281
rect 16764 37204 16816 37256
rect 18052 37204 18104 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 20904 37204 20956 37256
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 26884 37204 26936 37256
rect 28632 37204 28684 37256
rect 30932 37204 30984 37256
rect 32496 37204 32548 37256
rect 34796 37204 34848 37256
rect 10784 37068 10836 37120
rect 15200 37136 15252 37188
rect 38016 37204 38068 37256
rect 37740 37136 37792 37188
rect 12808 37068 12860 37120
rect 12900 37068 12952 37120
rect 14924 37111 14976 37120
rect 14924 37077 14933 37111
rect 14933 37077 14967 37111
rect 14967 37077 14976 37111
rect 14924 37068 14976 37077
rect 16948 37111 17000 37120
rect 16948 37077 16957 37111
rect 16957 37077 16991 37111
rect 16991 37077 17000 37111
rect 16948 37068 17000 37077
rect 19984 37068 20036 37120
rect 22100 37068 22152 37120
rect 23848 37068 23900 37120
rect 25136 37068 25188 37120
rect 27068 37068 27120 37120
rect 29000 37068 29052 37120
rect 31024 37111 31076 37120
rect 31024 37077 31033 37111
rect 31033 37077 31067 37111
rect 31067 37077 31076 37111
rect 31024 37068 31076 37077
rect 32220 37068 32272 37120
rect 34520 37068 34572 37120
rect 36084 37068 36136 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 3884 36864 3936 36916
rect 4896 36864 4948 36916
rect 6000 36864 6052 36916
rect 8576 36864 8628 36916
rect 5816 36839 5868 36848
rect 1584 36771 1636 36780
rect 1584 36737 1593 36771
rect 1593 36737 1627 36771
rect 1627 36737 1636 36771
rect 1584 36728 1636 36737
rect 4896 36771 4948 36780
rect 4896 36737 4905 36771
rect 4905 36737 4939 36771
rect 4939 36737 4948 36771
rect 5816 36805 5825 36839
rect 5825 36805 5859 36839
rect 5859 36805 5868 36839
rect 5816 36796 5868 36805
rect 6184 36796 6236 36848
rect 9220 36796 9272 36848
rect 10600 36796 10652 36848
rect 10784 36864 10836 36916
rect 20076 36864 20128 36916
rect 32496 36907 32548 36916
rect 32496 36873 32505 36907
rect 32505 36873 32539 36907
rect 32539 36873 32548 36907
rect 32496 36864 32548 36873
rect 39304 36864 39356 36916
rect 4896 36728 4948 36737
rect 5724 36728 5776 36780
rect 11060 36796 11112 36848
rect 11520 36728 11572 36780
rect 13084 36728 13136 36780
rect 14924 36728 14976 36780
rect 15200 36728 15252 36780
rect 16488 36728 16540 36780
rect 31024 36728 31076 36780
rect 2136 36660 2188 36712
rect 3608 36660 3660 36712
rect 5540 36660 5592 36712
rect 6552 36703 6604 36712
rect 6552 36669 6561 36703
rect 6561 36669 6595 36703
rect 6595 36669 6604 36703
rect 6552 36660 6604 36669
rect 7012 36660 7064 36712
rect 8300 36703 8352 36712
rect 8300 36669 8309 36703
rect 8309 36669 8343 36703
rect 8343 36669 8352 36703
rect 8300 36660 8352 36669
rect 8576 36703 8628 36712
rect 8576 36669 8585 36703
rect 8585 36669 8619 36703
rect 8619 36669 8628 36703
rect 8576 36660 8628 36669
rect 8668 36660 8720 36712
rect 9312 36660 9364 36712
rect 10508 36660 10560 36712
rect 6460 36592 6512 36644
rect 7196 36524 7248 36576
rect 13544 36660 13596 36712
rect 27896 36703 27948 36712
rect 27896 36669 27905 36703
rect 27905 36669 27939 36703
rect 27939 36669 27948 36703
rect 27896 36660 27948 36669
rect 16028 36592 16080 36644
rect 37924 36728 37976 36780
rect 10968 36524 11020 36576
rect 13176 36524 13228 36576
rect 14096 36567 14148 36576
rect 14096 36533 14105 36567
rect 14105 36533 14139 36567
rect 14139 36533 14148 36567
rect 14096 36524 14148 36533
rect 15292 36567 15344 36576
rect 15292 36533 15301 36567
rect 15301 36533 15335 36567
rect 15335 36533 15344 36567
rect 15292 36524 15344 36533
rect 15936 36524 15988 36576
rect 25320 36524 25372 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2596 36320 2648 36372
rect 3884 36184 3936 36236
rect 3056 36116 3108 36168
rect 14096 36320 14148 36372
rect 15936 36320 15988 36372
rect 1952 36091 2004 36100
rect 1952 36057 1961 36091
rect 1961 36057 1995 36091
rect 1995 36057 2004 36091
rect 1952 36048 2004 36057
rect 5080 36048 5132 36100
rect 5448 36252 5500 36304
rect 8300 36252 8352 36304
rect 9588 36252 9640 36304
rect 10968 36252 11020 36304
rect 12072 36295 12124 36304
rect 12072 36261 12081 36295
rect 12081 36261 12115 36295
rect 12115 36261 12124 36295
rect 12072 36252 12124 36261
rect 13176 36295 13228 36304
rect 13176 36261 13185 36295
rect 13185 36261 13219 36295
rect 13219 36261 13228 36295
rect 13176 36252 13228 36261
rect 14004 36252 14056 36304
rect 5448 36116 5500 36168
rect 6828 36159 6880 36168
rect 6828 36125 6837 36159
rect 6837 36125 6871 36159
rect 6871 36125 6880 36159
rect 6828 36116 6880 36125
rect 7748 36116 7800 36168
rect 6644 36048 6696 36100
rect 11520 36227 11572 36236
rect 11520 36193 11529 36227
rect 11529 36193 11563 36227
rect 11563 36193 11572 36227
rect 11520 36184 11572 36193
rect 15292 36184 15344 36236
rect 8484 36116 8536 36168
rect 9220 36116 9272 36168
rect 9496 36116 9548 36168
rect 10968 36116 11020 36168
rect 27896 36252 27948 36304
rect 5540 35980 5592 36032
rect 7932 35980 7984 36032
rect 9220 35980 9272 36032
rect 11704 36048 11756 36100
rect 12808 36048 12860 36100
rect 16856 36048 16908 36100
rect 38200 36091 38252 36100
rect 38200 36057 38209 36091
rect 38209 36057 38243 36091
rect 38243 36057 38252 36091
rect 38200 36048 38252 36057
rect 10876 35980 10928 36032
rect 38108 36023 38160 36032
rect 38108 35989 38117 36023
rect 38117 35989 38151 36023
rect 38151 35989 38160 36023
rect 38108 35980 38160 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4068 35776 4120 35828
rect 1952 35751 2004 35760
rect 1952 35717 1961 35751
rect 1961 35717 1995 35751
rect 1995 35717 2004 35751
rect 1952 35708 2004 35717
rect 2228 35708 2280 35760
rect 6000 35708 6052 35760
rect 6092 35708 6144 35760
rect 3976 35683 4028 35692
rect 3976 35649 3985 35683
rect 3985 35649 4019 35683
rect 4019 35649 4028 35683
rect 3976 35640 4028 35649
rect 5540 35640 5592 35692
rect 9588 35708 9640 35760
rect 15936 35776 15988 35828
rect 24584 35776 24636 35828
rect 38292 35776 38344 35828
rect 14464 35751 14516 35760
rect 14464 35717 14473 35751
rect 14473 35717 14507 35751
rect 14507 35717 14516 35751
rect 14464 35708 14516 35717
rect 9956 35640 10008 35692
rect 12348 35681 12400 35692
rect 12348 35647 12357 35681
rect 12357 35647 12391 35681
rect 12391 35647 12400 35681
rect 23112 35683 23164 35692
rect 12348 35640 12400 35647
rect 23112 35649 23121 35683
rect 23121 35649 23155 35683
rect 23155 35649 23164 35683
rect 23112 35640 23164 35649
rect 37556 35640 37608 35692
rect 6828 35572 6880 35624
rect 7288 35615 7340 35624
rect 7288 35581 7297 35615
rect 7297 35581 7331 35615
rect 7331 35581 7340 35615
rect 7288 35572 7340 35581
rect 8208 35572 8260 35624
rect 8392 35572 8444 35624
rect 9036 35615 9088 35624
rect 9036 35581 9045 35615
rect 9045 35581 9079 35615
rect 9079 35581 9088 35615
rect 9036 35572 9088 35581
rect 4620 35504 4672 35556
rect 4712 35436 4764 35488
rect 5908 35479 5960 35488
rect 5908 35445 5917 35479
rect 5917 35445 5951 35479
rect 5951 35445 5960 35479
rect 5908 35436 5960 35445
rect 9680 35504 9732 35556
rect 16304 35572 16356 35624
rect 10784 35504 10836 35556
rect 14372 35504 14424 35556
rect 13452 35479 13504 35488
rect 13452 35445 13461 35479
rect 13461 35445 13495 35479
rect 13495 35445 13504 35479
rect 13452 35436 13504 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 664 35232 716 35284
rect 3884 35096 3936 35148
rect 5632 35096 5684 35148
rect 7748 35232 7800 35284
rect 10968 35232 11020 35284
rect 13452 35232 13504 35284
rect 15936 35232 15988 35284
rect 6828 35096 6880 35148
rect 8300 35096 8352 35148
rect 8576 35096 8628 35148
rect 9036 35096 9088 35148
rect 10416 35164 10468 35216
rect 10784 35096 10836 35148
rect 4712 35028 4764 35080
rect 2688 34960 2740 35012
rect 1860 34892 1912 34944
rect 3424 34960 3476 35012
rect 3700 34892 3752 34944
rect 8576 34960 8628 35012
rect 9128 34960 9180 35012
rect 8852 34892 8904 34944
rect 9404 35003 9456 35012
rect 9404 34969 9413 35003
rect 9413 34969 9447 35003
rect 9447 34969 9456 35003
rect 9404 34960 9456 34969
rect 9864 34960 9916 35012
rect 15016 34960 15068 35012
rect 10784 34892 10836 34944
rect 15108 34892 15160 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2044 34688 2096 34740
rect 2412 34688 2464 34740
rect 3884 34688 3936 34740
rect 5540 34688 5592 34740
rect 5172 34620 5224 34672
rect 9036 34688 9088 34740
rect 10968 34688 11020 34740
rect 11152 34688 11204 34740
rect 11336 34688 11388 34740
rect 11980 34663 12032 34672
rect 11980 34629 11989 34663
rect 11989 34629 12023 34663
rect 12023 34629 12032 34663
rect 11980 34620 12032 34629
rect 13452 34688 13504 34740
rect 1676 34348 1728 34400
rect 3516 34484 3568 34536
rect 4804 34484 4856 34536
rect 5908 34484 5960 34536
rect 6828 34484 6880 34536
rect 8392 34416 8444 34468
rect 9956 34484 10008 34536
rect 12348 34527 12400 34536
rect 12348 34493 12357 34527
rect 12357 34493 12391 34527
rect 12391 34493 12400 34527
rect 12348 34484 12400 34493
rect 13820 34484 13872 34536
rect 37832 34484 37884 34536
rect 38292 34527 38344 34536
rect 38292 34493 38301 34527
rect 38301 34493 38335 34527
rect 38335 34493 38344 34527
rect 38292 34484 38344 34493
rect 12440 34416 12492 34468
rect 3884 34348 3936 34400
rect 4620 34348 4672 34400
rect 6920 34348 6972 34400
rect 8852 34391 8904 34400
rect 8852 34357 8861 34391
rect 8861 34357 8895 34391
rect 8895 34357 8904 34391
rect 8852 34348 8904 34357
rect 9956 34348 10008 34400
rect 10232 34348 10284 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 8300 34144 8352 34196
rect 11060 34144 11112 34196
rect 1676 34051 1728 34060
rect 1676 34017 1685 34051
rect 1685 34017 1719 34051
rect 1719 34017 1728 34051
rect 1676 34008 1728 34017
rect 3792 34008 3844 34060
rect 3884 34008 3936 34060
rect 5172 34051 5224 34060
rect 5172 34017 5181 34051
rect 5181 34017 5215 34051
rect 5215 34017 5224 34051
rect 14004 34076 14056 34128
rect 38292 34119 38344 34128
rect 38292 34085 38301 34119
rect 38301 34085 38335 34119
rect 38335 34085 38344 34119
rect 38292 34076 38344 34085
rect 5172 34008 5224 34017
rect 8392 34008 8444 34060
rect 14740 34008 14792 34060
rect 4436 33983 4488 33992
rect 4436 33949 4445 33983
rect 4445 33949 4479 33983
rect 4479 33949 4488 33983
rect 4436 33940 4488 33949
rect 6644 33940 6696 33992
rect 13544 33983 13596 33992
rect 2964 33872 3016 33924
rect 5080 33872 5132 33924
rect 5724 33872 5776 33924
rect 8208 33872 8260 33924
rect 9312 33872 9364 33924
rect 9864 33872 9916 33924
rect 11796 33915 11848 33924
rect 11796 33881 11805 33915
rect 11805 33881 11839 33915
rect 11839 33881 11848 33915
rect 11796 33872 11848 33881
rect 12348 33915 12400 33924
rect 12348 33881 12357 33915
rect 12357 33881 12391 33915
rect 12391 33881 12400 33915
rect 12348 33872 12400 33881
rect 7472 33804 7524 33856
rect 7564 33804 7616 33856
rect 10416 33804 10468 33856
rect 11152 33804 11204 33856
rect 13544 33949 13553 33983
rect 13553 33949 13587 33983
rect 13587 33949 13596 33983
rect 13544 33940 13596 33949
rect 14924 33983 14976 33992
rect 14924 33949 14933 33983
rect 14933 33949 14967 33983
rect 14967 33949 14976 33983
rect 14924 33940 14976 33949
rect 14832 33872 14884 33924
rect 14188 33804 14240 33856
rect 14280 33847 14332 33856
rect 14280 33813 14289 33847
rect 14289 33813 14323 33847
rect 14323 33813 14332 33847
rect 14280 33804 14332 33813
rect 14556 33804 14608 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 3792 33600 3844 33652
rect 6552 33600 6604 33652
rect 7748 33600 7800 33652
rect 9128 33600 9180 33652
rect 9312 33600 9364 33652
rect 2044 33532 2096 33584
rect 3608 33532 3660 33584
rect 8668 33532 8720 33584
rect 9036 33532 9088 33584
rect 2596 33464 2648 33516
rect 3976 33507 4028 33516
rect 3976 33473 3985 33507
rect 3985 33473 4019 33507
rect 4019 33473 4028 33507
rect 3976 33464 4028 33473
rect 4436 33464 4488 33516
rect 6828 33464 6880 33516
rect 7012 33464 7064 33516
rect 8392 33507 8444 33516
rect 8392 33473 8401 33507
rect 8401 33473 8435 33507
rect 8435 33473 8444 33507
rect 8852 33507 8904 33516
rect 8392 33464 8444 33473
rect 8852 33473 8861 33507
rect 8861 33473 8895 33507
rect 8895 33473 8904 33507
rect 8852 33464 8904 33473
rect 10416 33464 10468 33516
rect 11980 33600 12032 33652
rect 12348 33600 12400 33652
rect 14188 33575 14240 33584
rect 14188 33541 14197 33575
rect 14197 33541 14231 33575
rect 14231 33541 14240 33575
rect 14188 33532 14240 33541
rect 2320 33396 2372 33448
rect 3148 33396 3200 33448
rect 4712 33439 4764 33448
rect 4712 33405 4721 33439
rect 4721 33405 4755 33439
rect 4755 33405 4764 33439
rect 4712 33396 4764 33405
rect 5632 33439 5684 33448
rect 5632 33405 5641 33439
rect 5641 33405 5675 33439
rect 5675 33405 5684 33439
rect 5632 33396 5684 33405
rect 7472 33396 7524 33448
rect 9220 33396 9272 33448
rect 9588 33396 9640 33448
rect 11980 33464 12032 33516
rect 13912 33464 13964 33516
rect 14280 33396 14332 33448
rect 2044 33260 2096 33312
rect 5540 33260 5592 33312
rect 6920 33260 6972 33312
rect 7656 33260 7708 33312
rect 7748 33260 7800 33312
rect 11980 33328 12032 33380
rect 13820 33328 13872 33380
rect 14924 33328 14976 33380
rect 10232 33260 10284 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4068 33099 4120 33108
rect 4068 33065 4077 33099
rect 4077 33065 4111 33099
rect 4111 33065 4120 33099
rect 4068 33056 4120 33065
rect 8576 33056 8628 33108
rect 8852 33056 8904 33108
rect 9588 33056 9640 33108
rect 10876 33099 10928 33108
rect 10876 33065 10885 33099
rect 10885 33065 10919 33099
rect 10919 33065 10928 33099
rect 10876 33056 10928 33065
rect 11796 33056 11848 33108
rect 6920 32988 6972 33040
rect 7748 32988 7800 33040
rect 3884 32920 3936 32972
rect 5172 32920 5224 32972
rect 4620 32852 4672 32904
rect 10140 32920 10192 32972
rect 10324 32920 10376 32972
rect 1860 32716 1912 32768
rect 4344 32784 4396 32836
rect 6828 32895 6880 32904
rect 6828 32861 6837 32895
rect 6837 32861 6871 32895
rect 6871 32861 6880 32895
rect 6828 32852 6880 32861
rect 11060 32852 11112 32904
rect 5172 32784 5224 32836
rect 8760 32784 8812 32836
rect 3240 32716 3292 32768
rect 3608 32716 3660 32768
rect 12532 32716 12584 32768
rect 23112 32716 23164 32768
rect 38200 32827 38252 32836
rect 38200 32793 38209 32827
rect 38209 32793 38243 32827
rect 38243 32793 38252 32827
rect 38200 32784 38252 32793
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 3884 32512 3936 32564
rect 2872 32444 2924 32496
rect 4620 32444 4672 32496
rect 4804 32444 4856 32496
rect 2780 32376 2832 32428
rect 5908 32512 5960 32564
rect 2412 32308 2464 32360
rect 4344 32308 4396 32360
rect 6736 32444 6788 32496
rect 7196 32444 7248 32496
rect 14464 32444 14516 32496
rect 15016 32487 15068 32496
rect 15016 32453 15025 32487
rect 15025 32453 15059 32487
rect 15059 32453 15068 32487
rect 15016 32444 15068 32453
rect 16028 32444 16080 32496
rect 5264 32376 5316 32428
rect 5632 32419 5684 32428
rect 5632 32385 5641 32419
rect 5641 32385 5675 32419
rect 5675 32385 5684 32419
rect 5632 32376 5684 32385
rect 8852 32419 8904 32428
rect 8852 32385 8861 32419
rect 8861 32385 8895 32419
rect 8895 32385 8904 32419
rect 8852 32376 8904 32385
rect 13176 32419 13228 32428
rect 8576 32351 8628 32360
rect 8576 32317 8585 32351
rect 8585 32317 8619 32351
rect 8619 32317 8628 32351
rect 8576 32308 8628 32317
rect 5632 32172 5684 32224
rect 6736 32172 6788 32224
rect 13176 32385 13185 32419
rect 13185 32385 13219 32419
rect 13219 32385 13228 32419
rect 13176 32376 13228 32385
rect 15568 32308 15620 32360
rect 15936 32240 15988 32292
rect 16212 32172 16264 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 8208 31968 8260 32020
rect 8852 31968 8904 32020
rect 9312 31968 9364 32020
rect 6276 31900 6328 31952
rect 6644 31900 6696 31952
rect 1952 31875 2004 31884
rect 1952 31841 1961 31875
rect 1961 31841 1995 31875
rect 1995 31841 2004 31875
rect 1952 31832 2004 31841
rect 3424 31875 3476 31884
rect 3424 31841 3433 31875
rect 3433 31841 3467 31875
rect 3467 31841 3476 31875
rect 3424 31832 3476 31841
rect 4160 31832 4212 31884
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 3608 31696 3660 31748
rect 4160 31628 4212 31680
rect 6276 31764 6328 31816
rect 6552 31832 6604 31884
rect 8576 31875 8628 31884
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 8576 31841 8585 31875
rect 8585 31841 8619 31875
rect 8619 31841 8628 31875
rect 8576 31832 8628 31841
rect 12256 31832 12308 31884
rect 12900 31764 12952 31816
rect 15752 31764 15804 31816
rect 23112 31764 23164 31816
rect 5172 31628 5224 31680
rect 6368 31696 6420 31748
rect 5908 31628 5960 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1676 31424 1728 31476
rect 3884 31424 3936 31476
rect 3792 31356 3844 31408
rect 4160 31424 4212 31476
rect 6736 31424 6788 31476
rect 7288 31424 7340 31476
rect 8024 31399 8076 31408
rect 8024 31365 8033 31399
rect 8033 31365 8067 31399
rect 8067 31365 8076 31399
rect 8024 31356 8076 31365
rect 11152 31356 11204 31408
rect 5632 31288 5684 31340
rect 6000 31288 6052 31340
rect 6736 31288 6788 31340
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 1492 31220 1544 31272
rect 3700 31084 3752 31136
rect 3884 31084 3936 31136
rect 4620 31220 4672 31272
rect 5264 31220 5316 31272
rect 6920 31152 6972 31204
rect 9312 31220 9364 31272
rect 8944 31152 8996 31204
rect 15108 31356 15160 31408
rect 20444 31331 20496 31340
rect 20444 31297 20453 31331
rect 20453 31297 20487 31331
rect 20487 31297 20496 31331
rect 20444 31288 20496 31297
rect 15384 31263 15436 31272
rect 15384 31229 15393 31263
rect 15393 31229 15427 31263
rect 15427 31229 15436 31263
rect 15384 31220 15436 31229
rect 16028 31220 16080 31272
rect 18052 31220 18104 31272
rect 17960 31152 18012 31204
rect 5724 31127 5776 31136
rect 5724 31093 5733 31127
rect 5733 31093 5767 31127
rect 5767 31093 5776 31127
rect 5724 31084 5776 31093
rect 6184 31084 6236 31136
rect 8760 31084 8812 31136
rect 9680 31084 9732 31136
rect 14648 31127 14700 31136
rect 14648 31093 14657 31127
rect 14657 31093 14691 31127
rect 14691 31093 14700 31127
rect 14648 31084 14700 31093
rect 38016 31084 38068 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2044 30880 2096 30932
rect 2964 30880 3016 30932
rect 3148 30923 3200 30932
rect 3148 30889 3157 30923
rect 3157 30889 3191 30923
rect 3191 30889 3200 30923
rect 3148 30880 3200 30889
rect 3240 30719 3292 30728
rect 3240 30685 3249 30719
rect 3249 30685 3283 30719
rect 3283 30685 3292 30719
rect 3240 30676 3292 30685
rect 3424 30676 3476 30728
rect 4528 30812 4580 30864
rect 5632 30880 5684 30932
rect 5724 30880 5776 30932
rect 13176 30880 13228 30932
rect 16028 30880 16080 30932
rect 16304 30923 16356 30932
rect 16304 30889 16313 30923
rect 16313 30889 16347 30923
rect 16347 30889 16356 30923
rect 16304 30880 16356 30889
rect 16856 30923 16908 30932
rect 16856 30889 16865 30923
rect 16865 30889 16899 30923
rect 16899 30889 16908 30923
rect 16856 30880 16908 30889
rect 37556 30923 37608 30932
rect 37556 30889 37565 30923
rect 37565 30889 37599 30923
rect 37599 30889 37608 30923
rect 37556 30880 37608 30889
rect 5172 30812 5224 30864
rect 5264 30812 5316 30864
rect 8024 30812 8076 30864
rect 6644 30744 6696 30796
rect 6828 30744 6880 30796
rect 6920 30744 6972 30796
rect 5172 30676 5224 30728
rect 5724 30676 5776 30728
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8116 30676 8168 30685
rect 20444 30812 20496 30864
rect 11980 30744 12032 30796
rect 12440 30744 12492 30796
rect 14556 30787 14608 30796
rect 14556 30753 14565 30787
rect 14565 30753 14599 30787
rect 14599 30753 14608 30787
rect 14556 30744 14608 30753
rect 16488 30676 16540 30728
rect 38016 30719 38068 30728
rect 3240 30540 3292 30592
rect 5080 30540 5132 30592
rect 6920 30540 6972 30592
rect 12348 30651 12400 30660
rect 12348 30617 12357 30651
rect 12357 30617 12391 30651
rect 12391 30617 12400 30651
rect 12348 30608 12400 30617
rect 14648 30651 14700 30660
rect 14648 30617 14657 30651
rect 14657 30617 14691 30651
rect 14691 30617 14700 30651
rect 14648 30608 14700 30617
rect 15292 30608 15344 30660
rect 38016 30685 38025 30719
rect 38025 30685 38059 30719
rect 38059 30685 38068 30719
rect 38016 30676 38068 30685
rect 38108 30608 38160 30660
rect 8300 30540 8352 30592
rect 9588 30540 9640 30592
rect 15476 30540 15528 30592
rect 38200 30583 38252 30592
rect 38200 30549 38209 30583
rect 38209 30549 38243 30583
rect 38243 30549 38252 30583
rect 38200 30540 38252 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1952 30336 2004 30388
rect 8116 30336 8168 30388
rect 12348 30379 12400 30388
rect 12348 30345 12357 30379
rect 12357 30345 12391 30379
rect 12391 30345 12400 30379
rect 12348 30336 12400 30345
rect 3148 30268 3200 30320
rect 3792 30268 3844 30320
rect 5448 30311 5500 30320
rect 5448 30277 5457 30311
rect 5457 30277 5491 30311
rect 5491 30277 5500 30311
rect 5448 30268 5500 30277
rect 5816 30268 5868 30320
rect 6736 30268 6788 30320
rect 3240 30200 3292 30252
rect 4528 30200 4580 30252
rect 4712 30243 4764 30252
rect 4712 30209 4721 30243
rect 4721 30209 4755 30243
rect 4755 30209 4764 30243
rect 4712 30200 4764 30209
rect 5724 30200 5776 30252
rect 2872 30132 2924 30184
rect 8668 30200 8720 30252
rect 6828 30132 6880 30184
rect 13084 30268 13136 30320
rect 13544 30268 13596 30320
rect 15752 30268 15804 30320
rect 16120 30311 16172 30320
rect 16120 30277 16129 30311
rect 16129 30277 16163 30311
rect 16163 30277 16172 30311
rect 16120 30268 16172 30277
rect 9220 30200 9272 30252
rect 12256 30200 12308 30252
rect 14372 30132 14424 30184
rect 14740 30132 14792 30184
rect 17500 30132 17552 30184
rect 9496 30064 9548 30116
rect 6460 29996 6512 30048
rect 6736 29996 6788 30048
rect 8208 29996 8260 30048
rect 13452 29996 13504 30048
rect 16672 29996 16724 30048
rect 17960 30039 18012 30048
rect 17960 30005 17969 30039
rect 17969 30005 18003 30039
rect 18003 30005 18012 30039
rect 17960 29996 18012 30005
rect 18420 30039 18472 30048
rect 18420 30005 18429 30039
rect 18429 30005 18463 30039
rect 18463 30005 18472 30039
rect 18420 29996 18472 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2688 29792 2740 29844
rect 4896 29835 4948 29844
rect 4896 29801 4905 29835
rect 4905 29801 4939 29835
rect 4939 29801 4948 29835
rect 4896 29792 4948 29801
rect 6092 29724 6144 29776
rect 3332 29656 3384 29708
rect 3608 29656 3660 29708
rect 2044 29588 2096 29640
rect 3240 29588 3292 29640
rect 4712 29588 4764 29640
rect 7288 29792 7340 29844
rect 7748 29792 7800 29844
rect 12532 29835 12584 29844
rect 12532 29801 12541 29835
rect 12541 29801 12575 29835
rect 12575 29801 12584 29835
rect 12532 29792 12584 29801
rect 16120 29792 16172 29844
rect 15292 29699 15344 29708
rect 15292 29665 15301 29699
rect 15301 29665 15335 29699
rect 15335 29665 15344 29699
rect 15292 29656 15344 29665
rect 16120 29656 16172 29708
rect 6736 29588 6788 29640
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 2412 29452 2464 29504
rect 10324 29520 10376 29572
rect 12256 29588 12308 29640
rect 13820 29588 13872 29640
rect 14464 29588 14516 29640
rect 16856 29588 16908 29640
rect 18420 29588 18472 29640
rect 37832 29588 37884 29640
rect 13360 29452 13412 29504
rect 14280 29452 14332 29504
rect 14832 29452 14884 29504
rect 17868 29520 17920 29572
rect 17408 29452 17460 29504
rect 18604 29452 18656 29504
rect 30012 29495 30064 29504
rect 30012 29461 30021 29495
rect 30021 29461 30055 29495
rect 30055 29461 30064 29495
rect 30012 29452 30064 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2320 29248 2372 29300
rect 2504 29248 2556 29300
rect 2044 28976 2096 29028
rect 2964 29180 3016 29232
rect 4804 29180 4856 29232
rect 6552 29248 6604 29300
rect 7288 29291 7340 29300
rect 7288 29257 7297 29291
rect 7297 29257 7331 29291
rect 7331 29257 7340 29291
rect 7288 29248 7340 29257
rect 13544 29291 13596 29300
rect 13544 29257 13553 29291
rect 13553 29257 13587 29291
rect 13587 29257 13596 29291
rect 13544 29248 13596 29257
rect 20352 29291 20404 29300
rect 20352 29257 20361 29291
rect 20361 29257 20395 29291
rect 20395 29257 20404 29291
rect 20352 29248 20404 29257
rect 6828 29180 6880 29232
rect 3240 29112 3292 29164
rect 3424 29155 3476 29164
rect 3424 29121 3433 29155
rect 3433 29121 3467 29155
rect 3467 29121 3476 29155
rect 3424 29112 3476 29121
rect 4712 29155 4764 29164
rect 4712 29121 4721 29155
rect 4721 29121 4755 29155
rect 4755 29121 4764 29155
rect 4712 29112 4764 29121
rect 8300 29223 8352 29232
rect 8300 29189 8309 29223
rect 8309 29189 8343 29223
rect 8343 29189 8352 29223
rect 8300 29180 8352 29189
rect 12072 29223 12124 29232
rect 12072 29189 12081 29223
rect 12081 29189 12115 29223
rect 12115 29189 12124 29223
rect 12072 29180 12124 29189
rect 14280 29223 14332 29232
rect 14280 29189 14289 29223
rect 14289 29189 14323 29223
rect 14323 29189 14332 29223
rect 14280 29180 14332 29189
rect 14372 29180 14424 29232
rect 15568 29180 15620 29232
rect 16304 29180 16356 29232
rect 17408 29223 17460 29232
rect 17408 29189 17417 29223
rect 17417 29189 17451 29223
rect 17451 29189 17460 29223
rect 17408 29180 17460 29189
rect 18052 29223 18104 29232
rect 18052 29189 18061 29223
rect 18061 29189 18095 29223
rect 18095 29189 18104 29223
rect 18052 29180 18104 29189
rect 18604 29223 18656 29232
rect 18604 29189 18613 29223
rect 18613 29189 18647 29223
rect 18647 29189 18656 29223
rect 18604 29180 18656 29189
rect 10324 29155 10376 29164
rect 10324 29121 10333 29155
rect 10333 29121 10367 29155
rect 10367 29121 10376 29155
rect 10324 29112 10376 29121
rect 12808 29112 12860 29164
rect 20076 29112 20128 29164
rect 38200 29155 38252 29164
rect 38200 29121 38209 29155
rect 38209 29121 38243 29155
rect 38243 29121 38252 29155
rect 38200 29112 38252 29121
rect 7012 29044 7064 29096
rect 8208 29087 8260 29096
rect 8208 29053 8217 29087
rect 8217 29053 8251 29087
rect 8251 29053 8260 29087
rect 8208 29044 8260 29053
rect 9128 29044 9180 29096
rect 11980 29087 12032 29096
rect 11980 29053 11989 29087
rect 11989 29053 12023 29087
rect 12023 29053 12032 29087
rect 11980 29044 12032 29053
rect 12624 29087 12676 29096
rect 12624 29053 12633 29087
rect 12633 29053 12667 29087
rect 12667 29053 12676 29087
rect 12624 29044 12676 29053
rect 14188 29087 14240 29096
rect 14188 29053 14197 29087
rect 14197 29053 14231 29087
rect 14231 29053 14240 29087
rect 14188 29044 14240 29053
rect 15476 29044 15528 29096
rect 16120 29044 16172 29096
rect 17500 29087 17552 29096
rect 17500 29053 17509 29087
rect 17509 29053 17543 29087
rect 17543 29053 17552 29087
rect 17500 29044 17552 29053
rect 3424 28976 3476 29028
rect 2964 28908 3016 28960
rect 9772 28976 9824 29028
rect 10876 28976 10928 29028
rect 14740 29019 14792 29028
rect 14740 28985 14749 29019
rect 14749 28985 14783 29019
rect 14783 28985 14792 29019
rect 14740 28976 14792 28985
rect 15200 28976 15252 29028
rect 30012 28976 30064 29028
rect 37280 28976 37332 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2780 28704 2832 28756
rect 5356 28704 5408 28756
rect 6276 28704 6328 28756
rect 7196 28747 7248 28756
rect 7196 28713 7205 28747
rect 7205 28713 7239 28747
rect 7239 28713 7248 28747
rect 7196 28704 7248 28713
rect 7288 28704 7340 28756
rect 11336 28747 11388 28756
rect 11336 28713 11345 28747
rect 11345 28713 11379 28747
rect 11379 28713 11388 28747
rect 11336 28704 11388 28713
rect 12072 28704 12124 28756
rect 14372 28704 14424 28756
rect 14832 28704 14884 28756
rect 18512 28704 18564 28756
rect 2228 28679 2280 28688
rect 2228 28645 2237 28679
rect 2237 28645 2271 28679
rect 2271 28645 2280 28679
rect 2228 28636 2280 28645
rect 2596 28636 2648 28688
rect 9864 28636 9916 28688
rect 12532 28636 12584 28688
rect 8484 28568 8536 28620
rect 12624 28568 12676 28620
rect 2780 28543 2832 28552
rect 2780 28509 2789 28543
rect 2789 28509 2823 28543
rect 2823 28509 2832 28543
rect 2780 28500 2832 28509
rect 3240 28500 3292 28552
rect 3424 28500 3476 28552
rect 4712 28543 4764 28552
rect 4712 28509 4721 28543
rect 4721 28509 4755 28543
rect 4755 28509 4764 28543
rect 4712 28500 4764 28509
rect 7288 28500 7340 28552
rect 9956 28500 10008 28552
rect 11888 28543 11940 28552
rect 11888 28509 11897 28543
rect 11897 28509 11931 28543
rect 11931 28509 11940 28543
rect 11888 28500 11940 28509
rect 12808 28500 12860 28552
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 17684 28636 17736 28688
rect 14740 28568 14792 28620
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 16856 28568 16908 28620
rect 17868 28568 17920 28620
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 17960 28500 18012 28552
rect 9128 28475 9180 28484
rect 9128 28441 9137 28475
rect 9137 28441 9171 28475
rect 9171 28441 9180 28475
rect 9128 28432 9180 28441
rect 9680 28475 9732 28484
rect 9680 28441 9689 28475
rect 9689 28441 9723 28475
rect 9723 28441 9732 28475
rect 9680 28432 9732 28441
rect 13268 28432 13320 28484
rect 14464 28475 14516 28484
rect 14464 28441 14473 28475
rect 14473 28441 14507 28475
rect 14507 28441 14516 28475
rect 14464 28432 14516 28441
rect 18420 28500 18472 28552
rect 20076 28543 20128 28552
rect 20076 28509 20085 28543
rect 20085 28509 20119 28543
rect 20119 28509 20128 28543
rect 20076 28500 20128 28509
rect 1860 28364 1912 28416
rect 7380 28364 7432 28416
rect 13176 28364 13228 28416
rect 15752 28364 15804 28416
rect 16212 28364 16264 28416
rect 18512 28432 18564 28484
rect 37832 28543 37884 28552
rect 37832 28509 37841 28543
rect 37841 28509 37875 28543
rect 37875 28509 37884 28543
rect 37832 28500 37884 28509
rect 36268 28432 36320 28484
rect 16764 28364 16816 28416
rect 18788 28407 18840 28416
rect 18788 28373 18797 28407
rect 18797 28373 18831 28407
rect 18831 28373 18840 28407
rect 18788 28364 18840 28373
rect 20444 28364 20496 28416
rect 38016 28407 38068 28416
rect 38016 28373 38025 28407
rect 38025 28373 38059 28407
rect 38059 28373 38068 28407
rect 38016 28364 38068 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3516 28203 3568 28212
rect 3516 28169 3525 28203
rect 3525 28169 3559 28203
rect 3559 28169 3568 28203
rect 3516 28160 3568 28169
rect 4620 28160 4672 28212
rect 7288 28160 7340 28212
rect 14464 28160 14516 28212
rect 7104 28092 7156 28144
rect 7564 28092 7616 28144
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 2780 28067 2832 28076
rect 2780 28033 2789 28067
rect 2789 28033 2823 28067
rect 2823 28033 2832 28067
rect 2780 28024 2832 28033
rect 3424 28024 3476 28076
rect 10232 28024 10284 28076
rect 11888 28092 11940 28144
rect 13636 28092 13688 28144
rect 13820 28092 13872 28144
rect 15752 28135 15804 28144
rect 15752 28101 15761 28135
rect 15761 28101 15795 28135
rect 15795 28101 15804 28135
rect 15752 28092 15804 28101
rect 15936 28092 15988 28144
rect 7380 27956 7432 28008
rect 12900 28024 12952 28076
rect 13360 28024 13412 28076
rect 13728 28067 13780 28076
rect 13728 28033 13737 28067
rect 13737 28033 13771 28067
rect 13771 28033 13780 28067
rect 13728 28024 13780 28033
rect 16304 28067 16356 28076
rect 16304 28033 16313 28067
rect 16313 28033 16347 28067
rect 16347 28033 16356 28067
rect 23664 28067 23716 28076
rect 16304 28024 16356 28033
rect 23664 28033 23673 28067
rect 23673 28033 23707 28067
rect 23707 28033 23716 28067
rect 23664 28024 23716 28033
rect 14280 27956 14332 28008
rect 15476 27956 15528 28008
rect 17868 27999 17920 28008
rect 12440 27888 12492 27940
rect 14556 27888 14608 27940
rect 15384 27888 15436 27940
rect 10048 27863 10100 27872
rect 10048 27829 10057 27863
rect 10057 27829 10091 27863
rect 10091 27829 10100 27863
rect 10048 27820 10100 27829
rect 10968 27820 11020 27872
rect 14188 27820 14240 27872
rect 17868 27965 17877 27999
rect 17877 27965 17911 27999
rect 17911 27965 17920 27999
rect 17868 27956 17920 27965
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 18696 27999 18748 28008
rect 18696 27965 18705 27999
rect 18705 27965 18739 27999
rect 18739 27965 18748 27999
rect 18696 27956 18748 27965
rect 19340 27999 19392 28008
rect 19340 27965 19349 27999
rect 19349 27965 19383 27999
rect 19383 27965 19392 27999
rect 19340 27956 19392 27965
rect 20352 27888 20404 27940
rect 17316 27820 17368 27872
rect 19984 27820 20036 27872
rect 34796 27888 34848 27940
rect 38292 27820 38344 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 10048 27616 10100 27668
rect 14648 27616 14700 27668
rect 16028 27616 16080 27668
rect 17316 27616 17368 27668
rect 1584 27591 1636 27600
rect 1584 27557 1593 27591
rect 1593 27557 1627 27591
rect 1627 27557 1636 27591
rect 1584 27548 1636 27557
rect 11244 27548 11296 27600
rect 14372 27548 14424 27600
rect 14740 27548 14792 27600
rect 17776 27548 17828 27600
rect 9128 27387 9180 27396
rect 9128 27353 9137 27387
rect 9137 27353 9171 27387
rect 9171 27353 9180 27387
rect 9128 27344 9180 27353
rect 9588 27344 9640 27396
rect 10876 27387 10928 27396
rect 10876 27353 10885 27387
rect 10885 27353 10919 27387
rect 10919 27353 10928 27387
rect 10876 27344 10928 27353
rect 10968 27387 11020 27396
rect 10968 27353 10977 27387
rect 10977 27353 11011 27387
rect 11011 27353 11020 27387
rect 10968 27344 11020 27353
rect 11336 27344 11388 27396
rect 12532 27480 12584 27532
rect 13360 27523 13412 27532
rect 13360 27489 13369 27523
rect 13369 27489 13403 27523
rect 13403 27489 13412 27523
rect 13360 27480 13412 27489
rect 15844 27480 15896 27532
rect 16488 27480 16540 27532
rect 16856 27523 16908 27532
rect 16856 27489 16865 27523
rect 16865 27489 16899 27523
rect 16899 27489 16908 27523
rect 16856 27480 16908 27489
rect 17132 27523 17184 27532
rect 17132 27489 17141 27523
rect 17141 27489 17175 27523
rect 17175 27489 17184 27523
rect 17132 27480 17184 27489
rect 17960 27523 18012 27532
rect 17960 27489 17969 27523
rect 17969 27489 18003 27523
rect 18003 27489 18012 27523
rect 17960 27480 18012 27489
rect 19340 27480 19392 27532
rect 14372 27412 14424 27464
rect 18512 27412 18564 27464
rect 12808 27344 12860 27396
rect 13084 27387 13136 27396
rect 13084 27353 13093 27387
rect 13093 27353 13127 27387
rect 13127 27353 13136 27387
rect 13084 27344 13136 27353
rect 13176 27387 13228 27396
rect 13176 27353 13185 27387
rect 13185 27353 13219 27387
rect 13219 27353 13228 27387
rect 13176 27344 13228 27353
rect 14280 27344 14332 27396
rect 15660 27344 15712 27396
rect 12716 27276 12768 27328
rect 15752 27276 15804 27328
rect 15936 27344 15988 27396
rect 16856 27344 16908 27396
rect 16764 27276 16816 27328
rect 18788 27344 18840 27396
rect 20076 27387 20128 27396
rect 20076 27353 20085 27387
rect 20085 27353 20119 27387
rect 20119 27353 20128 27387
rect 20076 27344 20128 27353
rect 18328 27276 18380 27328
rect 18420 27276 18472 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8392 27072 8444 27124
rect 12348 27072 12400 27124
rect 13820 27072 13872 27124
rect 14188 27072 14240 27124
rect 13360 27004 13412 27056
rect 14556 27047 14608 27056
rect 14556 27013 14565 27047
rect 14565 27013 14599 27047
rect 14599 27013 14608 27047
rect 14556 27004 14608 27013
rect 17224 27072 17276 27124
rect 17408 27072 17460 27124
rect 37280 27072 37332 27124
rect 15660 27004 15712 27056
rect 16764 27004 16816 27056
rect 13544 26979 13596 26988
rect 10048 26911 10100 26920
rect 10048 26877 10057 26911
rect 10057 26877 10091 26911
rect 10091 26877 10100 26911
rect 10048 26868 10100 26877
rect 10600 26911 10652 26920
rect 10600 26877 10609 26911
rect 10609 26877 10643 26911
rect 10643 26877 10652 26911
rect 10600 26868 10652 26877
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 12256 26868 12308 26920
rect 11244 26800 11296 26852
rect 13084 26800 13136 26852
rect 12440 26732 12492 26784
rect 15200 26911 15252 26920
rect 15200 26877 15209 26911
rect 15209 26877 15243 26911
rect 15243 26877 15252 26911
rect 15200 26868 15252 26877
rect 18236 27004 18288 27056
rect 18420 27047 18472 27056
rect 18420 27013 18429 27047
rect 18429 27013 18463 27047
rect 18463 27013 18472 27047
rect 18420 27004 18472 27013
rect 18696 27004 18748 27056
rect 17316 26979 17368 26988
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 19616 27004 19668 27056
rect 20352 27047 20404 27056
rect 20352 27013 20361 27047
rect 20361 27013 20395 27047
rect 20395 27013 20404 27047
rect 20352 27004 20404 27013
rect 17316 26936 17368 26945
rect 38016 26979 38068 26988
rect 18144 26911 18196 26920
rect 18144 26877 18153 26911
rect 18153 26877 18187 26911
rect 18187 26877 18196 26911
rect 18144 26868 18196 26877
rect 18236 26868 18288 26920
rect 20168 26868 20220 26920
rect 17408 26800 17460 26852
rect 17500 26800 17552 26852
rect 38016 26945 38025 26979
rect 38025 26945 38059 26979
rect 38059 26945 38068 26979
rect 38016 26936 38068 26945
rect 17040 26732 17092 26784
rect 18788 26732 18840 26784
rect 20352 26732 20404 26784
rect 38200 26775 38252 26784
rect 38200 26741 38209 26775
rect 38209 26741 38243 26775
rect 38243 26741 38252 26775
rect 38200 26732 38252 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11980 26528 12032 26580
rect 16948 26528 17000 26580
rect 17684 26528 17736 26580
rect 20076 26528 20128 26580
rect 9404 26392 9456 26444
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 14740 26460 14792 26512
rect 12624 26392 12676 26444
rect 15384 26435 15436 26444
rect 15384 26401 15393 26435
rect 15393 26401 15427 26435
rect 15427 26401 15436 26435
rect 15384 26392 15436 26401
rect 15660 26392 15712 26444
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 16488 26392 16540 26444
rect 18788 26435 18840 26444
rect 18788 26401 18797 26435
rect 18797 26401 18831 26435
rect 18831 26401 18840 26435
rect 18788 26392 18840 26401
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 2136 26256 2188 26308
rect 11244 26324 11296 26376
rect 11520 26299 11572 26308
rect 11520 26265 11529 26299
rect 11529 26265 11563 26299
rect 11563 26265 11572 26299
rect 12624 26299 12676 26308
rect 11520 26256 11572 26265
rect 12624 26265 12633 26299
rect 12633 26265 12667 26299
rect 12667 26265 12676 26299
rect 12624 26256 12676 26265
rect 12716 26299 12768 26308
rect 12716 26265 12725 26299
rect 12725 26265 12759 26299
rect 12759 26265 12768 26299
rect 12716 26256 12768 26265
rect 13452 26256 13504 26308
rect 1676 26231 1728 26240
rect 1676 26197 1685 26231
rect 1685 26197 1719 26231
rect 1719 26197 1728 26231
rect 1676 26188 1728 26197
rect 9404 26231 9456 26240
rect 9404 26197 9413 26231
rect 9413 26197 9447 26231
rect 9447 26197 9456 26231
rect 9404 26188 9456 26197
rect 15200 26256 15252 26308
rect 15660 26256 15712 26308
rect 16488 26256 16540 26308
rect 17500 26299 17552 26308
rect 17500 26265 17509 26299
rect 17509 26265 17543 26299
rect 17543 26265 17552 26299
rect 17500 26256 17552 26265
rect 17776 26256 17828 26308
rect 20352 26367 20404 26376
rect 20352 26333 20361 26367
rect 20361 26333 20395 26367
rect 20395 26333 20404 26367
rect 20352 26324 20404 26333
rect 19616 26299 19668 26308
rect 19616 26265 19625 26299
rect 19625 26265 19659 26299
rect 19659 26265 19668 26299
rect 19616 26256 19668 26265
rect 17684 26188 17736 26240
rect 38108 26324 38160 26376
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9404 25848 9456 25900
rect 11336 25916 11388 25968
rect 12624 25959 12676 25968
rect 12624 25925 12633 25959
rect 12633 25925 12667 25959
rect 12667 25925 12676 25959
rect 12624 25916 12676 25925
rect 16304 25984 16356 26036
rect 18328 25984 18380 26036
rect 20904 26027 20956 26036
rect 20904 25993 20913 26027
rect 20913 25993 20947 26027
rect 20947 25993 20956 26027
rect 20904 25984 20956 25993
rect 15752 25916 15804 25968
rect 16580 25916 16632 25968
rect 17960 25916 18012 25968
rect 19524 25916 19576 25968
rect 12900 25848 12952 25900
rect 14464 25848 14516 25900
rect 16856 25848 16908 25900
rect 20076 25848 20128 25900
rect 21456 25848 21508 25900
rect 15936 25823 15988 25832
rect 9772 25687 9824 25696
rect 9772 25653 9781 25687
rect 9781 25653 9815 25687
rect 9815 25653 9824 25687
rect 9772 25644 9824 25653
rect 11612 25712 11664 25764
rect 15936 25789 15945 25823
rect 15945 25789 15979 25823
rect 15979 25789 15988 25823
rect 15936 25780 15988 25789
rect 16764 25780 16816 25832
rect 17684 25823 17736 25832
rect 17684 25789 17693 25823
rect 17693 25789 17727 25823
rect 17727 25789 17736 25823
rect 17684 25780 17736 25789
rect 21640 25780 21692 25832
rect 12716 25644 12768 25696
rect 12900 25644 12952 25696
rect 17592 25712 17644 25764
rect 23664 25712 23716 25764
rect 18696 25644 18748 25696
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 11520 25440 11572 25492
rect 13268 25440 13320 25492
rect 16028 25440 16080 25492
rect 19524 25483 19576 25492
rect 19524 25449 19533 25483
rect 19533 25449 19567 25483
rect 19567 25449 19576 25483
rect 19524 25440 19576 25449
rect 20076 25440 20128 25492
rect 21640 25483 21692 25492
rect 21640 25449 21649 25483
rect 21649 25449 21683 25483
rect 21683 25449 21692 25483
rect 21640 25440 21692 25449
rect 28632 25483 28684 25492
rect 28632 25449 28641 25483
rect 28641 25449 28675 25483
rect 28675 25449 28684 25483
rect 28632 25440 28684 25449
rect 36268 25483 36320 25492
rect 36268 25449 36277 25483
rect 36277 25449 36311 25483
rect 36311 25449 36320 25483
rect 36268 25440 36320 25449
rect 11612 25372 11664 25424
rect 12532 25372 12584 25424
rect 12808 25372 12860 25424
rect 15844 25372 15896 25424
rect 8208 25304 8260 25356
rect 9956 25236 10008 25288
rect 13084 25304 13136 25356
rect 18144 25347 18196 25356
rect 18144 25313 18153 25347
rect 18153 25313 18187 25347
rect 18187 25313 18196 25347
rect 18144 25304 18196 25313
rect 38016 25347 38068 25356
rect 38016 25313 38025 25347
rect 38025 25313 38059 25347
rect 38059 25313 38068 25347
rect 38016 25304 38068 25313
rect 5540 25168 5592 25220
rect 7380 25211 7432 25220
rect 7380 25177 7389 25211
rect 7389 25177 7423 25211
rect 7423 25177 7432 25211
rect 7380 25168 7432 25177
rect 11152 25236 11204 25288
rect 13912 25236 13964 25288
rect 14924 25236 14976 25288
rect 11428 25211 11480 25220
rect 10968 25100 11020 25152
rect 11428 25177 11437 25211
rect 11437 25177 11471 25211
rect 11471 25177 11480 25211
rect 11428 25168 11480 25177
rect 12716 25211 12768 25220
rect 12716 25177 12725 25211
rect 12725 25177 12759 25211
rect 12759 25177 12768 25211
rect 12716 25168 12768 25177
rect 15016 25100 15068 25152
rect 15568 25100 15620 25152
rect 16028 25168 16080 25220
rect 16672 25168 16724 25220
rect 19892 25236 19944 25288
rect 19984 25236 20036 25288
rect 21456 25236 21508 25288
rect 18696 25211 18748 25220
rect 18696 25177 18705 25211
rect 18705 25177 18739 25211
rect 18739 25177 18748 25211
rect 18696 25168 18748 25177
rect 19340 25168 19392 25220
rect 36268 25236 36320 25288
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 37648 25168 37700 25220
rect 16212 25100 16264 25152
rect 18604 25100 18656 25152
rect 38016 25100 38068 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7380 24896 7432 24948
rect 13820 24896 13872 24948
rect 14924 24896 14976 24948
rect 38292 24939 38344 24948
rect 9864 24871 9916 24880
rect 9864 24837 9873 24871
rect 9873 24837 9907 24871
rect 9907 24837 9916 24871
rect 9864 24828 9916 24837
rect 2136 24760 2188 24812
rect 9956 24760 10008 24812
rect 10784 24760 10836 24812
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 11428 24828 11480 24880
rect 11980 24803 12032 24812
rect 10968 24760 11020 24769
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 14648 24871 14700 24880
rect 14648 24837 14657 24871
rect 14657 24837 14691 24871
rect 14691 24837 14700 24871
rect 14648 24828 14700 24837
rect 13912 24760 13964 24812
rect 38292 24905 38301 24939
rect 38301 24905 38335 24939
rect 38335 24905 38344 24939
rect 38292 24896 38344 24905
rect 12808 24735 12860 24744
rect 12808 24701 12817 24735
rect 12817 24701 12851 24735
rect 12851 24701 12860 24735
rect 12808 24692 12860 24701
rect 14280 24692 14332 24744
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 15844 24692 15896 24744
rect 16580 24760 16632 24812
rect 16672 24692 16724 24744
rect 2320 24624 2372 24676
rect 12716 24624 12768 24676
rect 13820 24624 13872 24676
rect 18144 24871 18196 24880
rect 18144 24837 18153 24871
rect 18153 24837 18187 24871
rect 18187 24837 18196 24871
rect 18144 24828 18196 24837
rect 18604 24828 18656 24880
rect 19340 24828 19392 24880
rect 19984 24760 20036 24812
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 17868 24692 17920 24744
rect 15108 24556 15160 24608
rect 16488 24556 16540 24608
rect 21456 24692 21508 24744
rect 32404 24692 32456 24744
rect 28540 24556 28592 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 5540 24352 5592 24404
rect 10876 24352 10928 24404
rect 13084 24352 13136 24404
rect 14556 24352 14608 24404
rect 15108 24352 15160 24404
rect 17960 24352 18012 24404
rect 20076 24352 20128 24404
rect 26884 24395 26936 24404
rect 26884 24361 26893 24395
rect 26893 24361 26927 24395
rect 26927 24361 26936 24395
rect 26884 24352 26936 24361
rect 2044 24216 2096 24268
rect 1860 24191 1912 24200
rect 1860 24157 1869 24191
rect 1869 24157 1903 24191
rect 1903 24157 1912 24191
rect 1860 24148 1912 24157
rect 4620 24148 4672 24200
rect 9036 24148 9088 24200
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 12808 24080 12860 24132
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 12716 24012 12768 24064
rect 15108 24216 15160 24268
rect 15200 24216 15252 24268
rect 16212 24216 16264 24268
rect 17776 24259 17828 24268
rect 17776 24225 17785 24259
rect 17785 24225 17819 24259
rect 17819 24225 17828 24259
rect 17776 24216 17828 24225
rect 14188 24148 14240 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 15016 24148 15068 24200
rect 13084 24123 13136 24132
rect 13084 24089 13093 24123
rect 13093 24089 13127 24123
rect 13127 24089 13136 24123
rect 13084 24080 13136 24089
rect 13176 24123 13228 24132
rect 13176 24089 13185 24123
rect 13185 24089 13219 24123
rect 13219 24089 13228 24123
rect 16672 24148 16724 24200
rect 13176 24080 13228 24089
rect 17776 24080 17828 24132
rect 19340 24080 19392 24132
rect 14464 24012 14516 24064
rect 20076 24055 20128 24064
rect 20076 24021 20085 24055
rect 20085 24021 20119 24055
rect 20119 24021 20128 24055
rect 20076 24012 20128 24021
rect 27528 24012 27580 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 12348 23808 12400 23860
rect 14188 23851 14240 23860
rect 14188 23817 14197 23851
rect 14197 23817 14231 23851
rect 14231 23817 14240 23851
rect 14188 23808 14240 23817
rect 17776 23808 17828 23860
rect 19340 23851 19392 23860
rect 15568 23783 15620 23792
rect 10416 23672 10468 23724
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 14648 23672 14700 23724
rect 15568 23749 15577 23783
rect 15577 23749 15611 23783
rect 15611 23749 15620 23783
rect 15568 23740 15620 23749
rect 16120 23783 16172 23792
rect 16120 23749 16129 23783
rect 16129 23749 16163 23783
rect 16163 23749 16172 23783
rect 16120 23740 16172 23749
rect 17040 23783 17092 23792
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 17592 23740 17644 23792
rect 19340 23817 19349 23851
rect 19349 23817 19383 23851
rect 19383 23817 19392 23851
rect 19340 23808 19392 23817
rect 17868 23672 17920 23724
rect 20076 23672 20128 23724
rect 38016 23715 38068 23724
rect 38016 23681 38025 23715
rect 38025 23681 38059 23715
rect 38059 23681 38068 23715
rect 38016 23672 38068 23681
rect 15292 23536 15344 23588
rect 15568 23604 15620 23656
rect 16948 23647 17000 23656
rect 16948 23613 16957 23647
rect 16957 23613 16991 23647
rect 16991 23613 17000 23647
rect 16948 23604 17000 23613
rect 12808 23468 12860 23520
rect 16672 23468 16724 23520
rect 18052 23536 18104 23588
rect 20352 23536 20404 23588
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 27528 23468 27580 23520
rect 29828 23468 29880 23520
rect 38200 23511 38252 23520
rect 38200 23477 38209 23511
rect 38209 23477 38243 23511
rect 38243 23477 38252 23511
rect 38200 23468 38252 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1860 23264 1912 23316
rect 13176 23264 13228 23316
rect 14556 23264 14608 23316
rect 11244 23196 11296 23248
rect 12900 23128 12952 23180
rect 14188 23128 14240 23180
rect 14832 23128 14884 23180
rect 14004 23060 14056 23112
rect 4620 22924 4672 22976
rect 16028 23196 16080 23248
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 16396 23128 16448 23180
rect 16948 23128 17000 23180
rect 18328 23060 18380 23112
rect 23388 23060 23440 23112
rect 15200 22992 15252 23044
rect 16028 23035 16080 23044
rect 16028 23001 16037 23035
rect 16037 23001 16071 23035
rect 16071 23001 16080 23035
rect 16028 22992 16080 23001
rect 17040 23035 17092 23044
rect 17040 23001 17049 23035
rect 17049 23001 17083 23035
rect 17083 23001 17092 23035
rect 17040 22992 17092 23001
rect 18052 23035 18104 23044
rect 18052 23001 18061 23035
rect 18061 23001 18095 23035
rect 18095 23001 18104 23035
rect 18052 22992 18104 23001
rect 28908 22992 28960 23044
rect 17684 22924 17736 22976
rect 18788 22924 18840 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 11336 22720 11388 22772
rect 13912 22720 13964 22772
rect 15936 22720 15988 22772
rect 18328 22720 18380 22772
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 14280 22652 14332 22704
rect 14924 22695 14976 22704
rect 14924 22661 14933 22695
rect 14933 22661 14967 22695
rect 14967 22661 14976 22695
rect 14924 22652 14976 22661
rect 15384 22652 15436 22704
rect 17960 22695 18012 22704
rect 17960 22661 17969 22695
rect 17969 22661 18003 22695
rect 18003 22661 18012 22695
rect 17960 22652 18012 22661
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 15200 22559 15252 22568
rect 15200 22525 15209 22559
rect 15209 22525 15243 22559
rect 15243 22525 15252 22559
rect 15200 22516 15252 22525
rect 14004 22448 14056 22500
rect 17684 22584 17736 22636
rect 27528 22720 27580 22772
rect 17960 22516 18012 22568
rect 18788 22516 18840 22568
rect 17040 22448 17092 22500
rect 17684 22448 17736 22500
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14556 22176 14608 22228
rect 18052 22176 18104 22228
rect 14280 22040 14332 22092
rect 16948 22040 17000 22092
rect 14556 21972 14608 22024
rect 14924 21972 14976 22024
rect 1676 21879 1728 21888
rect 1676 21845 1685 21879
rect 1685 21845 1719 21879
rect 1719 21845 1728 21879
rect 1676 21836 1728 21845
rect 14464 21836 14516 21888
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 17684 21904 17736 21956
rect 25320 22040 25372 22092
rect 38292 21972 38344 22024
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 37740 21879 37792 21888
rect 37740 21845 37749 21879
rect 37749 21845 37783 21879
rect 37783 21845 37792 21879
rect 37740 21836 37792 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 14372 21632 14424 21684
rect 14556 21632 14608 21684
rect 15384 21675 15436 21684
rect 15384 21641 15393 21675
rect 15393 21641 15427 21675
rect 15427 21641 15436 21675
rect 15384 21632 15436 21641
rect 17960 21632 18012 21684
rect 15108 21564 15160 21616
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 16580 21428 16632 21480
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 17776 21428 17828 21480
rect 16212 21360 16264 21412
rect 37924 21360 37976 21412
rect 18604 21335 18656 21344
rect 18604 21301 18613 21335
rect 18613 21301 18647 21335
rect 18647 21301 18656 21335
rect 18604 21292 18656 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13912 21088 13964 21140
rect 14924 21131 14976 21140
rect 14924 21097 14933 21131
rect 14933 21097 14967 21131
rect 14967 21097 14976 21131
rect 14924 21088 14976 21097
rect 16948 21131 17000 21140
rect 16948 21097 16957 21131
rect 16957 21097 16991 21131
rect 16991 21097 17000 21131
rect 16948 21088 17000 21097
rect 17776 21131 17828 21140
rect 17776 21097 17785 21131
rect 17785 21097 17819 21131
rect 17819 21097 17828 21131
rect 17776 21088 17828 21097
rect 14464 20884 14516 20936
rect 16580 20995 16632 21004
rect 16580 20961 16589 20995
rect 16589 20961 16623 20995
rect 16623 20961 16632 20995
rect 16580 20952 16632 20961
rect 18604 20952 18656 21004
rect 1584 20816 1636 20868
rect 11980 20816 12032 20868
rect 18696 20884 18748 20936
rect 11704 20748 11756 20800
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 15108 20544 15160 20596
rect 16948 20544 17000 20596
rect 17408 20544 17460 20596
rect 28908 20544 28960 20596
rect 38016 20587 38068 20596
rect 38016 20553 38025 20587
rect 38025 20553 38059 20587
rect 38059 20553 38068 20587
rect 38016 20544 38068 20553
rect 1584 20519 1636 20528
rect 1584 20485 1593 20519
rect 1593 20485 1627 20519
rect 1627 20485 1636 20519
rect 1584 20476 1636 20485
rect 11704 20476 11756 20528
rect 15108 20408 15160 20460
rect 15292 20340 15344 20392
rect 16028 20408 16080 20460
rect 17132 20408 17184 20460
rect 14464 20204 14516 20256
rect 16580 20204 16632 20256
rect 37832 20451 37884 20460
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 18788 20204 18840 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 15476 20000 15528 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17868 20000 17920 20052
rect 16580 19907 16632 19916
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 16488 19796 16540 19848
rect 15200 19660 15252 19712
rect 17684 19660 17736 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 17960 19499 18012 19508
rect 17960 19465 17969 19499
rect 17969 19465 18003 19499
rect 18003 19465 18012 19499
rect 17960 19456 18012 19465
rect 17684 19388 17736 19440
rect 24584 19388 24636 19440
rect 14556 19320 14608 19372
rect 17132 19363 17184 19372
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 19432 19320 19484 19372
rect 38200 19363 38252 19372
rect 38200 19329 38209 19363
rect 38209 19329 38243 19363
rect 38243 19329 38252 19363
rect 38200 19320 38252 19329
rect 37924 19252 37976 19304
rect 37740 19116 37792 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 17132 18912 17184 18964
rect 9128 18708 9180 18760
rect 1584 18640 1636 18692
rect 9772 18640 9824 18692
rect 2780 18572 2832 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19432 17824 19484 17876
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 12992 16940 13044 16992
rect 38016 16940 38068 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 15200 16396 15252 16448
rect 15384 16396 15436 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 10876 16124 10928 16176
rect 12900 16124 12952 16176
rect 9864 16099 9916 16108
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 12256 16056 12308 16108
rect 13728 16056 13780 16108
rect 23204 16056 23256 16108
rect 9404 15920 9456 15972
rect 15384 15920 15436 15972
rect 33692 15920 33744 15972
rect 7472 15852 7524 15904
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1860 15648 1912 15700
rect 9404 15648 9456 15700
rect 9864 15648 9916 15700
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 16396 15648 16448 15700
rect 16396 15444 16448 15496
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 17684 14220 17736 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 37832 13880 37884 13932
rect 38292 13855 38344 13864
rect 38292 13821 38301 13855
rect 38301 13821 38335 13855
rect 38335 13821 38344 13855
rect 38292 13812 38344 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 38292 13515 38344 13524
rect 38292 13481 38301 13515
rect 38301 13481 38335 13515
rect 38335 13481 38344 13515
rect 38292 13472 38344 13481
rect 2780 13268 2832 13320
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 38200 11747 38252 11756
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 20076 11500 20128 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 16488 11339 16540 11348
rect 16488 11305 16497 11339
rect 16497 11305 16531 11339
rect 16531 11305 16540 11339
rect 16488 11296 16540 11305
rect 20444 11160 20496 11212
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 17132 11024 17184 11033
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 15016 10795 15068 10804
rect 15016 10761 15025 10795
rect 15025 10761 15059 10795
rect 15059 10761 15068 10795
rect 15016 10752 15068 10761
rect 17224 10795 17276 10804
rect 17224 10761 17233 10795
rect 17233 10761 17267 10795
rect 17267 10761 17276 10795
rect 17224 10752 17276 10761
rect 18788 10795 18840 10804
rect 18788 10761 18797 10795
rect 18797 10761 18831 10795
rect 18831 10761 18840 10795
rect 18788 10752 18840 10761
rect 15660 10616 15712 10668
rect 17408 10616 17460 10668
rect 38200 10659 38252 10668
rect 38200 10625 38209 10659
rect 38209 10625 38243 10659
rect 38243 10625 38252 10659
rect 38200 10616 38252 10625
rect 16396 10480 16448 10532
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 16396 10208 16448 10260
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 16764 9596 16816 9648
rect 17500 9528 17552 9580
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 14372 8916 14424 8968
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 38108 8619 38160 8628
rect 38108 8585 38117 8619
rect 38117 8585 38151 8619
rect 38151 8585 38160 8619
rect 38108 8576 38160 8585
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 23204 8007 23256 8016
rect 23204 7973 23213 8007
rect 23213 7973 23247 8007
rect 23247 7973 23256 8007
rect 23204 7964 23256 7973
rect 10600 7760 10652 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1584 7352 1636 7404
rect 14464 7148 14516 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 38016 6375 38068 6384
rect 38016 6341 38025 6375
rect 38025 6341 38059 6375
rect 38059 6341 38068 6375
rect 38016 6332 38068 6341
rect 38200 6307 38252 6316
rect 38200 6273 38209 6307
rect 38209 6273 38243 6307
rect 38243 6273 38252 6307
rect 38200 6264 38252 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37648 4700 37700 4752
rect 38200 4539 38252 4548
rect 38200 4505 38209 4539
rect 38209 4505 38243 4539
rect 38243 4505 38252 4539
rect 38200 4496 38252 4505
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 12808 3476 12860 3528
rect 15660 3408 15712 3460
rect 16028 3408 16080 3460
rect 21364 3408 21416 3460
rect 23756 3408 23808 3460
rect 36728 3476 36780 3528
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 17224 3340 17276 3392
rect 17500 3340 17552 3392
rect 38660 3408 38712 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5540 3136 5592 3188
rect 19432 3136 19484 3188
rect 24768 3136 24820 3188
rect 16304 3068 16356 3120
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 14556 3043 14608 3052
rect 12992 3000 13044 3009
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 17408 3043 17460 3052
rect 14188 2932 14240 2984
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 21364 3068 21416 3120
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 17224 2932 17276 2984
rect 17868 2932 17920 2984
rect 31024 2932 31076 2984
rect 34428 2864 34480 2916
rect 38108 2864 38160 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 10508 2796 10560 2848
rect 17500 2796 17552 2848
rect 19708 2796 19760 2848
rect 23572 2839 23624 2848
rect 23572 2805 23581 2839
rect 23581 2805 23615 2839
rect 23615 2805 23624 2839
rect 23572 2796 23624 2805
rect 27160 2796 27212 2848
rect 29644 2839 29696 2848
rect 29644 2805 29653 2839
rect 29653 2805 29687 2839
rect 29687 2805 29696 2839
rect 29644 2796 29696 2805
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 12992 2592 13044 2644
rect 17132 2592 17184 2644
rect 28540 2635 28592 2644
rect 20 2524 72 2576
rect 4620 2456 4672 2508
rect 8852 2456 8904 2508
rect 2320 2388 2372 2440
rect 2780 2388 2832 2440
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 5172 2252 5224 2304
rect 7104 2252 7156 2304
rect 8392 2252 8444 2304
rect 10324 2388 10376 2440
rect 23572 2524 23624 2576
rect 15476 2456 15528 2508
rect 19984 2456 20036 2508
rect 28540 2601 28549 2635
rect 28549 2601 28583 2635
rect 28583 2601 28592 2635
rect 28540 2592 28592 2601
rect 29828 2635 29880 2644
rect 29828 2601 29837 2635
rect 29837 2601 29871 2635
rect 29871 2601 29880 2635
rect 29828 2592 29880 2601
rect 32404 2635 32456 2644
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 33692 2635 33744 2644
rect 33692 2601 33701 2635
rect 33701 2601 33735 2635
rect 33735 2601 33744 2635
rect 33692 2592 33744 2601
rect 36728 2635 36780 2644
rect 36728 2601 36737 2635
rect 36737 2601 36771 2635
rect 36771 2601 36780 2635
rect 36728 2592 36780 2601
rect 31024 2524 31076 2576
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18328 2388 18380 2440
rect 19708 2388 19760 2440
rect 24492 2388 24544 2440
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 34428 2388 34480 2440
rect 36728 2388 36780 2440
rect 28356 2320 28408 2372
rect 29644 2320 29696 2372
rect 33508 2320 33560 2372
rect 38200 2363 38252 2372
rect 38200 2329 38209 2363
rect 38209 2329 38243 2363
rect 38243 2329 38252 2363
rect 38200 2320 38252 2329
rect 12256 2252 12308 2304
rect 17408 2252 17460 2304
rect 19340 2252 19392 2304
rect 21272 2252 21324 2304
rect 22560 2252 22612 2304
rect 26424 2252 26476 2304
rect 31760 2295 31812 2304
rect 31760 2261 31769 2295
rect 31769 2261 31803 2295
rect 31803 2261 31812 2295
rect 31760 2252 31812 2261
rect 35440 2252 35492 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 2594 39200 2650 39800
rect 3882 39200 3938 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 676 35290 704 39200
rect 2504 37188 2556 37194
rect 2504 37130 2556 37136
rect 1492 37120 1544 37126
rect 1492 37062 1544 37068
rect 664 35284 716 35290
rect 664 35226 716 35232
rect 1504 31278 1532 37062
rect 1582 36816 1638 36825
rect 1582 36751 1584 36760
rect 1636 36751 1638 36760
rect 1584 36722 1636 36728
rect 1492 31272 1544 31278
rect 1492 31214 1544 31220
rect 1596 27606 1624 36722
rect 2136 36712 2188 36718
rect 2136 36654 2188 36660
rect 1950 36272 2006 36281
rect 1950 36207 2006 36216
rect 1964 36106 1992 36207
rect 1952 36100 2004 36106
rect 1952 36042 2004 36048
rect 1964 35766 1992 36042
rect 1952 35760 2004 35766
rect 1952 35702 2004 35708
rect 1860 34944 1912 34950
rect 1912 34904 1992 34932
rect 1860 34886 1912 34892
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34066 1716 34342
rect 1676 34060 1728 34066
rect 1676 34002 1728 34008
rect 1860 32768 1912 32774
rect 1860 32710 1912 32716
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31482 1716 31758
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29345 1716 29446
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1872 28422 1900 32710
rect 1964 31890 1992 34904
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2056 33697 2084 34682
rect 2042 33688 2098 33697
rect 2042 33623 2098 33632
rect 2056 33590 2084 33623
rect 2044 33584 2096 33590
rect 2044 33526 2096 33532
rect 2044 33312 2096 33318
rect 2044 33254 2096 33260
rect 1952 31884 2004 31890
rect 1952 31826 2004 31832
rect 1964 30394 1992 31826
rect 2056 30938 2084 33254
rect 2044 30932 2096 30938
rect 2044 30874 2096 30880
rect 1952 30388 2004 30394
rect 1952 30330 2004 30336
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 2056 29034 2084 29582
rect 2044 29028 2096 29034
rect 2044 28970 2096 28976
rect 1860 28416 1912 28422
rect 1860 28358 1912 28364
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1584 27600 1636 27606
rect 1584 27542 1636 27548
rect 1872 26382 1900 28358
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1676 26240 1728 26246
rect 1676 26182 1728 26188
rect 1688 25945 1716 26182
rect 1674 25936 1730 25945
rect 1674 25871 1730 25880
rect 2056 24274 2084 28970
rect 2148 26314 2176 36654
rect 2228 35760 2280 35766
rect 2228 35702 2280 35708
rect 2240 28694 2268 35702
rect 2412 34740 2464 34746
rect 2412 34682 2464 34688
rect 2320 33448 2372 33454
rect 2320 33390 2372 33396
rect 2332 29306 2360 33390
rect 2424 32366 2452 34682
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 2424 29510 2452 32302
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2516 29306 2544 37130
rect 2608 36378 2636 39200
rect 3896 37262 3924 39200
rect 4066 38856 4122 38865
rect 4066 38791 4122 38800
rect 3884 37256 3936 37262
rect 3884 37198 3936 37204
rect 3148 37188 3200 37194
rect 3148 37130 3200 37136
rect 2596 36372 2648 36378
rect 2596 36314 2648 36320
rect 3056 36168 3108 36174
rect 3056 36110 3108 36116
rect 2688 35012 2740 35018
rect 2688 34954 2740 34960
rect 2596 33516 2648 33522
rect 2596 33458 2648 33464
rect 2320 29300 2372 29306
rect 2320 29242 2372 29248
rect 2504 29300 2556 29306
rect 2504 29242 2556 29248
rect 2608 28694 2636 33458
rect 2700 29850 2728 34954
rect 2964 33924 3016 33930
rect 2964 33866 3016 33872
rect 2872 32496 2924 32502
rect 2872 32438 2924 32444
rect 2780 32428 2832 32434
rect 2780 32370 2832 32376
rect 2792 31385 2820 32370
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 2792 28762 2820 31311
rect 2884 30190 2912 32438
rect 2976 30938 3004 33866
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 3068 30818 3096 36110
rect 3160 33454 3188 37130
rect 3896 36922 3924 37198
rect 3884 36916 3936 36922
rect 3884 36858 3936 36864
rect 3608 36712 3660 36718
rect 3608 36654 3660 36660
rect 3424 35012 3476 35018
rect 3424 34954 3476 34960
rect 3148 33448 3200 33454
rect 3148 33390 3200 33396
rect 3240 32768 3292 32774
rect 3160 32728 3240 32756
rect 3160 30938 3188 32728
rect 3240 32710 3292 32716
rect 3436 32314 3464 34954
rect 3516 34536 3568 34542
rect 3516 34478 3568 34484
rect 3252 32286 3464 32314
rect 3252 31754 3280 32286
rect 3422 31920 3478 31929
rect 3422 31855 3424 31864
rect 3476 31855 3478 31864
rect 3424 31826 3476 31832
rect 3252 31726 3372 31754
rect 3148 30932 3200 30938
rect 3148 30874 3200 30880
rect 3068 30790 3188 30818
rect 3160 30326 3188 30790
rect 3240 30728 3292 30734
rect 3240 30670 3292 30676
rect 3252 30598 3280 30670
rect 3240 30592 3292 30598
rect 3240 30534 3292 30540
rect 3148 30320 3200 30326
rect 3148 30262 3200 30268
rect 3252 30258 3280 30534
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 3252 29646 3280 30194
rect 3344 29714 3372 31726
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3332 29708 3384 29714
rect 3332 29650 3384 29656
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 2976 28966 3004 29174
rect 3252 29170 3280 29582
rect 3436 29170 3464 30670
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3424 29164 3476 29170
rect 3424 29106 3476 29112
rect 2964 28960 3016 28966
rect 2964 28902 3016 28908
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2228 28688 2280 28694
rect 2228 28630 2280 28636
rect 2596 28688 2648 28694
rect 2596 28630 2648 28636
rect 3252 28558 3280 29106
rect 3436 29034 3464 29106
rect 3424 29028 3476 29034
rect 3424 28970 3476 28976
rect 3436 28558 3464 28970
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3424 28552 3476 28558
rect 3424 28494 3476 28500
rect 2792 28082 2820 28494
rect 3436 28082 3464 28494
rect 3528 28218 3556 34478
rect 3620 33590 3648 36654
rect 3896 36242 3924 36858
rect 3884 36236 3936 36242
rect 3884 36178 3936 36184
rect 3896 35714 3924 36178
rect 4080 35834 4108 38791
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4528 37324 4580 37330
rect 4528 37266 4580 37272
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 4540 37210 4568 37266
rect 4540 37182 4660 37210
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 3896 35698 4016 35714
rect 3896 35692 4028 35698
rect 3896 35686 3976 35692
rect 3896 35154 3924 35686
rect 3976 35634 4028 35640
rect 4632 35562 4660 37182
rect 5448 37188 5500 37194
rect 5448 37130 5500 37136
rect 4896 36916 4948 36922
rect 4896 36858 4948 36864
rect 4908 36786 4936 36858
rect 4896 36780 4948 36786
rect 4896 36722 4948 36728
rect 5460 36310 5488 37130
rect 5540 36712 5592 36718
rect 5538 36680 5540 36689
rect 5592 36680 5594 36689
rect 5538 36615 5594 36624
rect 5448 36304 5500 36310
rect 5448 36246 5500 36252
rect 5448 36168 5500 36174
rect 5078 36136 5134 36145
rect 5448 36110 5500 36116
rect 5078 36071 5080 36080
rect 5132 36071 5134 36080
rect 5080 36042 5132 36048
rect 4620 35556 4672 35562
rect 4620 35498 4672 35504
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3884 35148 3936 35154
rect 3884 35090 3936 35096
rect 3700 34944 3752 34950
rect 3700 34886 3752 34892
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 3620 32774 3648 33526
rect 3608 32768 3660 32774
rect 3608 32710 3660 32716
rect 3608 31748 3660 31754
rect 3608 31690 3660 31696
rect 3620 29714 3648 31690
rect 3712 31142 3740 34886
rect 3896 34746 3924 35090
rect 4724 35086 4752 35430
rect 4712 35080 4764 35086
rect 4712 35022 4764 35028
rect 3884 34740 3936 34746
rect 3884 34682 3936 34688
rect 3896 34406 3924 34682
rect 5172 34672 5224 34678
rect 5172 34614 5224 34620
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 3884 34400 3936 34406
rect 3884 34342 3936 34348
rect 4620 34400 4672 34406
rect 4620 34342 4672 34348
rect 3896 34066 3924 34342
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 3792 34060 3844 34066
rect 3792 34002 3844 34008
rect 3884 34060 3936 34066
rect 3884 34002 3936 34008
rect 3804 33658 3832 34002
rect 3792 33652 3844 33658
rect 3792 33594 3844 33600
rect 3896 33504 3924 34002
rect 4436 33992 4488 33998
rect 4436 33934 4488 33940
rect 4448 33522 4476 33934
rect 3976 33516 4028 33522
rect 3896 33476 3976 33504
rect 3896 32978 3924 33476
rect 3976 33458 4028 33464
rect 4436 33516 4488 33522
rect 4436 33458 4488 33464
rect 4066 33416 4122 33425
rect 4066 33351 4122 33360
rect 4080 33114 4108 33351
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3884 32972 3936 32978
rect 3884 32914 3936 32920
rect 3896 32570 3924 32914
rect 4632 32910 4660 34342
rect 4712 33448 4764 33454
rect 4712 33390 4764 33396
rect 4620 32904 4672 32910
rect 4620 32846 4672 32852
rect 4344 32836 4396 32842
rect 4344 32778 4396 32784
rect 3884 32564 3936 32570
rect 3884 32506 3936 32512
rect 3896 31754 3924 32506
rect 4356 32366 4384 32778
rect 4620 32496 4672 32502
rect 4620 32438 4672 32444
rect 4344 32360 4396 32366
rect 4344 32302 4396 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4080 31890 4200 31906
rect 4080 31884 4212 31890
rect 4080 31878 4160 31884
rect 4080 31754 4108 31878
rect 4160 31826 4212 31832
rect 3896 31726 4108 31754
rect 3896 31482 3924 31726
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 4172 31482 4200 31622
rect 3884 31476 3936 31482
rect 3884 31418 3936 31424
rect 4160 31476 4212 31482
rect 4160 31418 4212 31424
rect 3792 31408 3844 31414
rect 4632 31385 4660 32438
rect 3792 31350 3844 31356
rect 4618 31376 4674 31385
rect 3700 31136 3752 31142
rect 3700 31078 3752 31084
rect 3804 30326 3832 31350
rect 4618 31311 4674 31320
rect 4632 31278 4660 31311
rect 4620 31272 4672 31278
rect 3882 31240 3938 31249
rect 4620 31214 4672 31220
rect 3882 31175 3938 31184
rect 3896 31142 3924 31175
rect 3884 31136 3936 31142
rect 3884 31078 3936 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4528 30864 4580 30870
rect 4528 30806 4580 30812
rect 3792 30320 3844 30326
rect 3792 30262 3844 30268
rect 4540 30258 4568 30806
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3608 29708 3660 29714
rect 3608 29650 3660 29656
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28218 4660 31214
rect 4724 30258 4752 33390
rect 4816 32502 4844 34478
rect 5184 34184 5212 34614
rect 5000 34156 5212 34184
rect 4804 32496 4856 32502
rect 4804 32438 4856 32444
rect 5000 32314 5028 34156
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5080 33924 5132 33930
rect 5080 33866 5132 33872
rect 4816 32286 5028 32314
rect 4712 30252 4764 30258
rect 4712 30194 4764 30200
rect 4724 29646 4752 30194
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 4724 29170 4752 29582
rect 4816 29238 4844 32286
rect 4894 32192 4950 32201
rect 4894 32127 4950 32136
rect 4908 29850 4936 32127
rect 5092 30598 5120 33866
rect 5184 32978 5212 34002
rect 5172 32972 5224 32978
rect 5172 32914 5224 32920
rect 5172 32836 5224 32842
rect 5172 32778 5224 32784
rect 5184 32201 5212 32778
rect 5264 32428 5316 32434
rect 5264 32370 5316 32376
rect 5170 32192 5226 32201
rect 5170 32127 5226 32136
rect 5276 31804 5304 32370
rect 5184 31776 5304 31804
rect 5184 31686 5212 31776
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5184 30870 5212 31622
rect 5354 31512 5410 31521
rect 5354 31447 5410 31456
rect 5264 31272 5316 31278
rect 5264 31214 5316 31220
rect 5276 30870 5304 31214
rect 5172 30864 5224 30870
rect 5172 30806 5224 30812
rect 5264 30864 5316 30870
rect 5264 30806 5316 30812
rect 5184 30734 5212 30806
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 5080 30592 5132 30598
rect 5080 30534 5132 30540
rect 4896 29844 4948 29850
rect 4896 29786 4948 29792
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4712 29164 4764 29170
rect 4712 29106 4764 29112
rect 4724 28558 4752 29106
rect 5368 28762 5396 31447
rect 5460 30326 5488 36110
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5552 35698 5580 35974
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5644 35154 5672 37266
rect 5828 37126 5856 39200
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 6000 37256 6052 37262
rect 6000 37198 6052 37204
rect 7196 37256 7248 37262
rect 7196 37198 7248 37204
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5828 36854 5856 37062
rect 6012 36922 6040 37198
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 5816 36848 5868 36854
rect 5816 36790 5868 36796
rect 6184 36848 6236 36854
rect 6184 36790 6236 36796
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 5632 35148 5684 35154
rect 5632 35090 5684 35096
rect 5540 34740 5592 34746
rect 5540 34682 5592 34688
rect 5552 33318 5580 34682
rect 5736 34184 5764 36722
rect 6000 35760 6052 35766
rect 6000 35702 6052 35708
rect 6092 35760 6144 35766
rect 6092 35702 6144 35708
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5920 34542 5948 35430
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5736 34156 5856 34184
rect 5724 33924 5776 33930
rect 5724 33866 5776 33872
rect 5632 33448 5684 33454
rect 5632 33390 5684 33396
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5644 32434 5672 33390
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 5644 31346 5672 32166
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5736 31226 5764 33866
rect 5644 31198 5764 31226
rect 5644 30938 5672 31198
rect 5724 31136 5776 31142
rect 5724 31078 5776 31084
rect 5736 30938 5764 31078
rect 5632 30932 5684 30938
rect 5632 30874 5684 30880
rect 5724 30932 5776 30938
rect 5724 30874 5776 30880
rect 5724 30728 5776 30734
rect 5724 30670 5776 30676
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5736 30258 5764 30670
rect 5828 30326 5856 34156
rect 5908 32564 5960 32570
rect 5908 32506 5960 32512
rect 5920 31686 5948 32506
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 6012 31346 6040 35702
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 5816 30320 5868 30326
rect 5816 30262 5868 30268
rect 5724 30252 5776 30258
rect 5724 30194 5776 30200
rect 6104 29782 6132 35702
rect 6196 31521 6224 36790
rect 7024 36718 7052 37130
rect 7208 36938 7236 37198
rect 7116 36910 7236 36938
rect 6552 36712 6604 36718
rect 6552 36654 6604 36660
rect 7012 36712 7064 36718
rect 7012 36654 7064 36660
rect 6460 36644 6512 36650
rect 6460 36586 6512 36592
rect 6276 31952 6328 31958
rect 6276 31894 6328 31900
rect 6288 31822 6316 31894
rect 6276 31816 6328 31822
rect 6276 31758 6328 31764
rect 6368 31748 6420 31754
rect 6368 31690 6420 31696
rect 6182 31512 6238 31521
rect 6182 31447 6238 31456
rect 6182 31240 6238 31249
rect 6182 31175 6238 31184
rect 6196 31142 6224 31175
rect 6184 31136 6236 31142
rect 6184 31078 6236 31084
rect 6380 30818 6408 31690
rect 6288 30790 6408 30818
rect 6092 29776 6144 29782
rect 6092 29718 6144 29724
rect 6288 28762 6316 30790
rect 6472 30054 6500 36586
rect 6564 33658 6592 36654
rect 6828 36168 6880 36174
rect 6828 36110 6880 36116
rect 6644 36100 6696 36106
rect 6644 36042 6696 36048
rect 6656 33998 6684 36042
rect 6840 35630 6868 36110
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6840 35154 6868 35566
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6552 33652 6604 33658
rect 6552 33594 6604 33600
rect 6840 33522 6868 34478
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6840 33130 6868 33458
rect 6932 33318 6960 34342
rect 7012 33516 7064 33522
rect 7012 33458 7064 33464
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 6840 33102 6960 33130
rect 6932 33046 6960 33102
rect 6920 33040 6972 33046
rect 6920 32982 6972 32988
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6748 32230 6776 32438
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6644 31952 6696 31958
rect 6550 31920 6606 31929
rect 6644 31894 6696 31900
rect 6550 31855 6552 31864
rect 6604 31855 6606 31864
rect 6552 31826 6604 31832
rect 6656 31754 6684 31894
rect 6564 31726 6684 31754
rect 6460 30048 6512 30054
rect 6460 29990 6512 29996
rect 6564 29306 6592 31726
rect 6748 31482 6776 32166
rect 6840 31822 6868 32846
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 6644 30796 6696 30802
rect 6644 30738 6696 30744
rect 6656 30410 6684 30738
rect 6748 30546 6776 31282
rect 6840 30802 6868 31758
rect 6920 31204 6972 31210
rect 6920 31146 6972 31152
rect 6932 30802 6960 31146
rect 6828 30796 6880 30802
rect 6828 30738 6880 30744
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 6920 30592 6972 30598
rect 6748 30540 6920 30546
rect 6748 30534 6972 30540
rect 6748 30518 6960 30534
rect 6656 30382 6776 30410
rect 6748 30326 6776 30382
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6736 30048 6788 30054
rect 6736 29990 6788 29996
rect 6748 29646 6776 29990
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6552 29300 6604 29306
rect 6552 29242 6604 29248
rect 6840 29238 6868 30126
rect 6828 29232 6880 29238
rect 6828 29174 6880 29180
rect 7024 29102 7052 33458
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 5356 28756 5408 28762
rect 5356 28698 5408 28704
rect 6276 28756 6328 28762
rect 6276 28698 6328 28704
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 4620 28212 4672 28218
rect 4620 28154 4672 28160
rect 7116 28150 7144 36910
rect 7194 36680 7250 36689
rect 7194 36615 7250 36624
rect 7208 36582 7236 36615
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7300 35630 7328 37402
rect 7760 36174 7788 39200
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8760 37256 8812 37262
rect 8760 37198 8812 37204
rect 8588 36922 8616 37198
rect 8576 36916 8628 36922
rect 8576 36858 8628 36864
rect 8588 36718 8616 36858
rect 8300 36712 8352 36718
rect 8300 36654 8352 36660
rect 8576 36712 8628 36718
rect 8576 36654 8628 36660
rect 8668 36712 8720 36718
rect 8668 36654 8720 36660
rect 8312 36310 8340 36654
rect 8300 36304 8352 36310
rect 8300 36246 8352 36252
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7930 36136 7986 36145
rect 7288 35624 7340 35630
rect 7288 35566 7340 35572
rect 7760 35290 7788 36110
rect 7930 36071 7986 36080
rect 7944 36038 7972 36071
rect 7932 36032 7984 36038
rect 7932 35974 7984 35980
rect 8208 35624 8260 35630
rect 8208 35566 8260 35572
rect 8220 35465 8248 35566
rect 8206 35456 8262 35465
rect 8206 35391 8262 35400
rect 8312 35306 8340 36246
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 8220 35278 8340 35306
rect 8220 34082 8248 35278
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8312 34202 8340 35090
rect 8404 34474 8432 35566
rect 8392 34468 8444 34474
rect 8392 34410 8444 34416
rect 8300 34196 8352 34202
rect 8352 34156 8432 34184
rect 8300 34138 8352 34144
rect 8220 34054 8340 34082
rect 8404 34066 8432 34156
rect 8208 33924 8260 33930
rect 8208 33866 8260 33872
rect 7472 33856 7524 33862
rect 7472 33798 7524 33804
rect 7564 33856 7616 33862
rect 7564 33798 7616 33804
rect 7484 33454 7512 33798
rect 7576 33697 7604 33798
rect 7562 33688 7618 33697
rect 7562 33623 7618 33632
rect 7748 33652 7800 33658
rect 7748 33594 7800 33600
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7760 33318 7788 33594
rect 7656 33312 7708 33318
rect 7656 33254 7708 33260
rect 7748 33312 7800 33318
rect 7748 33254 7800 33260
rect 7196 32496 7248 32502
rect 7196 32438 7248 32444
rect 7208 28762 7236 32438
rect 7288 31476 7340 31482
rect 7288 31418 7340 31424
rect 7300 31385 7328 31418
rect 7286 31376 7342 31385
rect 7286 31311 7342 31320
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7300 29306 7328 29786
rect 7288 29300 7340 29306
rect 7288 29242 7340 29248
rect 7300 28762 7328 29242
rect 7668 28994 7696 33254
rect 7748 33040 7800 33046
rect 7748 32982 7800 32988
rect 7760 29850 7788 32982
rect 8220 32026 8248 33866
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8312 31754 8340 34054
rect 8392 34060 8444 34066
rect 8392 34002 8444 34008
rect 8404 33522 8432 34002
rect 8392 33516 8444 33522
rect 8392 33458 8444 33464
rect 8312 31726 8432 31754
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 8036 30870 8064 31350
rect 8024 30864 8076 30870
rect 8024 30806 8076 30812
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8128 30394 8156 30670
rect 8300 30592 8352 30598
rect 8300 30534 8352 30540
rect 8116 30388 8168 30394
rect 8116 30330 8168 30336
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 8220 29102 8248 29990
rect 8312 29238 8340 30534
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 8208 29096 8260 29102
rect 8208 29038 8260 29044
rect 7576 28966 7696 28994
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7300 28558 7328 28698
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7300 28218 7328 28494
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 7392 28014 7420 28358
rect 7576 28150 7604 28966
rect 7564 28144 7616 28150
rect 7564 28086 7616 28092
rect 7380 28008 7432 28014
rect 7380 27950 7432 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2136 26308 2188 26314
rect 2136 26250 2188 26256
rect 2148 24818 2176 26250
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 8220 25362 8248 29038
rect 8404 27130 8432 31726
rect 8496 28626 8524 36110
rect 8588 35154 8616 36654
rect 8576 35148 8628 35154
rect 8576 35090 8628 35096
rect 8576 35012 8628 35018
rect 8576 34954 8628 34960
rect 8588 33114 8616 34954
rect 8680 33590 8708 36654
rect 8668 33584 8720 33590
rect 8668 33526 8720 33532
rect 8772 33402 8800 37198
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9036 35624 9088 35630
rect 9036 35566 9088 35572
rect 9048 35154 9076 35566
rect 9036 35148 9088 35154
rect 9036 35090 9088 35096
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8864 34406 8892 34886
rect 9048 34746 9076 35090
rect 9140 35018 9168 37062
rect 9220 36848 9272 36854
rect 9220 36790 9272 36796
rect 9232 36174 9260 36790
rect 9312 36712 9364 36718
rect 9312 36654 9364 36660
rect 9324 36281 9352 36654
rect 9588 36304 9640 36310
rect 9310 36272 9366 36281
rect 9588 36246 9640 36252
rect 9310 36207 9366 36216
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 9496 36168 9548 36174
rect 9496 36110 9548 36116
rect 9220 36032 9272 36038
rect 9220 35974 9272 35980
rect 9128 35012 9180 35018
rect 9232 35000 9260 35974
rect 9404 35012 9456 35018
rect 9232 34972 9404 35000
rect 9128 34954 9180 34960
rect 9404 34954 9456 34960
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 9312 33924 9364 33930
rect 9312 33866 9364 33872
rect 9324 33658 9352 33866
rect 9128 33652 9180 33658
rect 9128 33594 9180 33600
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9036 33584 9088 33590
rect 8956 33544 9036 33572
rect 8852 33516 8904 33522
rect 8852 33458 8904 33464
rect 8680 33374 8800 33402
rect 8576 33108 8628 33114
rect 8576 33050 8628 33056
rect 8576 32360 8628 32366
rect 8576 32302 8628 32308
rect 8588 31890 8616 32302
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8680 30258 8708 33374
rect 8864 33114 8892 33458
rect 8852 33108 8904 33114
rect 8852 33050 8904 33056
rect 8760 32836 8812 32842
rect 8760 32778 8812 32784
rect 8772 31754 8800 32778
rect 8864 32434 8892 33050
rect 8852 32428 8904 32434
rect 8852 32370 8904 32376
rect 8864 32026 8892 32370
rect 8852 32020 8904 32026
rect 8852 31962 8904 31968
rect 8772 31726 8892 31754
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 8772 31142 8800 31282
rect 8760 31136 8812 31142
rect 8760 31078 8812 31084
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 5540 25220 5592 25226
rect 5540 25162 5592 25168
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2320 24676 2372 24682
rect 2320 24618 2372 24624
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23905 1716 24006
rect 1674 23896 1730 23905
rect 1674 23831 1730 23840
rect 1872 23322 1900 24142
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1676 21888 1728 21894
rect 1674 21856 1676 21865
rect 1728 21856 1730 21865
rect 1674 21791 1730 21800
rect 1584 20868 1636 20874
rect 1584 20810 1636 20816
rect 1596 20534 1624 20810
rect 1584 20528 1636 20534
rect 1582 20496 1584 20505
rect 1636 20496 1638 20505
rect 1582 20431 1638 20440
rect 1584 18692 1636 18698
rect 1584 18634 1636 18640
rect 1596 18465 1624 18634
rect 1582 18456 1638 18465
rect 1582 18391 1584 18400
rect 1636 18391 1638 18400
rect 1584 18362 1636 18368
rect 1676 16448 1728 16454
rect 1674 16416 1676 16425
rect 1728 16416 1730 16425
rect 1674 16351 1730 16360
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1674 14376 1730 14385
rect 1674 14311 1676 14320
rect 1728 14311 1730 14320
rect 1676 14282 1728 14288
rect 1688 14074 1716 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 13025 1716 13126
rect 1674 13016 1730 13025
rect 1674 12951 1730 12960
rect 1676 11008 1728 11014
rect 1674 10976 1676 10985
rect 1728 10976 1730 10985
rect 1674 10911 1730 10920
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 1688 8838 1716 8871
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1872 5710 1900 15642
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1676 5568 1728 5574
rect 1674 5536 1676 5545
rect 1728 5536 1730 5545
rect 1674 5471 1730 5480
rect 2332 3738 2360 24618
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 5552 24410 5580 25162
rect 7392 24954 7420 25162
rect 7380 24948 7432 24954
rect 7380 24890 7432 24896
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 22982 4660 24142
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 13326 2820 18566
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2332 2446 2360 3674
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2446 2820 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 22918
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 5552 2446 5580 3130
rect 7484 2446 7512 15846
rect 8864 2514 8892 31726
rect 8956 31210 8984 33544
rect 9036 33526 9088 33532
rect 9140 33402 9168 33594
rect 9048 33374 9168 33402
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 9048 24206 9076 33374
rect 9232 30258 9260 33390
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 9324 31278 9352 31962
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 9140 28490 9168 29038
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 9140 27402 9168 28426
rect 9128 27396 9180 27402
rect 9128 27338 9180 27344
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9140 18766 9168 27338
rect 9416 26450 9444 34954
rect 9508 30122 9536 36110
rect 9600 35766 9628 36246
rect 9588 35760 9640 35766
rect 9588 35702 9640 35708
rect 9692 35562 9720 39200
rect 10140 37460 10192 37466
rect 10140 37402 10192 37408
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 9954 35728 10010 35737
rect 9954 35663 9956 35672
rect 10008 35663 10010 35672
rect 9956 35634 10008 35640
rect 9680 35556 9732 35562
rect 9680 35498 9732 35504
rect 9864 35012 9916 35018
rect 9784 34972 9864 35000
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9600 33114 9628 33390
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9600 27402 9628 30534
rect 9692 28490 9720 31078
rect 9784 29034 9812 34972
rect 9864 34954 9916 34960
rect 9956 34536 10008 34542
rect 10008 34496 10088 34524
rect 9956 34478 10008 34484
rect 9956 34400 10008 34406
rect 9956 34342 10008 34348
rect 9864 33924 9916 33930
rect 9864 33866 9916 33872
rect 9772 29028 9824 29034
rect 9772 28970 9824 28976
rect 9876 28694 9904 33866
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9968 28558 9996 34342
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 10060 27962 10088 34496
rect 10152 32978 10180 37402
rect 10508 37324 10560 37330
rect 10508 37266 10560 37272
rect 10520 37074 10548 37266
rect 10600 37188 10652 37194
rect 10600 37130 10652 37136
rect 10428 37046 10548 37074
rect 10428 35222 10456 37046
rect 10612 36938 10640 37130
rect 10784 37120 10836 37126
rect 10784 37062 10836 37068
rect 10520 36910 10640 36938
rect 10796 36922 10824 37062
rect 10784 36916 10836 36922
rect 10520 36718 10548 36910
rect 10784 36858 10836 36864
rect 10600 36848 10652 36854
rect 10652 36796 10732 36802
rect 10600 36790 10732 36796
rect 10612 36774 10732 36790
rect 10508 36712 10560 36718
rect 10508 36654 10560 36660
rect 10416 35216 10468 35222
rect 10416 35158 10468 35164
rect 10704 35034 10732 36774
rect 10888 36038 10916 37402
rect 10980 37346 11008 39200
rect 10980 37330 11100 37346
rect 10980 37324 11112 37330
rect 10980 37318 11060 37324
rect 11060 37266 11112 37272
rect 12072 37324 12124 37330
rect 12072 37266 12124 37272
rect 11520 37256 11572 37262
rect 11520 37198 11572 37204
rect 11060 36848 11112 36854
rect 11060 36790 11112 36796
rect 10968 36576 11020 36582
rect 10968 36518 11020 36524
rect 10980 36310 11008 36518
rect 10968 36304 11020 36310
rect 10968 36246 11020 36252
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 10876 36032 10928 36038
rect 10876 35974 10928 35980
rect 10784 35556 10836 35562
rect 10784 35498 10836 35504
rect 10796 35154 10824 35498
rect 10980 35442 11008 36110
rect 10888 35414 11008 35442
rect 10784 35148 10836 35154
rect 10784 35090 10836 35096
rect 10704 35006 10824 35034
rect 10796 34950 10824 35006
rect 10784 34944 10836 34950
rect 10784 34886 10836 34892
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 10244 33318 10272 34342
rect 10416 33856 10468 33862
rect 10416 33798 10468 33804
rect 10428 33522 10456 33798
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10232 33312 10284 33318
rect 10232 33254 10284 33260
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10244 28082 10272 33254
rect 10324 32972 10376 32978
rect 10324 32914 10376 32920
rect 10336 31754 10364 32914
rect 10336 31726 10456 31754
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 10336 29170 10364 29514
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 9968 27934 10088 27962
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9404 26444 9456 26450
rect 9404 26386 9456 26392
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9416 25906 9444 26182
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9784 18698 9812 25638
rect 9968 25294 9996 27934
rect 10048 27872 10100 27878
rect 10048 27814 10100 27820
rect 10060 27674 10088 27814
rect 10048 27668 10100 27674
rect 10048 27610 10100 27616
rect 10048 26920 10100 26926
rect 10046 26888 10048 26897
rect 10100 26888 10102 26897
rect 10046 26823 10102 26832
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9876 16114 9904 24822
rect 9968 24818 9996 25230
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 10428 23730 10456 31726
rect 10598 27024 10654 27033
rect 10598 26959 10654 26968
rect 10612 26926 10640 26959
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10796 24818 10824 34886
rect 10888 33114 10916 35414
rect 10968 35284 11020 35290
rect 10968 35226 11020 35232
rect 10980 34746 11008 35226
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 11072 34202 11100 36790
rect 11532 36786 11560 37198
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 11532 36242 11560 36722
rect 12084 36310 12112 37266
rect 12912 37126 12940 39200
rect 14844 37262 14872 39200
rect 16776 37466 16804 39200
rect 18064 37466 18092 39200
rect 16764 37460 16816 37466
rect 16764 37402 16816 37408
rect 18052 37460 18104 37466
rect 18052 37402 18104 37408
rect 16776 37262 16804 37402
rect 18064 37262 18092 37402
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 12992 37256 13044 37262
rect 12992 37198 13044 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 16764 37256 16816 37262
rect 16764 37198 16816 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 12072 36304 12124 36310
rect 12072 36246 12124 36252
rect 11520 36236 11572 36242
rect 11520 36178 11572 36184
rect 12820 36106 12848 37062
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 12808 36100 12860 36106
rect 12808 36042 12860 36048
rect 11150 35456 11206 35465
rect 11150 35391 11206 35400
rect 11164 34746 11192 35391
rect 11152 34740 11204 34746
rect 11152 34682 11204 34688
rect 11336 34740 11388 34746
rect 11336 34682 11388 34688
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 11072 32910 11100 34138
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 11164 31414 11192 33798
rect 11152 31408 11204 31414
rect 11152 31350 11204 31356
rect 10876 29028 10928 29034
rect 10876 28970 10928 28976
rect 10888 27402 10916 28970
rect 11348 28762 11376 34682
rect 11336 28756 11388 28762
rect 11336 28698 11388 28704
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10980 27402 11008 27814
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10888 24410 10916 27338
rect 11256 26858 11284 27542
rect 11348 27402 11376 28698
rect 11336 27396 11388 27402
rect 11336 27338 11388 27344
rect 11244 26852 11296 26858
rect 11244 26794 11296 26800
rect 11256 26466 11284 26794
rect 11164 26438 11284 26466
rect 11164 25294 11192 26438
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10980 24818 11008 25094
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 11256 23254 11284 26318
rect 11348 25974 11376 27338
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11532 25498 11560 26250
rect 11612 25764 11664 25770
rect 11612 25706 11664 25712
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11624 25430 11652 25706
rect 11612 25424 11664 25430
rect 11612 25366 11664 25372
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11440 24886 11468 25162
rect 11428 24880 11480 24886
rect 11428 24822 11480 24828
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11348 22778 11376 24006
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11716 22094 11744 36042
rect 12348 35692 12400 35698
rect 12348 35634 12400 35640
rect 11980 34672 12032 34678
rect 11980 34614 12032 34620
rect 11796 33924 11848 33930
rect 11796 33866 11848 33872
rect 11808 33114 11836 33866
rect 11992 33658 12020 34614
rect 12360 34542 12388 35634
rect 12348 34536 12400 34542
rect 12348 34478 12400 34484
rect 12360 33930 12388 34478
rect 12440 34468 12492 34474
rect 12440 34410 12492 34416
rect 12348 33924 12400 33930
rect 12348 33866 12400 33872
rect 12360 33658 12388 33866
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 12348 33652 12400 33658
rect 12348 33594 12400 33600
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11992 33386 12020 33458
rect 11980 33380 12032 33386
rect 11980 33322 12032 33328
rect 11796 33108 11848 33114
rect 11796 33050 11848 33056
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 11980 30796 12032 30802
rect 11980 30738 12032 30744
rect 11992 29102 12020 30738
rect 12268 30258 12296 31826
rect 12452 30802 12480 34410
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12440 30796 12492 30802
rect 12440 30738 12492 30744
rect 12348 30660 12400 30666
rect 12348 30602 12400 30608
rect 12360 30394 12388 30602
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12268 29646 12296 30194
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 12084 28762 12112 29174
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11900 28150 11928 28494
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 12452 28098 12480 30738
rect 12544 29850 12572 32710
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12544 28694 12572 29786
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12636 28626 12664 29038
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12452 28070 12572 28098
rect 12440 27940 12492 27946
rect 12440 27882 12492 27888
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11992 24818 12020 26522
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11716 22066 12020 22094
rect 11992 20874 12020 22066
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 20534 11744 20742
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9416 15706 9444 15914
rect 9876 15706 9904 16050
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10520 2854 10548 15846
rect 10888 15706 10916 16118
rect 12268 16114 12296 26862
rect 12360 24206 12388 27066
rect 12452 26790 12480 27882
rect 12544 27538 12572 28070
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12636 26466 12664 28562
rect 12820 28558 12848 29106
rect 12912 28558 12940 31758
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12912 28082 12940 28494
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12544 26450 12664 26466
rect 12544 26444 12676 26450
rect 12544 26438 12624 26444
rect 12544 25430 12572 26438
rect 12624 26386 12676 26392
rect 12728 26314 12756 27270
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12636 25974 12664 26250
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12532 25424 12584 25430
rect 12532 25366 12584 25372
rect 12728 25226 12756 25638
rect 12820 25430 12848 27338
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12912 25702 12940 25842
rect 12900 25696 12952 25702
rect 12900 25638 12952 25644
rect 12808 25424 12860 25430
rect 12808 25366 12860 25372
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12820 24750 12848 25366
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12716 24676 12768 24682
rect 12716 24618 12768 24624
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23866 12388 24142
rect 12728 24070 12756 24618
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12820 23526 12848 24074
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 12912 16182 12940 23122
rect 13004 16998 13032 37198
rect 15200 37188 15252 37194
rect 15200 37130 15252 37136
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 14936 36786 14964 37062
rect 15212 36786 15240 37130
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 13096 30326 13124 36722
rect 13544 36712 13596 36718
rect 13544 36654 13596 36660
rect 13176 36576 13228 36582
rect 13176 36518 13228 36524
rect 13188 36310 13216 36518
rect 13176 36304 13228 36310
rect 13176 36246 13228 36252
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13464 35290 13492 35430
rect 13452 35284 13504 35290
rect 13452 35226 13504 35232
rect 13464 34746 13492 35226
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13556 33998 13584 36654
rect 14096 36576 14148 36582
rect 14096 36518 14148 36524
rect 14108 36378 14136 36518
rect 14096 36372 14148 36378
rect 14096 36314 14148 36320
rect 14004 36304 14056 36310
rect 14004 36246 14056 36252
rect 14016 35894 14044 36246
rect 14016 35866 14136 35894
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13832 33386 13860 34478
rect 14004 34128 14056 34134
rect 14004 34070 14056 34076
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13820 33380 13872 33386
rect 13820 33322 13872 33328
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13188 30938 13216 32370
rect 13176 30932 13228 30938
rect 13176 30874 13228 30880
rect 13084 30320 13136 30326
rect 13084 30262 13136 30268
rect 13544 30320 13596 30326
rect 13544 30262 13596 30268
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13268 28484 13320 28490
rect 13268 28426 13320 28432
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13188 27402 13216 28358
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 13176 27396 13228 27402
rect 13176 27338 13228 27344
rect 13096 26858 13124 27338
rect 13084 26852 13136 26858
rect 13084 26794 13136 26800
rect 13096 25362 13124 26794
rect 13280 25498 13308 28426
rect 13372 28082 13400 29446
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13360 27532 13412 27538
rect 13360 27474 13412 27480
rect 13372 27062 13400 27474
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 13464 26314 13492 29990
rect 13556 29306 13584 30262
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13832 28234 13860 29582
rect 13648 28206 13860 28234
rect 13648 28150 13676 28206
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13556 26897 13584 26930
rect 13542 26888 13598 26897
rect 13542 26823 13598 26832
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13096 24138 13124 24346
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13188 23322 13216 24074
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 13740 16114 13768 28018
rect 13832 27130 13860 28086
rect 13820 27124 13872 27130
rect 13820 27066 13872 27072
rect 13924 25294 13952 33458
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13820 24948 13872 24954
rect 13820 24890 13872 24896
rect 13832 24682 13860 24890
rect 13924 24818 13952 25230
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13924 22778 13952 24754
rect 14016 23118 14044 34070
rect 14108 26874 14136 35866
rect 14464 35760 14516 35766
rect 14462 35728 14464 35737
rect 14516 35728 14518 35737
rect 14462 35663 14518 35672
rect 14372 35556 14424 35562
rect 14372 35498 14424 35504
rect 14188 33856 14240 33862
rect 14188 33798 14240 33804
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14200 33590 14228 33798
rect 14188 33584 14240 33590
rect 14188 33526 14240 33532
rect 14292 33454 14320 33798
rect 14280 33448 14332 33454
rect 14280 33390 14332 33396
rect 14384 30190 14412 35498
rect 14740 34060 14792 34066
rect 14740 34002 14792 34008
rect 14556 33856 14608 33862
rect 14556 33798 14608 33804
rect 14464 32496 14516 32502
rect 14464 32438 14516 32444
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14292 29238 14320 29446
rect 14384 29322 14412 30126
rect 14476 29646 14504 32438
rect 14568 30802 14596 33798
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14660 30666 14688 31078
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14752 30190 14780 34002
rect 14936 33998 14964 36722
rect 16028 36644 16080 36650
rect 16028 36586 16080 36592
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15936 36576 15988 36582
rect 15936 36518 15988 36524
rect 15304 36242 15332 36518
rect 15948 36378 15976 36518
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15292 36236 15344 36242
rect 15292 36178 15344 36184
rect 15948 35834 15976 36314
rect 15936 35828 15988 35834
rect 15936 35770 15988 35776
rect 15948 35290 15976 35770
rect 15936 35284 15988 35290
rect 15936 35226 15988 35232
rect 15016 35012 15068 35018
rect 15016 34954 15068 34960
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14832 33924 14884 33930
rect 14832 33866 14884 33872
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14384 29294 14504 29322
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 14200 27878 14228 29038
rect 14384 28762 14412 29174
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14476 28642 14504 29294
rect 14752 29034 14780 30126
rect 14844 29510 14872 33866
rect 14924 33380 14976 33386
rect 14924 33322 14976 33328
rect 14832 29504 14884 29510
rect 14832 29446 14884 29452
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14384 28614 14504 28642
rect 14740 28620 14792 28626
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14292 27402 14320 27950
rect 14384 27606 14412 28614
rect 14740 28562 14792 28568
rect 14464 28484 14516 28490
rect 14464 28426 14516 28432
rect 14476 28218 14504 28426
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14384 27470 14412 27542
rect 14372 27464 14424 27470
rect 14424 27424 14504 27452
rect 14372 27406 14424 27412
rect 14280 27396 14332 27402
rect 14280 27338 14332 27344
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14200 27033 14228 27066
rect 14186 27024 14242 27033
rect 14186 26959 14242 26968
rect 14108 26846 14412 26874
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14200 23866 14228 24142
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14200 23186 14228 23666
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 14016 22506 14044 23054
rect 14292 22710 14320 24686
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 14016 22094 14044 22442
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14292 22098 14320 22374
rect 13924 22066 14044 22094
rect 14280 22092 14332 22098
rect 13924 21146 13952 22066
rect 14280 22034 14332 22040
rect 14384 21690 14412 26846
rect 14476 25906 14504 27424
rect 14568 27062 14596 27882
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14660 24886 14688 27610
rect 14752 27606 14780 28562
rect 14740 27600 14792 27606
rect 14740 27542 14792 27548
rect 14752 26518 14780 27542
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14568 24410 14596 24686
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14476 24070 14504 24142
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14568 23322 14596 24346
rect 14844 23746 14872 28698
rect 14936 25294 14964 33322
rect 15028 32502 15056 34954
rect 15108 34944 15160 34950
rect 15108 34886 15160 34892
rect 15016 32496 15068 32502
rect 15016 32438 15068 32444
rect 15120 31414 15148 34886
rect 16040 32502 16068 36586
rect 16304 35624 16356 35630
rect 16304 35566 16356 35572
rect 16028 32496 16080 32502
rect 16028 32438 16080 32444
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15304 29714 15332 30602
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15212 26926 15240 28970
rect 15396 28626 15424 31214
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15488 29102 15516 30534
rect 15580 29238 15608 32302
rect 15936 32292 15988 32298
rect 15936 32234 15988 32240
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 15764 30326 15792 31758
rect 15752 30320 15804 30326
rect 15752 30262 15804 30268
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15488 28014 15516 29038
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15764 28150 15792 28358
rect 15948 28150 15976 32234
rect 16040 31278 16068 32438
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 16040 28558 16068 30874
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 16132 29850 16160 30262
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 16132 29102 16160 29650
rect 16120 29096 16172 29102
rect 16120 29038 16172 29044
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15200 26920 15252 26926
rect 15200 26862 15252 26868
rect 15396 26450 15424 27882
rect 16040 27674 16068 28494
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15856 27418 15884 27474
rect 15856 27402 15976 27418
rect 15660 27396 15712 27402
rect 15856 27396 15988 27402
rect 15856 27390 15936 27396
rect 15660 27338 15712 27344
rect 15936 27338 15988 27344
rect 15672 27062 15700 27338
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15672 26314 15700 26386
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14936 24954 14964 25230
rect 15016 25152 15068 25158
rect 15016 25094 15068 25100
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14660 23730 14872 23746
rect 14648 23724 14872 23730
rect 14700 23718 14872 23724
rect 14648 23666 14700 23672
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14568 22234 14596 23258
rect 14936 23202 14964 24890
rect 15028 24206 15056 25094
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 24410 15148 24550
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15212 24274 15240 26250
rect 15764 25974 15792 27270
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 15856 25430 15884 26386
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 15844 25424 15896 25430
rect 15844 25366 15896 25372
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 15200 24268 15252 24274
rect 15200 24210 15252 24216
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15120 24154 15148 24210
rect 15120 24126 15240 24154
rect 14844 23186 14964 23202
rect 14832 23180 14964 23186
rect 14884 23174 14964 23180
rect 14832 23122 14884 23128
rect 15212 23050 15240 24126
rect 15580 23798 15608 25094
rect 15856 24750 15884 25366
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15304 23186 15332 23530
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14936 22094 14964 22646
rect 15212 22574 15240 22986
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 14936 22066 15056 22094
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 14476 20942 14504 21830
rect 14568 21690 14596 21966
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14936 21146 14964 21966
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14476 20262 14504 20878
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 8974 14412 9862
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10612 2650 10640 7754
rect 14476 7206 14504 20198
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12820 2922 12848 3470
rect 14568 3058 14596 19314
rect 15028 10810 15056 22066
rect 15396 21690 15424 22646
rect 15580 22094 15608 23598
rect 15488 22066 15608 22094
rect 15856 22094 15884 24686
rect 15948 22778 15976 25774
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 16040 25226 16068 25434
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 16132 23798 16160 29038
rect 16224 28422 16252 32166
rect 16316 30938 16344 35566
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16500 30734 16528 36722
rect 16856 36100 16908 36106
rect 16856 36042 16908 36048
rect 16868 30938 16896 36042
rect 16856 30932 16908 30938
rect 16856 30874 16908 30880
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16304 29232 16356 29238
rect 16304 29174 16356 29180
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16316 28082 16344 29174
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16316 26042 16344 28018
rect 16488 27532 16540 27538
rect 16488 27474 16540 27480
rect 16500 26450 16528 27474
rect 16684 27146 16712 29990
rect 16868 29646 16896 30874
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16776 27334 16804 28358
rect 16868 27538 16896 28562
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 16868 27402 16896 27474
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16684 27118 16804 27146
rect 16776 27062 16804 27118
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16304 26036 16356 26042
rect 16304 25978 16356 25984
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24274 16252 25094
rect 16500 24614 16528 26250
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 16592 24818 16620 25910
rect 16776 25838 16804 26998
rect 16868 25906 16896 27338
rect 16960 26586 16988 37062
rect 18156 35894 18184 37266
rect 19996 37126 20024 39200
rect 20352 37392 20404 37398
rect 20352 37334 20404 37340
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20088 36922 20116 37198
rect 20076 36916 20128 36922
rect 20076 36858 20128 36864
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 18156 35866 18368 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 18340 31754 18368 35866
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 18340 31726 18552 31754
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17960 31204 18012 31210
rect 17960 31146 18012 31152
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17420 29238 17448 29446
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17512 29102 17540 30126
rect 17972 30054 18000 31146
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17500 29096 17552 29102
rect 17500 29038 17552 29044
rect 17684 28688 17736 28694
rect 17684 28630 17736 28636
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17328 27674 17356 27814
rect 17316 27668 17368 27674
rect 17316 27610 17368 27616
rect 17132 27532 17184 27538
rect 17184 27492 17264 27520
rect 17132 27474 17184 27480
rect 17236 27130 17264 27492
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16684 24750 16712 25162
rect 16672 24744 16724 24750
rect 16672 24686 16724 24692
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16684 24206 16712 24686
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16028 23248 16080 23254
rect 16028 23190 16080 23196
rect 16040 23050 16068 23190
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 15856 22066 16160 22094
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15120 20602 15148 21558
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15120 20466 15148 20538
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15212 16454 15240 19654
rect 15304 19514 15332 20334
rect 15488 20058 15516 22066
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 20466 16068 20742
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 16132 16574 16160 22066
rect 16224 21418 16252 22578
rect 16212 21412 16264 21418
rect 16212 21354 16264 21360
rect 16132 16546 16344 16574
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 15978 15424 16390
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10470 15700 10610
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 3466 15700 10406
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 13004 2650 13032 2994
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2246
rect 5184 800 5212 2246
rect 7116 800 7144 2246
rect 8404 800 8432 2246
rect 10336 800 10364 2382
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 14200 800 14228 2926
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15488 800 15516 2450
rect 16040 2446 16068 3402
rect 16316 3126 16344 16546
rect 16408 15706 16436 23122
rect 16684 21962 16712 23462
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 21010 16620 21422
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 19922 16620 20198
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 10538 16436 15438
rect 16500 11354 16528 19790
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 10266 16436 10474
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16776 9654 16804 25774
rect 17052 23798 17080 26726
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16960 23186 16988 23598
rect 16948 23180 17000 23186
rect 16948 23122 17000 23128
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 17052 22506 17080 22986
rect 17040 22500 17092 22506
rect 17040 22442 17092 22448
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16960 21146 16988 22034
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16960 20602 16988 21082
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16960 20058 16988 20538
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17144 19378 17172 20402
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17144 18970 17172 19314
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 17144 2650 17172 11018
rect 17236 10810 17264 27066
rect 17328 26994 17356 27610
rect 17408 27124 17460 27130
rect 17408 27066 17460 27072
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17420 26858 17448 27066
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17512 26314 17540 26794
rect 17696 26586 17724 28630
rect 17880 28626 17908 29514
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17880 28014 17908 28562
rect 17972 28558 18000 29990
rect 18064 29238 18092 31214
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18432 29646 18460 29990
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 18052 29232 18104 29238
rect 18052 29174 18104 29180
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 17776 27600 17828 27606
rect 17828 27548 18000 27554
rect 17776 27542 18000 27548
rect 17788 27538 18000 27542
rect 17788 27532 18012 27538
rect 17788 27526 17960 27532
rect 17960 27474 18012 27480
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17500 26308 17552 26314
rect 17500 26250 17552 26256
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17684 26240 17736 26246
rect 17684 26182 17736 26188
rect 17696 25838 17724 26182
rect 17684 25832 17736 25838
rect 17684 25774 17736 25780
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17604 23798 17632 25706
rect 17788 24274 17816 26250
rect 17972 25974 18000 27474
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17788 23866 17816 24074
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17880 23730 17908 24686
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17696 22642 17724 22918
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 17696 21962 17724 22442
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17420 20602 17448 21422
rect 17696 21026 17724 21898
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17788 21146 17816 21422
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17696 20998 17816 21026
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17696 19446 17724 19654
rect 17684 19440 17736 19446
rect 17684 19382 17736 19388
rect 17696 14278 17724 19382
rect 17788 16574 17816 20998
rect 17880 20058 17908 23666
rect 17972 22710 18000 24346
rect 18064 23594 18092 29174
rect 18432 28558 18460 29582
rect 18524 28762 18552 31726
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 18616 29238 18644 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20364 29306 20392 37334
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20456 30870 20484 31282
rect 20444 30864 20496 30870
rect 20444 30806 20496 30812
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 18604 29232 18656 29238
rect 18604 29174 18656 29180
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 18512 28756 18564 28762
rect 18512 28698 18564 28704
rect 20088 28558 20116 29106
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 26926 18184 27950
rect 18524 27470 18552 28426
rect 18788 28416 18840 28422
rect 18788 28358 18840 28364
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18248 26926 18276 26998
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18156 25362 18184 26862
rect 18340 26042 18368 27270
rect 18432 27062 18460 27270
rect 18708 27062 18736 27950
rect 18800 27402 18828 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19352 27538 19380 27950
rect 20352 27940 20404 27946
rect 20352 27882 20404 27888
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18800 26450 18828 26726
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18156 24886 18184 25298
rect 18708 25226 18736 25638
rect 18696 25220 18748 25226
rect 18696 25162 18748 25168
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18616 24886 18644 25094
rect 19352 24886 19380 25162
rect 18144 24880 18196 24886
rect 18144 24822 18196 24828
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19352 23866 19380 24074
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 17972 21690 18000 22510
rect 18064 22234 18092 22986
rect 18340 22778 18368 23054
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18800 22574 18828 22918
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17972 19514 18000 21626
rect 18708 21554 18736 21830
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21010 18644 21286
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18708 20942 18736 21490
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17788 16546 17908 16574
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17420 9926 17448 10610
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 2990 17264 3334
rect 17420 3058 17448 9862
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17512 9382 17540 9522
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 3398 17540 9318
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17880 2990 17908 16546
rect 18800 10810 18828 20198
rect 19444 19666 19472 26386
rect 19628 26314 19656 26998
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19524 25968 19576 25974
rect 19524 25910 19576 25916
rect 19536 25498 19564 25910
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19996 25378 20024 27814
rect 20076 27396 20128 27402
rect 20076 27338 20128 27344
rect 20088 26586 20116 27338
rect 20364 27062 20392 27882
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20168 26920 20220 26926
rect 20168 26862 20220 26868
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 20088 25906 20116 26522
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25498 20116 25842
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19904 25350 20116 25378
rect 19904 25294 19932 25350
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24818 20024 25230
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 20088 24410 20116 25350
rect 20180 24818 20208 26862
rect 20352 26784 20404 26790
rect 20352 26726 20404 26732
rect 20364 26382 20392 26726
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20088 23730 20116 24006
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 20088 23526 20116 23666
rect 20364 23594 20392 26318
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19352 19638 19472 19666
rect 19352 16574 19380 19638
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 17882 19472 19314
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19352 16546 19472 16574
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17512 2446 17540 2790
rect 18340 2446 18368 10406
rect 19444 3194 19472 16546
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 2446 19748 2790
rect 19996 2514 20024 15846
rect 20088 11558 20116 23462
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17202 20392 17478
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20456 11218 20484 28358
rect 20916 26042 20944 37198
rect 21928 37074 21956 39200
rect 23860 37126 23888 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 22100 37120 22152 37126
rect 21928 37068 22100 37074
rect 21928 37062 22152 37068
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 21928 37046 22140 37062
rect 24596 35834 24624 37198
rect 25148 37126 25176 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 26884 37256 26936 37262
rect 26884 37198 26936 37204
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 25332 36582 25360 37198
rect 25320 36576 25372 36582
rect 25320 36518 25372 36524
rect 24584 35828 24636 35834
rect 24584 35770 24636 35776
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23124 32774 23152 35634
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 23124 31822 23152 32710
rect 23112 31816 23164 31822
rect 23112 31758 23164 31764
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 20904 26036 20956 26042
rect 20904 25978 20956 25984
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21468 25702 21496 25842
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21468 25294 21496 25638
rect 21652 25498 21680 25774
rect 23676 25770 23704 28018
rect 23664 25764 23716 25770
rect 23664 25706 23716 25712
rect 21640 25492 21692 25498
rect 21640 25434 21692 25440
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21468 24750 21496 25230
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23400 22778 23428 23054
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 25332 22098 25360 36518
rect 26896 24410 26924 37198
rect 27080 37126 27108 39200
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 27896 36712 27948 36718
rect 27896 36654 27948 36660
rect 27908 36310 27936 36654
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 28644 25498 28672 37198
rect 29012 37126 29040 39200
rect 30944 37262 30972 39200
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 32232 37126 32260 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 31036 36786 31064 37062
rect 32508 36922 32536 37198
rect 34440 37108 34468 39222
rect 36082 39200 36138 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 34520 37062 34572 37068
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 30024 29034 30052 29446
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 34808 27946 34836 37198
rect 36096 37126 36124 39200
rect 38028 37262 38056 39200
rect 38290 38176 38346 38185
rect 38290 38111 38346 38120
rect 38016 37256 38068 37262
rect 38016 37198 38068 37204
rect 37740 37188 37792 37194
rect 37740 37130 37792 37136
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 37556 35692 37608 35698
rect 37556 35634 37608 35640
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 37568 30938 37596 35634
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 36268 28484 36320 28490
rect 36268 28426 36320 28432
rect 34796 27940 34848 27946
rect 34796 27882 34848 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36280 25498 36308 28426
rect 37292 27130 37320 28970
rect 37280 27124 37332 27130
rect 37280 27066 37332 27072
rect 28632 25492 28684 25498
rect 28632 25434 28684 25440
rect 36268 25492 36320 25498
rect 36268 25434 36320 25440
rect 36280 25294 36308 25434
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 37648 25220 37700 25226
rect 37648 25162 37700 25168
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 26884 24404 26936 24410
rect 26884 24346 26936 24352
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27540 23526 27568 24006
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27540 22778 27568 23462
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 24584 19440 24636 19446
rect 24584 19382 24636 19388
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 23216 8022 23244 16050
rect 24596 8974 24624 19382
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 23756 3460 23808 3466
rect 23756 3402 23808 3408
rect 21376 3126 21404 3402
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 23768 3058 23796 3402
rect 24780 3194 24808 8774
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 23584 2582 23612 2790
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 27172 2446 27200 2790
rect 28552 2650 28580 24550
rect 29828 23520 29880 23526
rect 29828 23462 29880 23468
rect 28908 23044 28960 23050
rect 28908 22986 28960 22992
rect 28920 20602 28948 22986
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 17420 800 17448 2246
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2246
rect 22572 800 22600 2246
rect 24504 800 24532 2382
rect 29656 2378 29684 2790
rect 29840 2650 29868 23462
rect 31024 2984 31076 2990
rect 31024 2926 31076 2932
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 31036 2582 31064 2926
rect 32416 2650 32444 24686
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33692 15972 33744 15978
rect 33692 15914 33744 15920
rect 33704 2650 33732 15914
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 37660 4758 37688 25162
rect 37752 21894 37780 37130
rect 37924 36780 37976 36786
rect 37924 36722 37976 36728
rect 37832 34536 37884 34542
rect 37832 34478 37884 34484
rect 37844 29646 37872 34478
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37844 28558 37872 29582
rect 37832 28552 37884 28558
rect 37832 28494 37884 28500
rect 37936 26234 37964 36722
rect 38198 36136 38254 36145
rect 38198 36071 38200 36080
rect 38252 36071 38254 36080
rect 38200 36042 38252 36048
rect 38108 36032 38160 36038
rect 38108 35974 38160 35980
rect 38016 31136 38068 31142
rect 38016 31078 38068 31084
rect 38028 30734 38056 31078
rect 38120 30818 38148 35974
rect 38304 35834 38332 38111
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38292 35828 38344 35834
rect 38292 35770 38344 35776
rect 38292 34536 38344 34542
rect 38292 34478 38344 34484
rect 38304 34134 38332 34478
rect 38292 34128 38344 34134
rect 38290 34096 38292 34105
rect 38344 34096 38346 34105
rect 38290 34031 38346 34040
rect 38200 32836 38252 32842
rect 38200 32778 38252 32784
rect 38212 32745 38240 32778
rect 38198 32736 38254 32745
rect 38198 32671 38254 32680
rect 38120 30790 38332 30818
rect 38016 30728 38068 30734
rect 38016 30670 38068 30676
rect 38198 30696 38254 30705
rect 38108 30660 38160 30666
rect 38198 30631 38254 30640
rect 38108 30602 38160 30608
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38028 26994 38056 28358
rect 38016 26988 38068 26994
rect 38016 26930 38068 26936
rect 38120 26382 38148 30602
rect 38212 30598 38240 30631
rect 38200 30592 38252 30598
rect 38200 30534 38252 30540
rect 38200 29164 38252 29170
rect 38200 29106 38252 29112
rect 38212 28665 38240 29106
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38304 27878 38332 30790
rect 38292 27872 38344 27878
rect 38292 27814 38344 27820
rect 38200 26784 38252 26790
rect 38200 26726 38252 26732
rect 38212 26625 38240 26726
rect 38198 26616 38254 26625
rect 38198 26551 38254 26560
rect 38108 26376 38160 26382
rect 38108 26318 38160 26324
rect 38120 26234 38148 26318
rect 37844 26206 37964 26234
rect 38028 26206 38148 26234
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37844 20618 37872 26206
rect 38028 25362 38056 26206
rect 38016 25356 38068 25362
rect 38016 25298 38068 25304
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 38016 25152 38068 25158
rect 38016 25094 38068 25100
rect 38028 23730 38056 25094
rect 38304 24954 38332 25191
rect 38292 24948 38344 24954
rect 38292 24890 38344 24896
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 38200 23520 38252 23526
rect 38200 23462 38252 23468
rect 38212 23225 38240 23462
rect 38198 23216 38254 23225
rect 38198 23151 38254 23160
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 37924 21412 37976 21418
rect 37924 21354 37976 21360
rect 37752 20590 37872 20618
rect 37752 19174 37780 20590
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37740 19168 37792 19174
rect 37740 19110 37792 19116
rect 37844 13938 37872 20402
rect 37936 19310 37964 21354
rect 38028 20602 38056 21490
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38016 20596 38068 20602
rect 38016 20538 38068 20544
rect 38200 19372 38252 19378
rect 38200 19314 38252 19320
rect 37924 19304 37976 19310
rect 37924 19246 37976 19252
rect 38212 19145 38240 19314
rect 38198 19136 38254 19145
rect 38198 19071 38254 19080
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 37832 13932 37884 13938
rect 37832 13874 37884 13880
rect 38028 6390 38056 16934
rect 38304 16574 38332 21966
rect 38120 16546 38332 16574
rect 38120 8634 38148 16546
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38292 13864 38344 13870
rect 38292 13806 38344 13812
rect 38304 13705 38332 13806
rect 38290 13696 38346 13705
rect 38290 13631 38346 13640
rect 38304 13530 38332 13631
rect 38292 13524 38344 13530
rect 38292 13466 38344 13472
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38212 11665 38240 11698
rect 38198 11656 38254 11665
rect 38198 11591 38254 11600
rect 38200 10668 38252 10674
rect 38200 10610 38252 10616
rect 38212 10305 38240 10610
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38304 8265 38332 8434
rect 38290 8256 38346 8265
rect 38290 8191 38346 8200
rect 38016 6384 38068 6390
rect 38016 6326 38068 6332
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38212 6225 38240 6258
rect 38198 6216 38254 6225
rect 38198 6151 38254 6160
rect 37648 4752 37700 4758
rect 37648 4694 37700 4700
rect 38200 4548 38252 4554
rect 38200 4490 38252 4496
rect 38212 4185 38240 4490
rect 38198 4176 38254 4185
rect 38198 4111 38254 4120
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 34428 2916 34480 2922
rect 34428 2858 34480 2864
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 34440 2446 34468 2858
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36740 2650 36768 3470
rect 38660 3460 38712 3466
rect 38660 3402 38712 3408
rect 38108 2916 38160 2922
rect 38108 2858 38160 2864
rect 38120 2666 38148 2858
rect 38200 2848 38252 2854
rect 38198 2816 38200 2825
rect 38252 2816 38254 2825
rect 38198 2751 38254 2760
rect 36728 2644 36780 2650
rect 38120 2638 38240 2666
rect 36728 2586 36780 2592
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 26436 800 26464 2246
rect 28368 800 28396 2314
rect 29656 800 29684 2314
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 31772 1714 31800 2246
rect 31588 1686 31800 1714
rect 31588 800 31616 1686
rect 33520 800 33548 2314
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35452 800 35480 2246
rect 36740 800 36768 2382
rect 38212 2378 38240 2638
rect 38200 2372 38252 2378
rect 38200 2314 38252 2320
rect 38212 1465 38240 2314
rect 38198 1456 38254 1465
rect 38198 1391 38254 1400
rect 38672 800 38700 3402
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 5170 200 5226 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 14186 200 14242 800
rect 15474 200 15530 800
rect 17406 200 17462 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 38658 200 38714 800
<< via2 >>
rect 1582 36780 1638 36816
rect 1582 36760 1584 36780
rect 1584 36760 1636 36780
rect 1636 36760 1638 36780
rect 1950 36216 2006 36272
rect 1674 29280 1730 29336
rect 2042 33632 2098 33688
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 25880 1730 25936
rect 4066 38800 4122 38856
rect 2778 31320 2834 31376
rect 3422 31884 3478 31920
rect 3422 31864 3424 31884
rect 3424 31864 3476 31884
rect 3476 31864 3478 31884
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 5538 36660 5540 36680
rect 5540 36660 5592 36680
rect 5592 36660 5594 36680
rect 5538 36624 5594 36660
rect 5078 36100 5134 36136
rect 5078 36080 5080 36100
rect 5080 36080 5132 36100
rect 5132 36080 5134 36100
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4066 33360 4122 33416
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4618 31320 4674 31376
rect 3882 31184 3938 31240
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4894 32136 4950 32192
rect 5170 32136 5226 32192
rect 5354 31456 5410 31512
rect 6182 31456 6238 31512
rect 6182 31184 6238 31240
rect 6550 31884 6606 31920
rect 6550 31864 6552 31884
rect 6552 31864 6604 31884
rect 6604 31864 6606 31884
rect 7194 36624 7250 36680
rect 7930 36080 7986 36136
rect 8206 35400 8262 35456
rect 7562 33632 7618 33688
rect 7286 31320 7342 31376
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 9310 36216 9366 36272
rect 1674 23840 1730 23896
rect 1674 21836 1676 21856
rect 1676 21836 1728 21856
rect 1728 21836 1730 21856
rect 1674 21800 1730 21836
rect 1582 20476 1584 20496
rect 1584 20476 1636 20496
rect 1636 20476 1638 20496
rect 1582 20440 1638 20476
rect 1582 18420 1638 18456
rect 1582 18400 1584 18420
rect 1584 18400 1636 18420
rect 1636 18400 1638 18420
rect 1674 16396 1676 16416
rect 1676 16396 1728 16416
rect 1728 16396 1730 16416
rect 1674 16360 1730 16396
rect 1674 14340 1730 14376
rect 1674 14320 1676 14340
rect 1676 14320 1728 14340
rect 1728 14320 1730 14340
rect 1674 12960 1730 13016
rect 1674 10956 1676 10976
rect 1676 10956 1728 10976
rect 1728 10956 1730 10976
rect 1674 10920 1730 10956
rect 1674 8880 1730 8936
rect 1582 6840 1638 6896
rect 1674 5516 1676 5536
rect 1676 5516 1728 5536
rect 1728 5516 1730 5536
rect 1674 5480 1730 5516
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1674 3440 1730 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9954 35692 10010 35728
rect 9954 35672 9956 35692
rect 9956 35672 10008 35692
rect 10008 35672 10010 35692
rect 10046 26868 10048 26888
rect 10048 26868 10100 26888
rect 10100 26868 10102 26888
rect 10046 26832 10102 26868
rect 10598 26968 10654 27024
rect 11150 35400 11206 35456
rect 13542 26832 13598 26888
rect 14462 35708 14464 35728
rect 14464 35708 14516 35728
rect 14516 35708 14518 35728
rect 14462 35672 14518 35708
rect 14186 26968 14242 27024
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 1674 1400 1730 1456
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 38290 38120 38346 38176
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38198 36100 38254 36136
rect 38198 36080 38200 36100
rect 38200 36080 38252 36100
rect 38252 36080 38254 36100
rect 38290 34076 38292 34096
rect 38292 34076 38344 34096
rect 38344 34076 38346 34096
rect 38290 34040 38346 34076
rect 38198 32680 38254 32736
rect 38198 30640 38254 30696
rect 38198 28600 38254 28656
rect 38198 26560 38254 26616
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 38198 23160 38254 23216
rect 38198 21120 38254 21176
rect 38198 19080 38254 19136
rect 38198 15680 38254 15736
rect 38290 13640 38346 13696
rect 38198 11600 38254 11656
rect 38198 10240 38254 10296
rect 38290 8200 38346 8256
rect 38198 6160 38254 6216
rect 38198 4120 38254 4176
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 2796 38200 2816
rect 38200 2796 38252 2816
rect 38252 2796 38254 2816
rect 38198 2760 38254 2796
rect 38198 1400 38254 1456
<< metal3 >>
rect 200 38858 800 38888
rect 4061 38858 4127 38861
rect 200 38856 4127 38858
rect 200 38800 4066 38856
rect 4122 38800 4127 38856
rect 200 38798 4127 38800
rect 200 38768 800 38798
rect 4061 38795 4127 38798
rect 38285 38178 38351 38181
rect 39200 38178 39800 38208
rect 38285 38176 39800 38178
rect 38285 38120 38290 38176
rect 38346 38120 39800 38176
rect 38285 38118 39800 38120
rect 38285 38115 38351 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1577 36818 1643 36821
rect 200 36816 1643 36818
rect 200 36760 1582 36816
rect 1638 36760 1643 36816
rect 200 36758 1643 36760
rect 200 36728 800 36758
rect 1577 36755 1643 36758
rect 5533 36682 5599 36685
rect 7189 36682 7255 36685
rect 5533 36680 7255 36682
rect 5533 36624 5538 36680
rect 5594 36624 7194 36680
rect 7250 36624 7255 36680
rect 5533 36622 7255 36624
rect 5533 36619 5599 36622
rect 7189 36619 7255 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 1945 36274 2011 36277
rect 9305 36274 9371 36277
rect 1945 36272 9371 36274
rect 1945 36216 1950 36272
rect 2006 36216 9310 36272
rect 9366 36216 9371 36272
rect 1945 36214 9371 36216
rect 1945 36211 2011 36214
rect 9305 36211 9371 36214
rect 5073 36138 5139 36141
rect 7925 36138 7991 36141
rect 5073 36136 7991 36138
rect 5073 36080 5078 36136
rect 5134 36080 7930 36136
rect 7986 36080 7991 36136
rect 5073 36078 7991 36080
rect 5073 36075 5139 36078
rect 7925 36075 7991 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 9949 35730 10015 35733
rect 14457 35730 14523 35733
rect 9949 35728 14523 35730
rect 9949 35672 9954 35728
rect 10010 35672 14462 35728
rect 14518 35672 14523 35728
rect 9949 35670 14523 35672
rect 9949 35667 10015 35670
rect 14457 35667 14523 35670
rect 200 35368 800 35488
rect 8201 35458 8267 35461
rect 11145 35458 11211 35461
rect 8201 35456 11211 35458
rect 8201 35400 8206 35456
rect 8262 35400 11150 35456
rect 11206 35400 11211 35456
rect 8201 35398 11211 35400
rect 8201 35395 8267 35398
rect 11145 35395 11211 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 38285 34098 38351 34101
rect 39200 34098 39800 34128
rect 38285 34096 39800 34098
rect 38285 34040 38290 34096
rect 38346 34040 39800 34096
rect 38285 34038 39800 34040
rect 38285 34035 38351 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 2037 33690 2103 33693
rect 7557 33690 7623 33693
rect 2037 33688 7623 33690
rect 2037 33632 2042 33688
rect 2098 33632 7562 33688
rect 7618 33632 7623 33688
rect 2037 33630 7623 33632
rect 2037 33627 2103 33630
rect 7557 33627 7623 33630
rect 200 33418 800 33448
rect 4061 33418 4127 33421
rect 200 33416 4127 33418
rect 200 33360 4066 33416
rect 4122 33360 4127 33416
rect 200 33358 4127 33360
rect 200 33328 800 33358
rect 4061 33355 4127 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 38193 32738 38259 32741
rect 39200 32738 39800 32768
rect 38193 32736 39800 32738
rect 38193 32680 38198 32736
rect 38254 32680 39800 32736
rect 38193 32678 39800 32680
rect 38193 32675 38259 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4889 32194 4955 32197
rect 5165 32194 5231 32197
rect 4889 32192 5231 32194
rect 4889 32136 4894 32192
rect 4950 32136 5170 32192
rect 5226 32136 5231 32192
rect 4889 32134 5231 32136
rect 4889 32131 4955 32134
rect 5165 32131 5231 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 3417 31922 3483 31925
rect 6545 31922 6611 31925
rect 3417 31920 6611 31922
rect 3417 31864 3422 31920
rect 3478 31864 6550 31920
rect 6606 31864 6611 31920
rect 3417 31862 6611 31864
rect 3417 31859 3483 31862
rect 6545 31859 6611 31862
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 5349 31514 5415 31517
rect 6177 31514 6243 31517
rect 5349 31512 6243 31514
rect 5349 31456 5354 31512
rect 5410 31456 6182 31512
rect 6238 31456 6243 31512
rect 5349 31454 6243 31456
rect 5349 31451 5415 31454
rect 6177 31451 6243 31454
rect 200 31378 800 31408
rect 2773 31378 2839 31381
rect 200 31376 2839 31378
rect 200 31320 2778 31376
rect 2834 31320 2839 31376
rect 200 31318 2839 31320
rect 200 31288 800 31318
rect 2773 31315 2839 31318
rect 4613 31378 4679 31381
rect 7281 31378 7347 31381
rect 4613 31376 7347 31378
rect 4613 31320 4618 31376
rect 4674 31320 7286 31376
rect 7342 31320 7347 31376
rect 4613 31318 7347 31320
rect 4613 31315 4679 31318
rect 7281 31315 7347 31318
rect 3877 31242 3943 31245
rect 6177 31242 6243 31245
rect 3877 31240 6243 31242
rect 3877 31184 3882 31240
rect 3938 31184 6182 31240
rect 6238 31184 6243 31240
rect 3877 31182 6243 31184
rect 3877 31179 3943 31182
rect 6177 31179 6243 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 38193 30698 38259 30701
rect 39200 30698 39800 30728
rect 38193 30696 39800 30698
rect 38193 30640 38198 30696
rect 38254 30640 39800 30696
rect 38193 30638 39800 30640
rect 38193 30635 38259 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1669 29338 1735 29341
rect 200 29336 1735 29338
rect 200 29280 1674 29336
rect 1730 29280 1735 29336
rect 200 29278 1735 29280
rect 200 29248 800 29278
rect 1669 29275 1735 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1669 27978 1735 27981
rect 200 27976 1735 27978
rect 200 27920 1674 27976
rect 1730 27920 1735 27976
rect 200 27918 1735 27920
rect 200 27888 800 27918
rect 1669 27915 1735 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 10593 27026 10659 27029
rect 14181 27026 14247 27029
rect 10593 27024 14247 27026
rect 10593 26968 10598 27024
rect 10654 26968 14186 27024
rect 14242 26968 14247 27024
rect 10593 26966 14247 26968
rect 10593 26963 10659 26966
rect 14181 26963 14247 26966
rect 10041 26890 10107 26893
rect 13537 26890 13603 26893
rect 10041 26888 13603 26890
rect 10041 26832 10046 26888
rect 10102 26832 13542 26888
rect 13598 26832 13603 26888
rect 10041 26830 13603 26832
rect 10041 26827 10107 26830
rect 13537 26827 13603 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1669 25938 1735 25941
rect 200 25936 1735 25938
rect 200 25880 1674 25936
rect 1730 25880 1735 25936
rect 200 25878 1735 25880
rect 200 25848 800 25878
rect 1669 25875 1735 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1669 23898 1735 23901
rect 200 23896 1735 23898
rect 200 23840 1674 23896
rect 1730 23840 1735 23896
rect 200 23838 1735 23840
rect 200 23808 800 23838
rect 1669 23835 1735 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 38193 23218 38259 23221
rect 39200 23218 39800 23248
rect 38193 23216 39800 23218
rect 38193 23160 38198 23216
rect 38254 23160 39800 23216
rect 38193 23158 39800 23160
rect 38193 23155 38259 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 200 21858 800 21888
rect 1669 21858 1735 21861
rect 200 21856 1735 21858
rect 200 21800 1674 21856
rect 1730 21800 1735 21856
rect 200 21798 1735 21800
rect 200 21768 800 21798
rect 1669 21795 1735 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1577 20498 1643 20501
rect 200 20496 1643 20498
rect 200 20440 1582 20496
rect 1638 20440 1643 20496
rect 200 20438 1643 20440
rect 200 20408 800 20438
rect 1577 20435 1643 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1577 18458 1643 18461
rect 200 18456 1643 18458
rect 200 18400 1582 18456
rect 1638 18400 1643 18456
rect 200 18398 1643 18400
rect 200 18368 800 18398
rect 1577 18395 1643 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 39200 17688 39800 17808
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16418 800 16448
rect 1669 16418 1735 16421
rect 200 16416 1735 16418
rect 200 16360 1674 16416
rect 1730 16360 1735 16416
rect 200 16358 1735 16360
rect 200 16328 800 16358
rect 1669 16355 1735 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1669 14378 1735 14381
rect 200 14376 1735 14378
rect 200 14320 1674 14376
rect 1730 14320 1735 14376
rect 200 14318 1735 14320
rect 200 14288 800 14318
rect 1669 14315 1735 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 38285 13698 38351 13701
rect 39200 13698 39800 13728
rect 38285 13696 39800 13698
rect 38285 13640 38290 13696
rect 38346 13640 39800 13696
rect 38285 13638 39800 13640
rect 38285 13635 38351 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1669 13018 1735 13021
rect 200 13016 1735 13018
rect 200 12960 1674 13016
rect 1730 12960 1735 13016
rect 200 12958 1735 12960
rect 200 12928 800 12958
rect 1669 12955 1735 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 38193 11658 38259 11661
rect 39200 11658 39800 11688
rect 38193 11656 39800 11658
rect 38193 11600 38198 11656
rect 38254 11600 39800 11656
rect 38193 11598 39800 11600
rect 38193 11595 38259 11598
rect 39200 11568 39800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 200 10978 800 11008
rect 1669 10978 1735 10981
rect 200 10976 1735 10978
rect 200 10920 1674 10976
rect 1730 10920 1735 10976
rect 200 10918 1735 10920
rect 200 10888 800 10918
rect 1669 10915 1735 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 38285 8258 38351 8261
rect 39200 8258 39800 8288
rect 38285 8256 39800 8258
rect 38285 8200 38290 8256
rect 38346 8200 39800 8256
rect 38285 8198 39800 8200
rect 38285 8195 38351 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 38193 6218 38259 6221
rect 39200 6218 39800 6248
rect 38193 6216 39800 6218
rect 38193 6160 38198 6216
rect 38254 6160 39800 6216
rect 38193 6158 39800 6160
rect 38193 6155 38259 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 38193 1458 38259 1461
rect 38193 1456 39314 1458
rect 38193 1400 38198 1456
rect 38254 1400 39314 1456
rect 38193 1398 39314 1400
rect 38193 1395 38259 1398
rect 39254 1050 39314 1398
rect 39070 990 39314 1050
rect 39070 778 39130 990
rect 39200 778 39800 808
rect 39070 718 39800 778
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1667941163
transform 1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1667941163
transform -1 0 20700 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1667941163
transform -1 0 18860 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1667941163
transform -1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1667941163
transform 1 0 13616 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1667941163
transform 1 0 16836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1667941163
transform -1 0 21068 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1667941163
transform -1 0 13248 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1667941163
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1667941163
transform -1 0 12972 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1667941163
transform -1 0 12420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1667941163
transform -1 0 13800 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1667941163
transform -1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1667941163
transform -1 0 20792 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1667941163
transform 1 0 17848 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1667941163
transform -1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1667941163
transform -1 0 20792 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1667941163
transform 1 0 12420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1667941163
transform 1 0 13984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1667941163
transform 1 0 11776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1667941163
transform 1 0 9292 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1667941163
transform -1 0 9384 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 1667941163
transform 1 0 11316 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1667941163
transform -1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1667941163
transform -1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1667941163
transform -1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1667941163
transform 1 0 18308 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1667941163
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1667941163
transform -1 0 25668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1667941163
transform -1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1667941163
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1667941163
transform -1 0 20424 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1667941163
transform 1 0 9752 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1667941163
transform -1 0 9936 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1667941163
transform 1 0 10948 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1667941163
transform -1 0 9016 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1667941163
transform -1 0 5796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1667941163
transform 1 0 36248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1667941163
transform 1 0 20792 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1667941163
transform -1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1667941163
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1667941163
transform -1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1667941163
transform 1 0 12880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1667941163
transform -1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1667941163
transform -1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1667941163
transform 1 0 31648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1667941163
transform 1 0 8464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1667941163
transform 1 0 20240 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1667941163
transform -1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform 1 0 12972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform 1 0 5888 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform 1 0 6440 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform -1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 7176 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1667941163
transform 1 0 7728 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1667941163
transform -1 0 6900 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform 1 0 6992 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__CLK
timestamp 1667941163
transform 1 0 10488 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__CLK
timestamp 1667941163
transform 1 0 7912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__CLK
timestamp 1667941163
transform 1 0 7268 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__D
timestamp 1667941163
transform 1 0 8464 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__CLK
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__D
timestamp 1667941163
transform 1 0 13156 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__D
timestamp 1667941163
transform 1 0 7360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__CLK
timestamp 1667941163
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__D
timestamp 1667941163
transform 1 0 8372 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__CLK
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__CLK
timestamp 1667941163
transform 1 0 9384 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__CLK
timestamp 1667941163
transform -1 0 16652 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__D
timestamp 1667941163
transform -1 0 14260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__CLK
timestamp 1667941163
transform 1 0 12788 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__CLK
timestamp 1667941163
transform 1 0 6532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__CLK
timestamp 1667941163
transform 1 0 7912 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__CLK
timestamp 1667941163
transform -1 0 7360 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__CLK
timestamp 1667941163
transform -1 0 7912 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__D
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__CLK
timestamp 1667941163
transform 1 0 12972 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__D
timestamp 1667941163
transform -1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__CLK
timestamp 1667941163
transform 1 0 9292 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__D
timestamp 1667941163
transform 1 0 10212 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__CLK
timestamp 1667941163
transform 1 0 15824 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__CLK
timestamp 1667941163
transform 1 0 8464 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__CLK
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__CLK
timestamp 1667941163
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__D
timestamp 1667941163
transform 1 0 12328 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__CLK
timestamp 1667941163
transform 1 0 13340 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__D
timestamp 1667941163
transform 1 0 11040 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__CLK
timestamp 1667941163
transform 1 0 15272 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__D
timestamp 1667941163
transform 1 0 14260 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__CLK
timestamp 1667941163
transform 1 0 5060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__CLK
timestamp 1667941163
transform 1 0 9844 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__CLK
timestamp 1667941163
transform 1 0 12604 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__CLK
timestamp 1667941163
transform 1 0 15364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__D
timestamp 1667941163
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__CLK
timestamp 1667941163
transform 1 0 13616 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__D
timestamp 1667941163
transform 1 0 14996 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__CLK
timestamp 1667941163
transform 1 0 15548 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__D
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__CLK
timestamp 1667941163
transform 1 0 13064 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__CLK
timestamp 1667941163
transform 1 0 11500 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__CLK
timestamp 1667941163
transform 1 0 8464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__CLK
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__CLK
timestamp 1667941163
transform 1 0 7820 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__CLK
timestamp 1667941163
transform 1 0 7268 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__CLK
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform -1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform -1 0 20240 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1667941163
transform 1 0 21344 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1667941163
transform 1 0 2576 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform -1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1667941163
transform -1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1667941163
transform -1 0 24472 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1667941163
transform -1 0 27508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1667941163
transform -1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1667941163
transform 1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1667941163
transform -1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1667941163
transform -1 0 21252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1667941163
transform -1 0 27968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1667941163
transform -1 0 2668 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1667941163
transform -1 0 10120 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1667941163
transform 1 0 23736 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1667941163
transform -1 0 20608 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 10948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1667941163
transform -1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform 1 0 20608 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 25392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1667941163
transform 1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform -1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform -1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1667941163
transform -1 0 21344 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform -1 0 10672 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform -1 0 17020 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 14904 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 37628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 37628 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 37720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 37628 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 1748 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 13892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 37628 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 37628 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 37628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 37628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 37628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 14628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 12236 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 37628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 37628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 15732 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output47_A
timestamp 1667941163
transform 1 0 37444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1667941163
transform -1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1667941163
transform -1 0 14444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output69_A
timestamp 1667941163
transform -1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1667941163
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1667941163
transform -1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1667941163
transform 1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1667941163
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 1667941163
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1667941163
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1667941163
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1667941163
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_231
timestamp 1667941163
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_239
timestamp 1667941163
transform 1 0 23092 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_327
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1667941163
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_386
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_397
timestamp 1667941163
transform 1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1667941163
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_43
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_130
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1667941163
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1667941163
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_160
timestamp 1667941163
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1667941163
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_186
timestamp 1667941163
transform 1 0 18216 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_194
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1667941163
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_255
timestamp 1667941163
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_267
timestamp 1667941163
transform 1 0 25668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_292
timestamp 1667941163
transform 1 0 27968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1667941163
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_308
timestamp 1667941163
transform 1 0 29440 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_311
timestamp 1667941163
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_323
timestamp 1667941163
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1667941163
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_397
timestamp 1667941163
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_397
timestamp 1667941163
transform 1 0 37628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_241
timestamp 1667941163
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1667941163
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_398
timestamp 1667941163
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_288
timestamp 1667941163
transform 1 0 27600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1667941163
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1667941163
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_192
timestamp 1667941163
transform 1 0 18768 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_204
timestamp 1667941163
transform 1 0 19872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1667941163
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1667941163
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_179
timestamp 1667941163
transform 1 0 17572 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1667941163
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1667941163
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1667941163
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1667941163
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_194
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1667941163
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1667941163
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_397
timestamp 1667941163
transform 1 0 37628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_169
timestamp 1667941163
transform 1 0 16652 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1667941163
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1667941163
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1667941163
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1667941163
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1667941163
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_98
timestamp 1667941163
transform 1 0 10120 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_104
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_119
timestamp 1667941163
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_161
timestamp 1667941163
transform 1 0 15916 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_171
timestamp 1667941163
transform 1 0 16836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_183
timestamp 1667941163
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_100
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1667941163
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1667941163
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_127
timestamp 1667941163
transform 1 0 12788 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_139
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_201
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_212
timestamp 1667941163
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_397
timestamp 1667941163
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1667941163
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1667941163
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_154
timestamp 1667941163
transform 1 0 15272 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_211
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1667941163
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_7
timestamp 1667941163
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1667941163
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1667941163
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_56
timestamp 1667941163
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1667941163
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_174
timestamp 1667941163
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1667941163
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_177
timestamp 1667941163
transform 1 0 17388 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_191
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_203
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_397
timestamp 1667941163
transform 1 0 37628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_160
timestamp 1667941163
transform 1 0 15824 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1667941163
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1667941163
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_7
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_19
timestamp 1667941163
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_145
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_148
timestamp 1667941163
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1667941163
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_187
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_199
timestamp 1667941163
transform 1 0 19412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1667941163
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_313
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_402
timestamp 1667941163
transform 1 0 38088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1667941163
transform 1 0 38456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1667941163
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_152
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1667941163
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_183
timestamp 1667941163
transform 1 0 17940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_133
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1667941163
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_157
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1667941163
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_192
timestamp 1667941163
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_198
timestamp 1667941163
transform 1 0 19320 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_210
timestamp 1667941163
transform 1 0 20424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1667941163
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_155
timestamp 1667941163
transform 1 0 15364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1667941163
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1667941163
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_177
timestamp 1667941163
transform 1 0 17388 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_194
timestamp 1667941163
transform 1 0 18952 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_206
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1667941163
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_250
timestamp 1667941163
transform 1 0 24104 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_262
timestamp 1667941163
transform 1 0 25208 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1667941163
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_12
timestamp 1667941163
transform 1 0 2208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1667941163
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1667941163
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1667941163
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1667941163
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1667941163
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_157
timestamp 1667941163
transform 1 0 15548 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1667941163
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_187
timestamp 1667941163
transform 1 0 18308 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_207
timestamp 1667941163
transform 1 0 20148 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_219
timestamp 1667941163
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_231
timestamp 1667941163
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_117
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1667941163
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1667941163
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_144
timestamp 1667941163
transform 1 0 14352 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 1667941163
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1667941163
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_207
timestamp 1667941163
transform 1 0 20148 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_45
timestamp 1667941163
transform 1 0 5244 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_51
timestamp 1667941163
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_63
timestamp 1667941163
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 1667941163
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1667941163
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_125
timestamp 1667941163
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_151
timestamp 1667941163
transform 1 0 14996 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_159
timestamp 1667941163
transform 1 0 15732 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_169
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1667941163
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_188
timestamp 1667941163
transform 1 0 18400 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_208
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_220
timestamp 1667941163
transform 1 0 21344 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_232
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1667941163
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_281
timestamp 1667941163
transform 1 0 26956 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_287
timestamp 1667941163
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1667941163
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1667941163
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_17
timestamp 1667941163
transform 1 0 2668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_29
timestamp 1667941163
transform 1 0 3772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_41
timestamp 1667941163
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_72
timestamp 1667941163
transform 1 0 7728 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_84
timestamp 1667941163
transform 1 0 8832 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_92
timestamp 1667941163
transform 1 0 9568 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_96
timestamp 1667941163
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1667941163
transform 1 0 10580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_119
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1667941163
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_158
timestamp 1667941163
transform 1 0 15640 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1667941163
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_210
timestamp 1667941163
transform 1 0 20424 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_401
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1667941163
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1667941163
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1667941163
transform 1 0 12144 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_148
timestamp 1667941163
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1667941163
transform 1 0 15364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_172
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1667941163
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_214
timestamp 1667941163
transform 1 0 20792 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_225
timestamp 1667941163
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_231
timestamp 1667941163
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1667941163
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_300
timestamp 1667941163
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 1667941163
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_384
timestamp 1667941163
transform 1 0 36432 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_391
timestamp 1667941163
transform 1 0 37076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_90
timestamp 1667941163
transform 1 0 9384 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_96
timestamp 1667941163
transform 1 0 9936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_103
timestamp 1667941163
transform 1 0 10580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1667941163
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1667941163
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_139
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1667941163
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1667941163
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_195
timestamp 1667941163
transform 1 0 19044 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_209
timestamp 1667941163
transform 1 0 20332 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_216
timestamp 1667941163
transform 1 0 20976 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1667941163
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1667941163
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_98
timestamp 1667941163
transform 1 0 10120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1667941163
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_150
timestamp 1667941163
transform 1 0 14904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_171
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1667941163
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1667941163
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_216
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1667941163
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1667941163
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_92
timestamp 1667941163
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1667941163
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_104
timestamp 1667941163
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_122
timestamp 1667941163
transform 1 0 12328 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_129
timestamp 1667941163
transform 1 0 12972 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1667941163
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1667941163
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1667941163
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1667941163
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1667941163
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1667941163
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_7
timestamp 1667941163
transform 1 0 1748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1667941163
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_96
timestamp 1667941163
transform 1 0 9936 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_104
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_114
timestamp 1667941163
transform 1 0 11592 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1667941163
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_163
timestamp 1667941163
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_176
timestamp 1667941163
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1667941163
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_220
timestamp 1667941163
transform 1 0 21344 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_232
timestamp 1667941163
transform 1 0 22448 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_17
timestamp 1667941163
transform 1 0 2668 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_21
timestamp 1667941163
transform 1 0 3036 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_28
timestamp 1667941163
transform 1 0 3680 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_34
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_46
timestamp 1667941163
transform 1 0 5336 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_63
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_75
timestamp 1667941163
transform 1 0 8004 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_87
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_95
timestamp 1667941163
transform 1 0 9844 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_99
timestamp 1667941163
transform 1 0 10212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1667941163
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1667941163
transform 1 0 11960 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_122
timestamp 1667941163
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_126
timestamp 1667941163
transform 1 0 12696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_133
timestamp 1667941163
transform 1 0 13340 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_153
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1667941163
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_187
timestamp 1667941163
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1667941163
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_201
timestamp 1667941163
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1667941163
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1667941163
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1667941163
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_248
timestamp 1667941163
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_254
timestamp 1667941163
transform 1 0 24472 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_266
timestamp 1667941163
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_14
timestamp 1667941163
transform 1 0 2392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1667941163
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_34
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_38
timestamp 1667941163
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_42
timestamp 1667941163
transform 1 0 4968 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_50
timestamp 1667941163
transform 1 0 5704 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_54
timestamp 1667941163
transform 1 0 6072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_61
timestamp 1667941163
transform 1 0 6716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_68
timestamp 1667941163
transform 1 0 7360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_74
timestamp 1667941163
transform 1 0 7912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_96
timestamp 1667941163
transform 1 0 9936 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_105
timestamp 1667941163
transform 1 0 10764 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_113
timestamp 1667941163
transform 1 0 11500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_120
timestamp 1667941163
transform 1 0 12144 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_156
timestamp 1667941163
transform 1 0 15456 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_163
timestamp 1667941163
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1667941163
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_203
timestamp 1667941163
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1667941163
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_214
timestamp 1667941163
transform 1 0 20792 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_226
timestamp 1667941163
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_238
timestamp 1667941163
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1667941163
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_397
timestamp 1667941163
transform 1 0 37628 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_402
timestamp 1667941163
transform 1 0 38088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1667941163
transform 1 0 38456 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1667941163
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1667941163
transform 1 0 2392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1667941163
transform 1 0 3680 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_35
timestamp 1667941163
transform 1 0 4324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_42
timestamp 1667941163
transform 1 0 4968 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_50
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_62
timestamp 1667941163
transform 1 0 6808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_68
timestamp 1667941163
transform 1 0 7360 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_85
timestamp 1667941163
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_97
timestamp 1667941163
transform 1 0 10028 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_103
timestamp 1667941163
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_126
timestamp 1667941163
transform 1 0 12696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_150
timestamp 1667941163
transform 1 0 14904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1667941163
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1667941163
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_204
timestamp 1667941163
transform 1 0 19872 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_210
timestamp 1667941163
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_397
timestamp 1667941163
transform 1 0 37628 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_19
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_36
timestamp 1667941163
transform 1 0 4416 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_43
timestamp 1667941163
transform 1 0 5060 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1667941163
transform 1 0 6072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_60
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_66
timestamp 1667941163
transform 1 0 7176 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1667941163
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1667941163
transform 1 0 12604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_131
timestamp 1667941163
transform 1 0 13156 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1667941163
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_149
timestamp 1667941163
transform 1 0 14812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_166
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1667941163
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_176
timestamp 1667941163
transform 1 0 17296 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_187
timestamp 1667941163
transform 1 0 18308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1667941163
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_316
timestamp 1667941163
transform 1 0 30176 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1667941163
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_340
timestamp 1667941163
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_352
timestamp 1667941163
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_16
timestamp 1667941163
transform 1 0 2576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_23
timestamp 1667941163
transform 1 0 3220 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_34
timestamp 1667941163
transform 1 0 4232 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_38
timestamp 1667941163
transform 1 0 4600 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_42
timestamp 1667941163
transform 1 0 4968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1667941163
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_62
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_68
timestamp 1667941163
transform 1 0 7360 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_74
timestamp 1667941163
transform 1 0 7912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_86
timestamp 1667941163
transform 1 0 9016 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1667941163
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1667941163
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_151
timestamp 1667941163
transform 1 0 14996 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_173
timestamp 1667941163
transform 1 0 17020 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_184
timestamp 1667941163
transform 1 0 18032 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_190
timestamp 1667941163
transform 1 0 18584 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1667941163
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1667941163
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_10
timestamp 1667941163
transform 1 0 2024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_17
timestamp 1667941163
transform 1 0 2668 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1667941163
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_34
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_48
timestamp 1667941163
transform 1 0 5520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_72
timestamp 1667941163
transform 1 0 7728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1667941163
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_102
timestamp 1667941163
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_106
timestamp 1667941163
transform 1 0 10856 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1667941163
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_129
timestamp 1667941163
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1667941163
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_154
timestamp 1667941163
transform 1 0 15272 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_161
timestamp 1667941163
transform 1 0 15916 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_167
timestamp 1667941163
transform 1 0 16468 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_173
timestamp 1667941163
transform 1 0 17020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1667941163
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1667941163
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_393
timestamp 1667941163
transform 1 0 37260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_397
timestamp 1667941163
transform 1 0 37628 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_79
timestamp 1667941163
transform 1 0 8372 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_86
timestamp 1667941163
transform 1 0 9016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1667941163
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_98
timestamp 1667941163
transform 1 0 10120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_142
timestamp 1667941163
transform 1 0 14168 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_209
timestamp 1667941163
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1667941163
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1667941163
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_58
timestamp 1667941163
transform 1 0 6440 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_89
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_95
timestamp 1667941163
transform 1 0 9844 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_107
timestamp 1667941163
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_119
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_185
timestamp 1667941163
transform 1 0 18124 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp 1667941163
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_201
timestamp 1667941163
transform 1 0 19596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_213
timestamp 1667941163
transform 1 0 20700 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_225
timestamp 1667941163
transform 1 0 21804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_237
timestamp 1667941163
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1667941163
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_19
timestamp 1667941163
transform 1 0 2852 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_43
timestamp 1667941163
transform 1 0 5060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1667941163
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_63
timestamp 1667941163
transform 1 0 6900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_85
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1667941163
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_97
timestamp 1667941163
transform 1 0 10028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_103
timestamp 1667941163
transform 1 0 10580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_121
timestamp 1667941163
transform 1 0 12236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1667941163
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_134
timestamp 1667941163
transform 1 0 13432 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_146
timestamp 1667941163
transform 1 0 14536 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_162
timestamp 1667941163
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_35
timestamp 1667941163
transform 1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_39
timestamp 1667941163
transform 1 0 4692 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_63
timestamp 1667941163
transform 1 0 6900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_69
timestamp 1667941163
transform 1 0 7452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_75
timestamp 1667941163
transform 1 0 8004 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1667941163
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_89
timestamp 1667941163
transform 1 0 9292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_95
timestamp 1667941163
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1667941163
transform 1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_107
timestamp 1667941163
transform 1 0 10948 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_114
timestamp 1667941163
transform 1 0 11592 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_126
timestamp 1667941163
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_397
timestamp 1667941163
transform 1 0 37628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_32
timestamp 1667941163
transform 1 0 4048 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_42
timestamp 1667941163
transform 1 0 4968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1667941163
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_80
timestamp 1667941163
transform 1 0 8464 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_104
timestamp 1667941163
transform 1 0 10672 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1667941163
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1667941163
transform 1 0 11960 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_124
timestamp 1667941163
transform 1 0 12512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_136
timestamp 1667941163
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1667941163
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_37
timestamp 1667941163
transform 1 0 4508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_64
timestamp 1667941163
transform 1 0 6992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_70
timestamp 1667941163
transform 1 0 7544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_76
timestamp 1667941163
transform 1 0 8096 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_107
timestamp 1667941163
transform 1 0 10948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_113
timestamp 1667941163
transform 1 0 11500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_123
timestamp 1667941163
transform 1 0 12420 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_130
timestamp 1667941163
transform 1 0 13064 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_134
timestamp 1667941163
transform 1 0 13432 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_146
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1667941163
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_32
timestamp 1667941163
transform 1 0 4048 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1667941163
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1667941163
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_104
timestamp 1667941163
transform 1 0 10672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1667941163
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_131
timestamp 1667941163
transform 1 0 13156 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_143
timestamp 1667941163
transform 1 0 14260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_155
timestamp 1667941163
transform 1 0 15364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1667941163
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_35
timestamp 1667941163
transform 1 0 4324 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_43
timestamp 1667941163
transform 1 0 5060 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_67
timestamp 1667941163
transform 1 0 7268 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_73
timestamp 1667941163
transform 1 0 7820 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_76
timestamp 1667941163
transform 1 0 8096 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_107
timestamp 1667941163
transform 1 0 10948 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_115
timestamp 1667941163
transform 1 0 11684 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1667941163
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_126
timestamp 1667941163
transform 1 0 12696 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_132
timestamp 1667941163
transform 1 0 13248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_145
timestamp 1667941163
transform 1 0 14444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_157
timestamp 1667941163
transform 1 0 15548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_169
timestamp 1667941163
transform 1 0 16652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_181
timestamp 1667941163
transform 1 0 17756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1667941163
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_32
timestamp 1667941163
transform 1 0 4048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_40
timestamp 1667941163
transform 1 0 4784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_47
timestamp 1667941163
transform 1 0 5428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_61
timestamp 1667941163
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_65
timestamp 1667941163
transform 1 0 7084 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_87
timestamp 1667941163
transform 1 0 9108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_98
timestamp 1667941163
transform 1 0 10120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_104
timestamp 1667941163
transform 1 0 10672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1667941163
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_119
timestamp 1667941163
transform 1 0 12052 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_123
timestamp 1667941163
transform 1 0 12420 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_129
timestamp 1667941163
transform 1 0 12972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1667941163
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_147
timestamp 1667941163
transform 1 0 14628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_153
timestamp 1667941163
transform 1 0 15180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1667941163
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1667941163
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_248
timestamp 1667941163
transform 1 0 23920 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_260
timestamp 1667941163
transform 1 0 25024 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_272
timestamp 1667941163
transform 1 0 26128 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_35
timestamp 1667941163
transform 1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_39
timestamp 1667941163
transform 1 0 4692 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_63
timestamp 1667941163
transform 1 0 6900 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1667941163
transform 1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_76
timestamp 1667941163
transform 1 0 8096 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_107
timestamp 1667941163
transform 1 0 10948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_115
timestamp 1667941163
transform 1 0 11684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_127
timestamp 1667941163
transform 1 0 12788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_145
timestamp 1667941163
transform 1 0 14444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_151
timestamp 1667941163
transform 1 0 14996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1667941163
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_163
timestamp 1667941163
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_169
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_181
timestamp 1667941163
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1667941163
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_42
timestamp 1667941163
transform 1 0 4968 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_82
timestamp 1667941163
transform 1 0 8648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_106
timestamp 1667941163
transform 1 0 10856 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_135
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_150
timestamp 1667941163
transform 1 0 14904 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_156
timestamp 1667941163
transform 1 0 15456 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1667941163
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_186
timestamp 1667941163
transform 1 0 18216 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_198
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_210
timestamp 1667941163
transform 1 0 20424 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1667941163
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_295
timestamp 1667941163
transform 1 0 28244 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_307
timestamp 1667941163
transform 1 0 29348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_319
timestamp 1667941163
transform 1 0 30452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_331
timestamp 1667941163
transform 1 0 31556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_343
timestamp 1667941163
transform 1 0 32660 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_355
timestamp 1667941163
transform 1 0 33764 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_367
timestamp 1667941163
transform 1 0 34868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_379
timestamp 1667941163
transform 1 0 35972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_397
timestamp 1667941163
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1667941163
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1667941163
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_163
timestamp 1667941163
transform 1 0 16100 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_243
timestamp 1667941163
transform 1 0 23460 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_355
timestamp 1667941163
transform 1 0 33764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_359
timestamp 1667941163
transform 1 0 34132 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_397
timestamp 1667941163
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _115_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1667941163
transform 1 0 12880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1667941163
transform 1 0 12420 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1667941163
transform -1 0 12512 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1667941163
transform 1 0 13524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1667941163
transform 1 0 11316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1667941163
transform 1 0 13064 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1667941163
transform 1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1667941163
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1667941163
transform 1 0 12420 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1667941163
transform 1 0 18032 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1667941163
transform -1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130_
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1667941163
transform -1 0 19688 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132_
timestamp 1667941163
transform 1 0 11776 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp 1667941163
transform 1 0 14628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1667941163
transform -1 0 16100 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1667941163
transform 1 0 10120 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1667941163
transform -1 0 19964 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1667941163
transform 1 0 13800 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1667941163
transform 1 0 12696 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1667941163
transform 1 0 10488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1667941163
transform -1 0 20424 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1667941163
transform 1 0 14444 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1667941163
transform 1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1667941163
transform -1 0 10212 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1667941163
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1667941163
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1667941163
transform 1 0 13156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1667941163
transform -1 0 20332 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1667941163
transform -1 0 18308 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1667941163
transform 1 0 12512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1667941163
transform -1 0 19688 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1667941163
transform -1 0 19688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1667941163
transform 1 0 17480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1667941163
transform 1 0 12788 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1667941163
transform -1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1667941163
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1667941163
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1667941163
transform 1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1667941163
transform 1 0 8096 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1667941163
transform 1 0 13432 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1667941163
transform -1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1667941163
transform 1 0 8740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1667941163
transform 1 0 11868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1667941163
transform -1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1667941163
transform -1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1667941163
transform 1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1667941163
transform 1 0 10580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1667941163
transform -1 0 16192 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1667941163
transform -1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1667941163
transform -1 0 18768 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1667941163
transform -1 0 17940 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1667941163
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1667941163
transform -1 0 18308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1667941163
transform -1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1667941163
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1667941163
transform -1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1667941163
transform 1 0 10304 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1667941163
transform -1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1667941163
transform -1 0 30268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1667941163
transform -1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1667941163
transform -1 0 19872 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1667941163
transform -1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1667941163
transform -1 0 18676 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _196_
timestamp 1667941163
transform -1 0 12052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1667941163
transform 1 0 11500 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1667941163
transform 1 0 12052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1667941163
transform 1 0 4968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1667941163
transform 1 0 36800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _201_
timestamp 1667941163
transform -1 0 20424 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1667941163
transform 1 0 14904 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1667941163
transform -1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1667941163
transform -1 0 15916 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1667941163
transform -1 0 29256 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _206_
timestamp 1667941163
transform -1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1667941163
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1667941163
transform -1 0 19320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1667941163
transform -1 0 15088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _210_
timestamp 1667941163
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1667941163
transform -1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1667941163
transform -1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _213_
timestamp 1667941163
transform -1 0 19596 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _214_
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform 1 0 9844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform -1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform -1 0 21804 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 12420 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform -1 0 30176 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _224_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 28244 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _225_
timestamp 1667941163
transform -1 0 4968 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform 1 0 4692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform 1 0 5336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform 1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform 1 0 4784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform -1 0 3496 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 4232 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform -1 0 4324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 4140 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _236_
timestamp 1667941163
transform -1 0 5888 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform 1 0 2760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 5704 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 3680 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 4232 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform 1 0 5244 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _247_
timestamp 1667941163
transform -1 0 4508 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform 1 0 2392 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 2760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 1932 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 3312 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform 1 0 2944 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 2300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 2116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform 1 0 2116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform 1 0 2576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 5796 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 6808 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 6440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 6072 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _264_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10856 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1667941163
transform -1 0 10948 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _267_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 6900 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _268_
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _269_
timestamp 1667941163
transform -1 0 6900 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1667941163
transform -1 0 3496 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1667941163
transform -1 0 3496 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _273_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 9108 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _274_
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _275_
timestamp 1667941163
transform -1 0 8464 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1667941163
transform -1 0 8372 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1667941163
transform 1 0 5888 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _279_
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _280_
timestamp 1667941163
transform -1 0 4048 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _281_
timestamp 1667941163
transform -1 0 4968 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1667941163
transform -1 0 10672 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1667941163
transform 1 0 8832 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1667941163
transform 1 0 1656 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _285_
timestamp 1667941163
transform -1 0 8648 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _286_
timestamp 1667941163
transform -1 0 8648 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _287_
timestamp 1667941163
transform -1 0 5060 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp 1667941163
transform -1 0 3496 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp 1667941163
transform -1 0 10948 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _290_
timestamp 1667941163
transform 1 0 1656 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _291_
timestamp 1667941163
transform -1 0 4048 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _292_
timestamp 1667941163
transform -1 0 6072 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _293_
timestamp 1667941163
transform -1 0 7268 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1667941163
transform 1 0 4600 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _297_
timestamp 1667941163
transform -1 0 8924 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp 1667941163
transform 1 0 6808 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _299_
timestamp 1667941163
transform 1 0 1656 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1667941163
transform -1 0 28704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1667941163
transform -1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _310_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1667941163
transform 1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1667941163
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1667941163
transform -1 0 38088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1667941163
transform 1 0 14076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1667941163
transform 1 0 5152 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1667941163
transform -1 0 23920 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1667941163
transform -1 0 26956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1667941163
transform 1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1667941163
transform 1 0 14352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1667941163
transform -1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1667941163
transform 1 0 15548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1667941163
transform -1 0 20700 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1667941163
transform -1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _325_
timestamp 1667941163
transform 1 0 15824 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _326_
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _327_
timestamp 1667941163
transform -1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1667941163
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1667941163
transform 1 0 37720 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1667941163
transform -1 0 23368 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp 1667941163
transform -1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1667941163
transform -1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _333_
timestamp 1667941163
transform -1 0 10764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1667941163
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1667941163
transform -1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1667941163
transform -1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1667941163
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1667941163
transform -1 0 37628 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1667941163
transform -1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1667941163
transform 1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1667941163
transform 1 0 4416 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _344_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18308 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _345_
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _346_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17388 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _347_
timestamp 1667941163
transform -1 0 18676 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _348__86 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _348_
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _349_
timestamp 1667941163
transform 1 0 16376 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _350_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _351_
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _352_
timestamp 1667941163
transform 1 0 12972 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _353_
timestamp 1667941163
transform -1 0 20148 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _354_
timestamp 1667941163
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _355_
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _356_
timestamp 1667941163
transform -1 0 9936 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _357_
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _357__87
timestamp 1667941163
transform -1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _358_
timestamp 1667941163
transform 1 0 7176 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _359_
timestamp 1667941163
transform 1 0 8096 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _360_
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _361_
timestamp 1667941163
transform -1 0 13432 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _362_
timestamp 1667941163
transform 1 0 12512 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _363_
timestamp 1667941163
transform 1 0 11316 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _364_
timestamp 1667941163
transform -1 0 9936 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _365_
timestamp 1667941163
transform -1 0 14996 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _366_
timestamp 1667941163
transform 1 0 11868 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _367_
timestamp 1667941163
transform 1 0 10764 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _368_
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _369_
timestamp 1667941163
transform -1 0 18308 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _370_
timestamp 1667941163
transform -1 0 18952 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _371__88
timestamp 1667941163
transform 1 0 18676 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _371_
timestamp 1667941163
transform -1 0 18676 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _372_
timestamp 1667941163
transform 1 0 15364 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _373_
timestamp 1667941163
transform 1 0 14444 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _374_
timestamp 1667941163
transform -1 0 17848 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _375_
timestamp 1667941163
transform -1 0 16100 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _376_
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _377_
timestamp 1667941163
transform -1 0 18952 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _378_
timestamp 1667941163
transform 1 0 15272 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _379_
timestamp 1667941163
transform -1 0 17296 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _380_
timestamp 1667941163
transform 1 0 14444 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _381_
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _382_
timestamp 1667941163
transform -1 0 18400 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _383__89
timestamp 1667941163
transform -1 0 14904 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _383_
timestamp 1667941163
transform 1 0 15824 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _384_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _385_
timestamp 1667941163
transform 1 0 14628 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _386_
timestamp 1667941163
transform 1 0 14352 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _387_
timestamp 1667941163
transform -1 0 17664 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _388_
timestamp 1667941163
transform 1 0 15272 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _389_
timestamp 1667941163
transform -1 0 18952 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _390_
timestamp 1667941163
transform -1 0 15548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _391_
timestamp 1667941163
transform -1 0 17756 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _392_
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _393_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _394_
timestamp 1667941163
transform -1 0 19044 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _395__90
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _395_
timestamp 1667941163
transform -1 0 18492 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _396_
timestamp 1667941163
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _397_
timestamp 1667941163
transform -1 0 17664 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _398_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _399_
timestamp 1667941163
transform -1 0 18860 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _400_
timestamp 1667941163
transform -1 0 16376 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _401_
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _402_
timestamp 1667941163
transform -1 0 16100 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _403_
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _404_
timestamp 1667941163
transform 1 0 11592 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _405__91
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _405_
timestamp 1667941163
transform 1 0 13984 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _406_
timestamp 1667941163
transform 1 0 14076 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _407_
timestamp 1667941163
transform -1 0 16376 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _408_
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _409_
timestamp 1667941163
transform -1 0 14812 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _410_
timestamp 1667941163
transform 1 0 11776 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _411_
timestamp 1667941163
transform -1 0 16008 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _412_
timestamp 1667941163
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform 1 0 5704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform -1 0 38364 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform -1 0 38364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 38364 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform -1 0 38364 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform -1 0 38364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 36708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform -1 0 16376 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform -1 0 38364 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform -1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform -1 0 38364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 4416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform -1 0 38364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform -1 0 38364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform -1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 7820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 1932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform -1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform -1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 4324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform -1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 13340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 36524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform -1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 10120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 1932 0 1 13056
box -38 -48 406 592
<< labels >>
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal2 s 15474 200 15530 800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal3 s 200 16328 800 16448 0 FreeSans 480 0 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 78 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 79 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 80 nsew signal tristate
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 pReset
port 81 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 prog_clk
port 82 nsew signal input
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 83 nsew signal tristate
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 84 nsew signal tristate
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 85 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 86 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 86 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 86 nsew signal bidirectional
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 vssd1
port 87 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 87 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 8878 36142 8878 36142 0 _000_
rlabel metal2 9844 34986 9844 34986 0 _001_
rlabel metal1 7176 30090 7176 30090 0 _002_
rlabel metal2 5474 33218 5474 33218 0 _003_
rlabel metal1 5198 30906 5198 30906 0 _004_
rlabel metal3 5060 32164 5060 32164 0 _005_
rlabel metal2 2714 32402 2714 32402 0 _006_
rlabel metal1 3956 30294 3956 30294 0 _007_
rlabel metal2 2530 33218 2530 33218 0 _008_
rlabel metal1 5198 29750 5198 29750 0 _009_
rlabel metal2 4922 32300 4922 32300 0 _010_
rlabel metal1 5290 29070 5290 29070 0 _011_
rlabel metal1 4140 31654 4140 31654 0 _012_
rlabel metal1 5375 30634 5375 30634 0 _013_
rlabel metal1 5612 32198 5612 32198 0 _014_
rlabel metal1 3450 34510 3450 34510 0 _015_
rlabel metal2 2622 31076 2622 31076 0 _016_
rlabel metal2 5796 34170 5796 34170 0 _017_
rlabel metal1 1978 30906 1978 30906 0 _018_
rlabel metal2 9016 33558 9016 33558 0 _019_
rlabel metal1 2760 30906 2760 30906 0 _020_
rlabel metal1 4140 28730 4140 28730 0 _021_
rlabel metal2 7176 36924 7176 36924 0 _022_
rlabel metal1 3213 32470 3213 32470 0 _023_
rlabel metal1 2744 32810 2744 32810 0 _024_
rlabel metal2 8740 33388 8740 33388 0 _025_
rlabel metal2 3174 30549 3174 30549 0 _026_
rlabel metal2 2254 32198 2254 32198 0 _027_
rlabel metal1 2300 29274 2300 29274 0 _028_
rlabel metal2 3358 32300 3358 32300 0 _029_
rlabel metal2 13110 33524 13110 33524 0 _030_
rlabel metal1 7912 28662 7912 28662 0 _031_
rlabel metal1 6171 31790 6171 31790 0 _032_
rlabel metal1 7307 32470 7307 32470 0 _033_
rlabel metal1 6440 28730 6440 28730 0 _034_
rlabel metal1 4784 29682 4784 29682 0 _035_
rlabel metal1 16560 36210 16560 36210 0 _036_
rlabel metal1 4462 30226 4462 30226 0 _037_
rlabel metal1 3818 28526 3818 28526 0 _038_
rlabel metal1 2116 30226 2116 30226 0 _039_
rlabel metal1 18124 22202 18124 22202 0 _040_
rlabel metal1 15226 22678 15226 22678 0 _041_
rlabel metal2 17802 21284 17802 21284 0 _042_
rlabel metal1 18446 19312 18446 19312 0 _043_
rlabel metal1 17710 20978 17710 20978 0 _044_
rlabel metal2 16606 20060 16606 20060 0 _045_
rlabel metal2 12834 23800 12834 23800 0 _046_
rlabel metal2 15134 24480 15134 24480 0 _047_
rlabel metal1 13386 23290 13386 23290 0 _048_
rlabel metal1 17802 22746 17802 22746 0 _049_
rlabel metal1 15962 20434 15962 20434 0 _050_
rlabel metal1 14950 23086 14950 23086 0 _051_
rlabel metal2 9706 29784 9706 29784 0 _052_
rlabel metal1 13294 25976 13294 25976 0 _053_
rlabel metal1 7498 24922 7498 24922 0 _054_
rlabel metal2 8326 29886 8326 29886 0 _055_
rlabel metal2 12742 25432 12742 25432 0 _056_
rlabel metal1 12650 24820 12650 24820 0 _057_
rlabel metal2 12742 26792 12742 26792 0 _058_
rlabel metal1 11546 25160 11546 25160 0 _059_
rlabel metal1 9660 27370 9660 27370 0 _060_
rlabel metal2 13570 29784 13570 29784 0 _061_
rlabel metal1 12052 28730 12052 28730 0 _062_
rlabel metal2 10994 27608 10994 27608 0 _063_
rlabel metal1 13892 33898 13892 33898 0 _064_
rlabel metal1 14306 32266 14306 32266 0 _065_
rlabel metal1 18676 24854 18676 24854 0 _066_
rlabel metal2 18446 27166 18446 27166 0 _067_
rlabel metal2 15594 24446 15594 24446 0 _068_
rlabel metal2 14674 30872 14674 30872 0 _069_
rlabel metal1 16422 24786 16422 24786 0 _070_
rlabel metal1 15870 27336 15870 27336 0 _071_
rlabel metal1 14766 32198 14766 32198 0 _072_
rlabel metal2 18722 25432 18722 25432 0 _073_
rlabel metal1 14030 28730 14030 28730 0 _074_
rlabel metal1 19274 26010 19274 26010 0 _075_
rlabel metal2 14674 26248 14674 26248 0 _076_
rlabel metal2 13294 26962 13294 26962 0 _077_
rlabel metal1 16330 23834 16330 23834 0 _078_
rlabel metal1 15904 24106 15904 24106 0 _079_
rlabel metal2 14490 24106 14490 24106 0 _080_
rlabel metal1 14582 22066 14582 22066 0 _081_
rlabel metal1 13340 27098 13340 27098 0 _082_
rlabel metal1 17158 24854 17158 24854 0 _083_
rlabel metal2 13478 28152 13478 28152 0 _084_
rlabel metal1 19090 26282 19090 26282 0 _085_
rlabel metal2 15318 23358 15318 23358 0 _086_
rlabel metal2 17526 26554 17526 26554 0 _087_
rlabel metal2 15042 33728 15042 33728 0 _088_
rlabel metal2 14490 28322 14490 28322 0 _089_
rlabel metal2 19550 25704 19550 25704 0 _090_
rlabel metal1 18538 27370 18538 27370 0 _091_
rlabel metal2 15778 28254 15778 28254 0 _092_
rlabel metal2 17434 29342 17434 29342 0 _093_
rlabel metal2 17066 25262 17066 25262 0 _094_
rlabel metal2 18630 29342 18630 29342 0 _095_
rlabel metal1 13846 34918 13846 34918 0 _096_
rlabel metal1 11178 25466 11178 25466 0 _097_
rlabel metal1 15824 25942 15824 25942 0 _098_
rlabel metal1 18262 23800 18262 23800 0 _099_
rlabel metal1 11638 33082 11638 33082 0 _100_
rlabel metal2 14214 33694 14214 33694 0 _101_
rlabel metal2 14306 29342 14306 29342 0 _102_
rlabel metal1 15410 29818 15410 29818 0 _103_
rlabel metal2 12374 30498 12374 30498 0 _104_
rlabel metal2 14582 27472 14582 27472 0 _105_
rlabel metal1 11914 33626 11914 33626 0 _106_
rlabel metal1 15732 27030 15732 27030 0 _107_
rlabel metal2 13202 27880 13202 27880 0 _108_
rlabel metal1 8464 2278 8464 2278 0 ccff_head
rlabel metal2 1702 26061 1702 26061 0 ccff_tail
rlabel metal1 2208 32402 2208 32402 0 chany_bottom_in[0]
rlabel metal1 17894 37434 17894 37434 0 chany_bottom_in[10]
rlabel metal2 5842 36958 5842 36958 0 chany_bottom_in[11]
rlabel metal2 38226 6239 38226 6239 0 chany_bottom_in[12]
rlabel metal2 38226 32759 38226 32759 0 chany_bottom_in[13]
rlabel metal2 38318 8347 38318 8347 0 chany_bottom_in[14]
rlabel metal1 28520 2346 28520 2346 0 chany_bottom_in[15]
rlabel via2 38226 36091 38226 36091 0 chany_bottom_in[16]
rlabel via2 1610 36771 1610 36771 0 chany_bottom_in[17]
rlabel metal1 14260 2958 14260 2958 0 chany_bottom_in[18]
rlabel metal2 38226 28883 38226 28883 0 chany_bottom_in[1]
rlabel metal2 38226 1887 38226 1887 0 chany_bottom_in[2]
rlabel via2 38318 25245 38318 25245 0 chany_bottom_in[3]
rlabel via2 1702 14331 1702 14331 0 chany_bottom_in[4]
rlabel metal1 38134 37230 38134 37230 0 chany_bottom_in[5]
rlabel metal2 38318 13583 38318 13583 0 chany_bottom_in[6]
rlabel metal2 16790 38328 16790 38328 0 chany_bottom_in[7]
rlabel metal1 36846 2414 36846 2414 0 chany_bottom_in[8]
rlabel metal1 33672 2346 33672 2346 0 chany_bottom_in[9]
rlabel metal2 35466 1520 35466 1520 0 chany_bottom_out[0]
rlabel metal1 25346 37094 25346 37094 0 chany_bottom_out[10]
rlabel metal2 38226 26673 38226 26673 0 chany_bottom_out[11]
rlabel metal2 19366 1520 19366 1520 0 chany_bottom_out[12]
rlabel metal3 1188 23868 1188 23868 0 chany_bottom_out[13]
rlabel metal2 38226 15793 38226 15793 0 chany_bottom_out[14]
rlabel metal1 22172 37094 22172 37094 0 chany_bottom_out[15]
rlabel metal3 1188 29308 1188 29308 0 chany_bottom_out[16]
rlabel metal1 29486 37094 29486 37094 0 chany_bottom_out[17]
rlabel metal3 1188 3468 1188 3468 0 chany_bottom_out[18]
rlabel metal2 38226 30617 38226 30617 0 chany_bottom_out[1]
rlabel metal3 1188 1428 1188 1428 0 chany_bottom_out[2]
rlabel metal1 20148 37094 20148 37094 0 chany_bottom_out[3]
rlabel metal3 1188 8908 1188 8908 0 chany_bottom_out[4]
rlabel metal3 1188 21828 1188 21828 0 chany_bottom_out[5]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[6]
rlabel metal1 34822 37094 34822 37094 0 chany_bottom_out[7]
rlabel metal2 690 37240 690 37240 0 chany_bottom_out[8]
rlabel metal2 2622 37784 2622 37784 0 chany_bottom_out[9]
rlabel metal1 15916 2482 15916 2482 0 chany_top_in[0]
rlabel metal3 1142 6868 1142 6868 0 chany_top_in[10]
rlabel via2 38318 34085 38318 34085 0 chany_top_in[11]
rlabel via2 1610 20485 1610 20485 0 chany_top_in[12]
rlabel metal1 3312 2278 3312 2278 0 chany_top_in[13]
rlabel metal1 10396 2414 10396 2414 0 chany_top_in[14]
rlabel metal2 31786 1989 31786 1989 0 chany_top_in[15]
rlabel metal2 38226 11679 38226 11679 0 chany_top_in[16]
rlabel metal2 38226 4335 38226 4335 0 chany_top_in[17]
rlabel metal1 24564 2414 24564 2414 0 chany_top_in[18]
rlabel metal1 4554 35768 4554 35768 0 chany_top_in[1]
rlabel metal1 38456 3434 38456 3434 0 chany_top_in[2]
rlabel metal1 11408 37298 11408 37298 0 chany_top_in[3]
rlabel metal2 38226 10455 38226 10455 0 chany_top_in[4]
rlabel metal2 38226 19227 38226 19227 0 chany_top_in[5]
rlabel metal1 29808 2346 29808 2346 0 chany_top_in[6]
rlabel via2 1610 18411 1610 18411 0 chany_top_in[7]
rlabel metal1 7912 36142 7912 36142 0 chany_top_in[8]
rlabel metal1 14996 37230 14996 37230 0 chany_top_in[9]
rlabel metal2 4094 33235 4094 33235 0 chany_top_out[0]
rlabel metal2 46 1656 46 1656 0 chany_top_out[10]
rlabel metal2 22586 1520 22586 1520 0 chany_top_out[11]
rlabel metal1 13018 37094 13018 37094 0 chany_top_out[12]
rlabel metal1 24334 37094 24334 37094 0 chany_top_out[13]
rlabel metal1 36202 37094 36202 37094 0 chany_top_out[14]
rlabel metal3 1188 27948 1188 27948 0 chany_top_out[15]
rlabel metal2 5198 1520 5198 1520 0 chany_top_out[16]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[17]
rlabel metal1 38778 36890 38778 36890 0 chany_top_out[18]
rlabel metal3 1188 5508 1188 5508 0 chany_top_out[1]
rlabel metal2 17434 1520 17434 1520 0 chany_top_out[2]
rlabel metal3 38786 38148 38786 38148 0 chany_top_out[3]
rlabel via2 38226 2805 38226 2805 0 chany_top_out[4]
rlabel metal3 1188 10948 1188 10948 0 chany_top_out[5]
rlabel metal2 38226 21233 38226 21233 0 chany_top_out[6]
rlabel metal2 7130 1520 7130 1520 0 chany_top_out[7]
rlabel metal2 12282 1520 12282 1520 0 chany_top_out[8]
rlabel via2 1702 16405 1702 16405 0 chany_top_out[9]
rlabel metal2 38226 23341 38226 23341 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal2 21298 1520 21298 1520 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal1 32338 37094 32338 37094 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal1 14122 21114 14122 21114 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal2 17158 19142 17158 19142 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 18124 20910 18124 20910 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal1 9200 36006 9200 36006 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal1 10856 34918 10856 34918 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal1 8418 33558 8418 33558 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal2 12834 28832 12834 28832 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal1 8832 34442 8832 34442 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal1 13271 34646 13271 34646 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal1 1610 37094 1610 37094 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal1 3542 34918 3542 34918 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal2 1978 31110 1978 31110 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal1 13018 28050 13018 28050 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal1 10442 31858 10442 31858 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 14214 29614 14214 29614 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal1 8832 33898 8832 33898 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal1 10994 34170 10994 34170 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal1 13524 36686 13524 36686 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal2 20102 26962 20102 26962 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal1 13754 34510 13754 34510 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 20148 27438 20148 27438 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal2 13202 31654 13202 31654 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal1 12834 33898 12834 33898 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal1 12558 32300 12558 32300 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal2 20378 24956 20378 24956 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal1 7682 36686 7682 36686 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal2 6578 35156 6578 35156 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal1 8326 33422 8326 33422 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 10442 33286 10442 33286 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal1 9430 34374 9430 34374 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 14168 35530 14168 35530 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal1 15686 35598 15686 35598 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 14398 36074 14398 36074 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal1 12466 35122 12466 35122 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal2 9154 36040 9154 36040 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal2 13110 24242 13110 24242 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal2 15042 16429 15042 16429 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 29532 20570 29532 20570 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal2 23414 22916 23414 22916 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 19596 17850 19596 17850 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 17526 20570 17526 20570 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal2 15318 19924 15318 19924 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal1 16468 19822 16468 19822 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal2 15226 23341 15226 23341 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18032 21658 18032 21658 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 16974 21590 16974 21590 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 24886 2992 24886 2992 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 13110 27098 13110 27098 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 11960 30770 11960 30770 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal2 11454 25024 11454 25024 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal2 12650 26112 12650 26112 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal1 17158 31790 17158 31790 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal1 5336 24378 5336 24378 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal1 13018 25398 13018 25398 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 12788 26418 12788 26418 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 13478 25772 13478 25772 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7682 18734 7682 18734 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 17204 27506 17204 27506 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal1 16882 9622 16882 9622 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal1 14766 27846 14766 27846 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal2 30038 29240 30038 29240 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal1 12512 30770 12512 30770 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15180 30158 15180 30158 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 12374 33762 12374 33762 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 25599 26282 25599 26282 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal1 15456 29070 15456 29070 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal1 15594 20026 15594 20026 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal1 14812 33830 14812 33830 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 19090 25194 19090 25194 0 mux_right_ipin_0.INVTX1_6_.out
rlabel metal1 19090 24718 19090 24718 0 mux_right_ipin_0.INVTX1_7_.out
rlabel metal2 16882 26690 16882 26690 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16100 29070 16100 29070 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18170 27438 18170 27438 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 36570 25262 36570 25262 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17756 20026 17756 20026 0 mux_right_ipin_1.INVTX1_2_.out
rlabel metal1 16284 15674 16284 15674 0 mux_right_ipin_1.INVTX1_3_.out
rlabel metal2 14214 24004 14214 24004 0 mux_right_ipin_1.INVTX1_4_.out
rlabel metal2 14950 21556 14950 21556 0 mux_right_ipin_1.INVTX1_5_.out
rlabel metal2 18814 26588 18814 26588 0 mux_right_ipin_1.INVTX1_6_.out
rlabel metal1 18814 24106 18814 24106 0 mux_right_ipin_1.INVTX1_7_.out
rlabel metal2 15410 27166 15410 27166 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14628 24378 14628 24378 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17802 25262 17802 25262 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 19182 3060 19182 3060 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19228 29070 19228 29070 0 mux_right_ipin_2.INVTX1_2_.out
rlabel metal1 16054 22746 16054 22746 0 mux_right_ipin_2.INVTX1_3_.out
rlabel metal1 10718 26282 10718 26282 0 mux_right_ipin_2.INVTX1_6_.out
rlabel metal2 21666 25636 21666 25636 0 mux_right_ipin_2.INVTX1_7_.out
rlabel metal2 18078 30226 18078 30226 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15272 32334 15272 32334 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17986 26724 17986 26724 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32062 36754 32062 36754 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 9154 2482 9154 2482 0 net1
rlabel metal1 2024 24786 2024 24786 0 net10
rlabel metal1 14904 19346 14904 19346 0 net11
rlabel metal2 37306 28050 37306 28050 0 net12
rlabel metal1 21574 2890 21574 2890 0 net13
rlabel metal2 38042 25775 38042 25775 0 net14
rlabel metal1 21160 19414 21160 19414 0 net15
rlabel metal1 29210 37366 29210 37366 0 net16
rlabel metal1 37950 13906 37950 13906 0 net17
rlabel metal1 9936 15674 9936 15674 0 net18
rlabel metal2 23782 3230 23782 3230 0 net19
rlabel metal2 2438 32096 2438 32096 0 net2
rlabel metal1 15180 19686 15180 19686 0 net20
rlabel metal2 21390 3264 21390 3264 0 net21
rlabel metal1 14536 20230 14536 20230 0 net22
rlabel metal2 37858 31518 37858 31518 0 net23
rlabel metal1 18538 20230 18538 20230 0 net24
rlabel metal1 4462 2482 4462 2482 0 net25
rlabel metal2 10626 5202 10626 5202 0 net26
rlabel metal2 32430 13668 32430 13668 0 net27
rlabel metal1 23161 11526 23161 11526 0 net28
rlabel metal1 37858 4726 37858 4726 0 net29
rlabel metal2 18170 36589 18170 36589 0 net3
rlabel metal1 24886 2550 24886 2550 0 net30
rlabel metal2 20470 31076 20470 31076 0 net31
rlabel metal2 17250 3162 17250 3162 0 net32
rlabel metal2 15226 36958 15226 36958 0 net33
rlabel metal1 16629 15334 16629 15334 0 net34
rlabel metal1 37996 19278 37996 19278 0 net35
rlabel metal1 23782 22610 23782 22610 0 net36
rlabel metal1 24012 28050 24012 28050 0 net37
rlabel metal1 5474 35666 5474 35666 0 net38
rlabel metal1 14628 36754 14628 36754 0 net39
rlabel metal1 20148 16082 20148 16082 0 net4
rlabel metal1 29624 36754 29624 36754 0 net40
rlabel metal1 1794 32742 1794 32742 0 net41
rlabel metal1 35006 2414 35006 2414 0 net42
rlabel metal1 18170 21964 18170 21964 0 net43
rlabel metal2 38042 27676 38042 27676 0 net44
rlabel metal1 18906 2414 18906 2414 0 net45
rlabel metal1 1932 23290 1932 23290 0 net46
rlabel metal2 23230 12036 23230 12036 0 net47
rlabel metal1 21482 37230 21482 37230 0 net48
rlabel metal1 1886 29002 1886 29002 0 net49
rlabel metal1 20700 17170 20700 17170 0 net5
rlabel metal1 29210 37230 29210 37230 0 net50
rlabel metal2 12834 3196 12834 3196 0 net51
rlabel metal2 38042 30906 38042 30906 0 net52
rlabel metal1 12926 2958 12926 2958 0 net53
rlabel metal1 18584 36890 18584 36890 0 net54
rlabel metal2 14398 9418 14398 9418 0 net55
rlabel metal1 14628 21658 14628 21658 0 net56
rlabel metal1 27048 37230 27048 37230 0 net57
rlabel metal1 34868 37230 34868 37230 0 net58
rlabel metal1 4508 35054 4508 35054 0 net59
rlabel metal1 19044 31790 19044 31790 0 net6
rlabel metal2 14122 36448 14122 36448 0 net60
rlabel metal1 4462 32878 4462 32878 0 net61
rlabel metal1 2714 2414 2714 2414 0 net62
rlabel metal1 21390 2482 21390 2482 0 net63
rlabel metal1 16652 16966 16652 16966 0 net64
rlabel metal1 23966 35802 23966 35802 0 net65
rlabel metal1 37122 37162 37122 37162 0 net66
rlabel metal1 12926 26758 12926 26758 0 net67
rlabel metal2 5566 2788 5566 2788 0 net68
rlabel metal1 2116 2414 2116 2414 0 net69
rlabel metal1 38134 21998 38134 21998 0 net7
rlabel metal2 37766 19873 37766 19873 0 net70
rlabel metal1 2116 5678 2116 5678 0 net71
rlabel metal2 17526 2618 17526 2618 0 net72
rlabel metal2 37582 33286 37582 33286 0 net73
rlabel metal1 37766 3026 37766 3026 0 net74
rlabel metal1 2162 11118 2162 11118 0 net75
rlabel metal2 38042 21046 38042 21046 0 net76
rlabel metal1 8602 15878 8602 15878 0 net77
rlabel metal2 23598 2686 23598 2686 0 net78
rlabel metal1 14490 16490 14490 16490 0 net79
rlabel metal2 28566 13600 28566 13600 0 net8
rlabel metal2 38042 24412 38042 24412 0 net80
rlabel metal1 20884 2414 20884 2414 0 net81
rlabel metal2 32522 37060 32522 37060 0 net82
rlabel metal1 11178 35666 11178 35666 0 net83
rlabel metal2 27186 2618 27186 2618 0 net84
rlabel metal1 4462 18598 4462 18598 0 net85
rlabel metal2 16606 21216 16606 21216 0 net86
rlabel metal1 12558 25806 12558 25806 0 net87
rlabel metal1 18630 27030 18630 27030 0 net88
rlabel metal1 15594 24242 15594 24242 0 net89
rlabel metal2 38318 29325 38318 29325 0 net9
rlabel metal1 18860 27506 18860 27506 0 net90
rlabel metal1 14214 33422 14214 33422 0 net91
rlabel metal1 31096 37230 31096 37230 0 pReset
rlabel metal1 1978 34442 1978 34442 0 prog_clk
rlabel metal1 9798 35530 9798 35530 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
rlabel metal2 26450 1520 26450 1520 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel metal3 1188 12988 1188 12988 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
