magic
tech sky130A
magscale 1 2
timestamp 1674175245
<< viali >>
rect 1777 37213 1811 37247
rect 2421 37213 2455 37247
rect 3065 37213 3099 37247
rect 4169 37213 4203 37247
rect 4629 37213 4663 37247
rect 6561 37213 6595 37247
rect 7849 37213 7883 37247
rect 9321 37213 9355 37247
rect 10425 37213 10459 37247
rect 12541 37213 12575 37247
rect 14289 37213 14323 37247
rect 15577 37213 15611 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22201 37213 22235 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 26065 37213 26099 37247
rect 27997 37213 28031 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 35081 37213 35115 37247
rect 36921 37213 36955 37247
rect 38025 37213 38059 37247
rect 1593 37077 1627 37111
rect 2237 37077 2271 37111
rect 2881 37077 2915 37111
rect 3985 37077 4019 37111
rect 4813 37077 4847 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9137 37077 9171 37111
rect 10609 37077 10643 37111
rect 12357 37077 12391 37111
rect 14473 37077 14507 37111
rect 15761 37077 15795 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 22017 37077 22051 37111
rect 22661 37077 22695 37111
rect 24777 37077 24811 37111
rect 25881 37077 25915 37111
rect 27813 37077 27847 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 34897 37077 34931 37111
rect 36737 37077 36771 37111
rect 38209 37077 38243 37111
rect 9137 36873 9171 36907
rect 1777 36737 1811 36771
rect 9321 36737 9355 36771
rect 37657 36737 37691 36771
rect 38301 36737 38335 36771
rect 1593 36533 1627 36567
rect 37473 36533 37507 36567
rect 38117 36533 38151 36567
rect 15761 36329 15795 36363
rect 15945 36125 15979 36159
rect 38301 36125 38335 36159
rect 38117 35989 38151 36023
rect 10701 35241 10735 35275
rect 10609 35037 10643 35071
rect 38025 35037 38059 35071
rect 38209 34901 38243 34935
rect 16865 34697 16899 34731
rect 22845 34697 22879 34731
rect 17049 34561 17083 34595
rect 23029 34561 23063 34595
rect 7297 34153 7331 34187
rect 13277 34153 13311 34187
rect 14289 34153 14323 34187
rect 7481 33949 7515 33983
rect 13461 33949 13495 33983
rect 14473 33949 14507 33983
rect 19441 33609 19475 33643
rect 1593 33473 1627 33507
rect 14197 33473 14231 33507
rect 19625 33473 19659 33507
rect 23397 33473 23431 33507
rect 24869 33473 24903 33507
rect 38025 33473 38059 33507
rect 1777 33337 1811 33371
rect 38209 33337 38243 33371
rect 14289 33269 14323 33303
rect 23489 33269 23523 33303
rect 24961 33269 24995 33303
rect 9781 33065 9815 33099
rect 9965 32861 9999 32895
rect 16865 32861 16899 32895
rect 28181 32861 28215 32895
rect 31033 32861 31067 32895
rect 31677 32861 31711 32895
rect 16957 32725 16991 32759
rect 28273 32725 28307 32759
rect 31125 32725 31159 32759
rect 31769 32725 31803 32759
rect 16957 32521 16991 32555
rect 1777 32385 1811 32419
rect 7389 32385 7423 32419
rect 16865 32385 16899 32419
rect 19625 32385 19659 32419
rect 20361 32385 20395 32419
rect 38301 32385 38335 32419
rect 1593 32181 1627 32215
rect 7481 32181 7515 32215
rect 19717 32181 19751 32215
rect 20453 32181 20487 32215
rect 38117 32181 38151 32215
rect 33885 31977 33919 32011
rect 32137 31773 32171 31807
rect 32229 31773 32263 31807
rect 34069 31773 34103 31807
rect 33885 30889 33919 30923
rect 1593 30821 1627 30855
rect 9413 30821 9447 30855
rect 25053 30821 25087 30855
rect 1777 30685 1811 30719
rect 6009 30685 6043 30719
rect 9321 30685 9355 30719
rect 9965 30685 9999 30719
rect 23489 30685 23523 30719
rect 24961 30685 24995 30719
rect 25881 30685 25915 30719
rect 27721 30685 27755 30719
rect 34069 30685 34103 30719
rect 6101 30549 6135 30583
rect 10057 30549 10091 30583
rect 23581 30549 23615 30583
rect 25973 30549 26007 30583
rect 27813 30549 27847 30583
rect 8125 30209 8159 30243
rect 29285 30209 29319 30243
rect 38301 30209 38335 30243
rect 8217 30005 8251 30039
rect 29377 30005 29411 30039
rect 38117 30005 38151 30039
rect 1593 29257 1627 29291
rect 5273 29257 5307 29291
rect 22661 29257 22695 29291
rect 1777 29121 1811 29155
rect 5457 29121 5491 29155
rect 11713 29121 11747 29155
rect 22569 29121 22603 29155
rect 38301 29121 38335 29155
rect 11805 28985 11839 29019
rect 38117 28985 38151 29019
rect 15577 28713 15611 28747
rect 16865 28713 16899 28747
rect 15485 28509 15519 28543
rect 16773 28509 16807 28543
rect 8769 28169 8803 28203
rect 11805 28169 11839 28203
rect 13645 28169 13679 28203
rect 29009 28169 29043 28203
rect 8677 28033 8711 28067
rect 11713 28033 11747 28067
rect 13553 28033 13587 28067
rect 28917 28033 28951 28067
rect 19533 27557 19567 27591
rect 1593 27421 1627 27455
rect 19441 27421 19475 27455
rect 33241 27421 33275 27455
rect 38025 27421 38059 27455
rect 1777 27285 1811 27319
rect 33333 27285 33367 27319
rect 38209 27285 38243 27319
rect 28089 27081 28123 27115
rect 8033 26945 8067 26979
rect 27997 26945 28031 26979
rect 8125 26741 8159 26775
rect 7665 25857 7699 25891
rect 17601 25857 17635 25891
rect 18521 25857 18555 25891
rect 7757 25653 7791 25687
rect 17693 25653 17727 25687
rect 18337 25653 18371 25687
rect 10149 25449 10183 25483
rect 1777 25245 1811 25279
rect 10057 25245 10091 25279
rect 15853 25245 15887 25279
rect 17601 25245 17635 25279
rect 19441 25245 19475 25279
rect 31677 25245 31711 25279
rect 32321 25245 32355 25279
rect 38025 25245 38059 25279
rect 1593 25109 1627 25143
rect 15945 25109 15979 25143
rect 17693 25109 17727 25143
rect 18613 25109 18647 25143
rect 19533 25109 19567 25143
rect 31769 25109 31803 25143
rect 32413 25109 32447 25143
rect 38209 25109 38243 25143
rect 15485 24769 15519 24803
rect 16313 24769 16347 24803
rect 17049 24769 17083 24803
rect 17693 24769 17727 24803
rect 18337 24769 18371 24803
rect 18981 24769 19015 24803
rect 20545 24769 20579 24803
rect 21005 24769 21039 24803
rect 18797 24701 18831 24735
rect 16865 24633 16899 24667
rect 18153 24633 18187 24667
rect 15577 24565 15611 24599
rect 16129 24565 16163 24599
rect 17509 24565 17543 24599
rect 19165 24565 19199 24599
rect 20361 24565 20395 24599
rect 21097 24565 21131 24599
rect 15393 24361 15427 24395
rect 16681 24361 16715 24395
rect 33517 24361 33551 24395
rect 16221 24225 16255 24259
rect 17141 24225 17175 24259
rect 17325 24225 17359 24259
rect 18245 24225 18279 24259
rect 1593 24157 1627 24191
rect 15577 24157 15611 24191
rect 16037 24157 16071 24191
rect 18429 24157 18463 24191
rect 21005 24157 21039 24191
rect 21833 24157 21867 24191
rect 33701 24157 33735 24191
rect 38301 24157 38335 24191
rect 18889 24089 18923 24123
rect 19533 24089 19567 24123
rect 19625 24089 19659 24123
rect 20177 24089 20211 24123
rect 21097 24089 21131 24123
rect 1777 24021 1811 24055
rect 17785 24021 17819 24055
rect 21649 24021 21683 24055
rect 38117 24021 38151 24055
rect 3985 23817 4019 23851
rect 14381 23817 14415 23851
rect 16313 23817 16347 23851
rect 19349 23749 19383 23783
rect 19901 23749 19935 23783
rect 20913 23749 20947 23783
rect 21465 23749 21499 23783
rect 4169 23681 4203 23715
rect 13645 23681 13679 23715
rect 14565 23681 14599 23715
rect 15209 23681 15243 23715
rect 15669 23681 15703 23715
rect 15853 23681 15887 23715
rect 17049 23681 17083 23715
rect 18061 23681 18095 23715
rect 22017 23681 22051 23715
rect 13001 23613 13035 23647
rect 16865 23613 16899 23647
rect 18245 23613 18279 23647
rect 19257 23613 19291 23647
rect 20821 23613 20855 23647
rect 22661 23613 22695 23647
rect 15025 23545 15059 23579
rect 18429 23545 18463 23579
rect 13737 23477 13771 23511
rect 17233 23477 17267 23511
rect 22109 23477 22143 23511
rect 15209 23273 15243 23307
rect 16865 23273 16899 23307
rect 18705 23273 18739 23307
rect 11989 23205 12023 23239
rect 15945 23205 15979 23239
rect 22569 23205 22603 23239
rect 16681 23137 16715 23171
rect 18061 23137 18095 23171
rect 18245 23137 18279 23171
rect 19901 23137 19935 23171
rect 20085 23137 20119 23171
rect 22201 23137 22235 23171
rect 22385 23137 22419 23171
rect 12173 23069 12207 23103
rect 12817 23069 12851 23103
rect 14565 23069 14599 23103
rect 15393 23069 15427 23103
rect 15853 23069 15887 23103
rect 16497 23069 16531 23103
rect 21741 23069 21775 23103
rect 14657 23001 14691 23035
rect 21097 23001 21131 23035
rect 21189 23001 21223 23035
rect 12633 22933 12667 22967
rect 13553 22933 13587 22967
rect 20545 22933 20579 22967
rect 5549 22729 5583 22763
rect 17233 22729 17267 22763
rect 21281 22729 21315 22763
rect 32965 22729 32999 22763
rect 18061 22661 18095 22695
rect 18613 22661 18647 22695
rect 1777 22593 1811 22627
rect 5457 22593 5491 22627
rect 9321 22593 9355 22627
rect 9965 22593 9999 22627
rect 13093 22593 13127 22627
rect 13553 22593 13587 22627
rect 14381 22593 14415 22627
rect 14841 22593 14875 22627
rect 15669 22593 15703 22627
rect 16313 22593 16347 22627
rect 17417 22593 17451 22627
rect 19717 22593 19751 22627
rect 22201 22593 22235 22627
rect 33149 22593 33183 22627
rect 10701 22525 10735 22559
rect 12265 22525 12299 22559
rect 17969 22525 18003 22559
rect 19533 22525 19567 22559
rect 20637 22525 20671 22559
rect 20821 22525 20855 22559
rect 9413 22457 9447 22491
rect 14933 22457 14967 22491
rect 16129 22457 16163 22491
rect 22017 22457 22051 22491
rect 1593 22389 1627 22423
rect 10057 22389 10091 22423
rect 12909 22389 12943 22423
rect 13645 22389 13679 22423
rect 14197 22389 14231 22423
rect 15485 22389 15519 22423
rect 19901 22389 19935 22423
rect 12357 22185 12391 22219
rect 17325 22185 17359 22219
rect 18429 22185 18463 22219
rect 21833 22185 21867 22219
rect 9873 22049 9907 22083
rect 13093 22049 13127 22083
rect 15577 22049 15611 22083
rect 16957 22049 16991 22083
rect 18245 22049 18279 22083
rect 20729 22049 20763 22083
rect 9321 21981 9355 22015
rect 9781 21981 9815 22015
rect 10609 21981 10643 22015
rect 11069 21981 11103 22015
rect 11897 21981 11931 22015
rect 12541 21981 12575 22015
rect 15025 21981 15059 22015
rect 16221 21981 16255 22015
rect 17141 21981 17175 22015
rect 18061 21981 18095 22015
rect 20177 21981 20211 22015
rect 22017 21981 22051 22015
rect 27445 21981 27479 22015
rect 27537 21981 27571 22015
rect 13185 21913 13219 21947
rect 13737 21913 13771 21947
rect 15669 21913 15703 21947
rect 20821 21913 20855 21947
rect 21373 21913 21407 21947
rect 38117 21913 38151 21947
rect 9137 21845 9171 21879
rect 10425 21845 10459 21879
rect 11161 21845 11195 21879
rect 11713 21845 11747 21879
rect 14841 21845 14875 21879
rect 19993 21845 20027 21879
rect 38209 21845 38243 21879
rect 8493 21641 8527 21675
rect 15485 21641 15519 21675
rect 16129 21641 16163 21675
rect 7941 21573 7975 21607
rect 10517 21573 10551 21607
rect 10609 21573 10643 21607
rect 13921 21573 13955 21607
rect 17049 21573 17083 21607
rect 17601 21573 17635 21607
rect 7849 21505 7883 21539
rect 8677 21505 8711 21539
rect 9321 21505 9355 21539
rect 9965 21505 9999 21539
rect 11989 21505 12023 21539
rect 12633 21505 12667 21539
rect 13277 21505 13311 21539
rect 15669 21505 15703 21539
rect 18797 21505 18831 21539
rect 19257 21505 19291 21539
rect 20453 21505 20487 21539
rect 22201 21505 22235 21539
rect 13829 21437 13863 21471
rect 14105 21437 14139 21471
rect 16957 21437 16991 21471
rect 19441 21437 19475 21471
rect 20637 21437 20671 21471
rect 9137 21369 9171 21403
rect 11069 21369 11103 21403
rect 11805 21369 11839 21403
rect 18613 21369 18647 21403
rect 22017 21369 22051 21403
rect 9781 21301 9815 21335
rect 12449 21301 12483 21335
rect 13093 21301 13127 21335
rect 19625 21301 19659 21335
rect 20821 21301 20855 21335
rect 6929 21097 6963 21131
rect 13737 21097 13771 21131
rect 16313 21097 16347 21131
rect 18797 21097 18831 21131
rect 19625 21097 19659 21131
rect 7757 21029 7791 21063
rect 10701 21029 10735 21063
rect 12633 21029 12667 21063
rect 14749 21029 14783 21063
rect 21097 21029 21131 21063
rect 22477 21029 22511 21063
rect 10517 20961 10551 20995
rect 12173 20961 12207 20995
rect 13093 20961 13127 20995
rect 13277 20961 13311 20995
rect 14381 20961 14415 20995
rect 14565 20961 14599 20995
rect 17601 20961 17635 20995
rect 20913 20961 20947 20995
rect 1777 20893 1811 20927
rect 7113 20893 7147 20927
rect 7941 20893 7975 20927
rect 8401 20893 8435 20927
rect 10333 20893 10367 20927
rect 11989 20893 12023 20927
rect 15945 20893 15979 20927
rect 16129 20893 16163 20927
rect 18705 20893 18739 20927
rect 19809 20893 19843 20927
rect 20729 20893 20763 20927
rect 22017 20893 22051 20927
rect 22661 20893 22695 20927
rect 23121 20893 23155 20927
rect 25881 20893 25915 20927
rect 38025 20893 38059 20927
rect 9689 20825 9723 20859
rect 17141 20825 17175 20859
rect 17233 20825 17267 20859
rect 1593 20757 1627 20791
rect 21833 20757 21867 20791
rect 23213 20757 23247 20791
rect 25973 20757 26007 20791
rect 38209 20757 38243 20791
rect 7573 20553 7607 20587
rect 14473 20553 14507 20587
rect 22017 20553 22051 20587
rect 10333 20485 10367 20519
rect 10885 20485 10919 20519
rect 12173 20485 12207 20519
rect 13277 20485 13311 20519
rect 13369 20485 13403 20519
rect 17049 20485 17083 20519
rect 18889 20485 18923 20519
rect 19993 20485 20027 20519
rect 20085 20485 20119 20519
rect 20637 20485 20671 20519
rect 6929 20417 6963 20451
rect 7757 20417 7791 20451
rect 8217 20417 8251 20451
rect 9045 20417 9079 20451
rect 9689 20417 9723 20451
rect 14657 20417 14691 20451
rect 15117 20417 15151 20451
rect 18061 20417 18095 20451
rect 21097 20417 21131 20451
rect 22845 20417 22879 20451
rect 23489 20417 23523 20451
rect 10241 20349 10275 20383
rect 12081 20349 12115 20383
rect 15301 20349 15335 20383
rect 16957 20349 16991 20383
rect 17233 20349 17267 20383
rect 18797 20349 18831 20383
rect 8861 20281 8895 20315
rect 12633 20281 12667 20315
rect 13829 20281 13863 20315
rect 19349 20281 19383 20315
rect 7021 20213 7055 20247
rect 8309 20213 8343 20247
rect 9505 20213 9539 20247
rect 15761 20213 15795 20247
rect 18153 20213 18187 20247
rect 21189 20213 21223 20247
rect 22661 20213 22695 20247
rect 23305 20213 23339 20247
rect 8401 20009 8435 20043
rect 10333 20009 10367 20043
rect 11345 20009 11379 20043
rect 17601 20009 17635 20043
rect 19901 20009 19935 20043
rect 21097 20009 21131 20043
rect 9689 19873 9723 19907
rect 9873 19873 9907 19907
rect 12081 19873 12115 19907
rect 12541 19873 12575 19907
rect 15117 19873 15151 19907
rect 16221 19873 16255 19907
rect 16405 19873 16439 19907
rect 18245 19873 18279 19907
rect 20729 19873 20763 19907
rect 20913 19873 20947 19907
rect 21925 19873 21959 19907
rect 7113 19805 7147 19839
rect 7941 19805 7975 19839
rect 8585 19805 8619 19839
rect 11529 19805 11563 19839
rect 14565 19805 14599 19839
rect 15761 19805 15795 19839
rect 17509 19805 17543 19839
rect 18429 19805 18463 19839
rect 19533 19805 19567 19839
rect 19717 19805 19751 19839
rect 23029 19805 23063 19839
rect 29745 19805 29779 19839
rect 7205 19737 7239 19771
rect 12173 19737 12207 19771
rect 15209 19737 15243 19771
rect 22017 19737 22051 19771
rect 22569 19737 22603 19771
rect 7757 19669 7791 19703
rect 13553 19669 13587 19703
rect 14381 19669 14415 19703
rect 16865 19669 16899 19703
rect 18889 19669 18923 19703
rect 23121 19669 23155 19703
rect 29837 19669 29871 19703
rect 1593 19465 1627 19499
rect 6745 19465 6779 19499
rect 7389 19465 7423 19499
rect 12357 19465 12391 19499
rect 13645 19465 13679 19499
rect 14657 19465 14691 19499
rect 18705 19465 18739 19499
rect 1777 19329 1811 19363
rect 5825 19329 5859 19363
rect 5917 19329 5951 19363
rect 6929 19329 6963 19363
rect 7573 19329 7607 19363
rect 8033 19329 8067 19363
rect 8125 19329 8159 19363
rect 8861 19329 8895 19363
rect 9505 19329 9539 19363
rect 13001 19329 13035 19363
rect 17049 19329 17083 19363
rect 17693 19329 17727 19363
rect 18889 19329 18923 19363
rect 19993 19329 20027 19363
rect 20729 19329 20763 19363
rect 21373 19329 21407 19363
rect 22661 19329 22695 19363
rect 23305 19329 23339 19363
rect 9965 19261 9999 19295
rect 10150 19261 10184 19295
rect 11713 19261 11747 19295
rect 11897 19261 11931 19295
rect 13185 19261 13219 19295
rect 15301 19261 15335 19295
rect 15485 19261 15519 19295
rect 17233 19261 17267 19295
rect 19349 19261 19383 19295
rect 19533 19261 19567 19295
rect 20913 19261 20947 19295
rect 22017 19261 22051 19295
rect 22201 19261 22235 19295
rect 8677 19193 8711 19227
rect 10333 19193 10367 19227
rect 23121 19193 23155 19227
rect 9321 19125 9355 19159
rect 15945 19125 15979 19159
rect 7205 18921 7239 18955
rect 9965 18921 9999 18955
rect 10517 18921 10551 18955
rect 15025 18921 15059 18955
rect 15669 18921 15703 18955
rect 16313 18921 16347 18955
rect 18889 18921 18923 18955
rect 23029 18921 23063 18955
rect 33609 18921 33643 18955
rect 13553 18853 13587 18887
rect 17601 18853 17635 18887
rect 9321 18785 9355 18819
rect 11253 18785 11287 18819
rect 17049 18785 17083 18819
rect 19533 18785 19567 18819
rect 20821 18785 20855 18819
rect 21649 18785 21683 18819
rect 6653 18717 6687 18751
rect 7113 18717 7147 18751
rect 7757 18717 7791 18751
rect 8401 18717 8435 18751
rect 9505 18717 9539 18751
rect 10425 18717 10459 18751
rect 11069 18717 11103 18751
rect 12265 18717 12299 18751
rect 14565 18717 14599 18751
rect 15209 18717 15243 18751
rect 15853 18717 15887 18751
rect 16497 18717 16531 18751
rect 18245 18717 18279 18751
rect 18429 18717 18463 18751
rect 22937 18717 22971 18751
rect 33793 18717 33827 18751
rect 13001 18649 13035 18683
rect 13093 18649 13127 18683
rect 17141 18649 17175 18683
rect 20545 18649 20579 18683
rect 20637 18649 20671 18683
rect 6469 18581 6503 18615
rect 7849 18581 7883 18615
rect 8493 18581 8527 18615
rect 11713 18581 11747 18615
rect 12357 18581 12391 18615
rect 14381 18581 14415 18615
rect 22293 18581 22327 18615
rect 7205 18377 7239 18411
rect 9137 18377 9171 18411
rect 15117 18377 15151 18411
rect 18429 18377 18463 18411
rect 19625 18377 19659 18411
rect 21281 18377 21315 18411
rect 22017 18377 22051 18411
rect 33425 18377 33459 18411
rect 10609 18309 10643 18343
rect 17141 18309 17175 18343
rect 17693 18309 17727 18343
rect 20269 18309 20303 18343
rect 20821 18309 20855 18343
rect 1777 18241 1811 18275
rect 7389 18241 7423 18275
rect 8033 18241 8067 18275
rect 8677 18241 8711 18275
rect 9321 18241 9355 18275
rect 9965 18241 9999 18275
rect 12265 18241 12299 18275
rect 12909 18241 12943 18275
rect 16129 18241 16163 18275
rect 18337 18241 18371 18275
rect 21465 18241 21499 18275
rect 22201 18241 22235 18275
rect 22661 18241 22695 18275
rect 23305 18241 23339 18275
rect 33333 18241 33367 18275
rect 10517 18173 10551 18207
rect 12449 18173 12483 18207
rect 13369 18173 13403 18207
rect 13553 18173 13587 18207
rect 14473 18173 14507 18207
rect 14657 18173 14691 18207
rect 17049 18173 17083 18207
rect 18981 18173 19015 18207
rect 19165 18173 19199 18207
rect 20177 18173 20211 18207
rect 7849 18105 7883 18139
rect 9781 18105 9815 18139
rect 11069 18105 11103 18139
rect 13737 18105 13771 18139
rect 1593 18037 1627 18071
rect 8493 18037 8527 18071
rect 16221 18037 16255 18071
rect 22753 18037 22787 18071
rect 23397 18037 23431 18071
rect 8401 17833 8435 17867
rect 9229 17833 9263 17867
rect 11713 17833 11747 17867
rect 16221 17833 16255 17867
rect 19717 17833 19751 17867
rect 17325 17765 17359 17799
rect 21005 17765 21039 17799
rect 9965 17697 9999 17731
rect 10241 17697 10275 17731
rect 11253 17697 11287 17731
rect 12725 17697 12759 17731
rect 13001 17697 13035 17731
rect 17049 17697 17083 17731
rect 18337 17697 18371 17731
rect 20453 17697 20487 17731
rect 5181 17629 5215 17663
rect 7297 17629 7331 17663
rect 8585 17629 8619 17663
rect 9413 17629 9447 17663
rect 11069 17629 11103 17663
rect 14289 17629 14323 17663
rect 14473 17629 14507 17663
rect 16405 17629 16439 17663
rect 16865 17629 16899 17663
rect 18153 17629 18187 17663
rect 19901 17629 19935 17663
rect 21557 17629 21591 17663
rect 21741 17629 21775 17663
rect 22661 17629 22695 17663
rect 23489 17629 23523 17663
rect 5273 17561 5307 17595
rect 10057 17561 10091 17595
rect 12817 17561 12851 17595
rect 14933 17561 14967 17595
rect 20545 17561 20579 17595
rect 7113 17493 7147 17527
rect 7757 17493 7791 17527
rect 15577 17493 15611 17527
rect 18797 17493 18831 17527
rect 22201 17493 22235 17527
rect 22753 17493 22787 17527
rect 23305 17493 23339 17527
rect 7389 17289 7423 17323
rect 8033 17289 8067 17323
rect 16957 17289 16991 17323
rect 19441 17289 19475 17323
rect 21097 17289 21131 17323
rect 12449 17221 12483 17255
rect 13001 17221 13035 17255
rect 15301 17221 15335 17255
rect 20085 17221 20119 17255
rect 6929 17153 6963 17187
rect 7573 17153 7607 17187
rect 8217 17153 8251 17187
rect 8677 17153 8711 17187
rect 10701 17153 10735 17187
rect 13461 17153 13495 17187
rect 13645 17153 13679 17187
rect 15853 17153 15887 17187
rect 17141 17153 17175 17187
rect 17601 17153 17635 17187
rect 21281 17153 21315 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 38025 17153 38059 17187
rect 9321 17085 9355 17119
rect 9505 17085 9539 17119
rect 10517 17085 10551 17119
rect 12357 17085 12391 17119
rect 15209 17085 15243 17119
rect 17785 17085 17819 17119
rect 18797 17085 18831 17119
rect 18981 17085 19015 17119
rect 19993 17085 20027 17119
rect 23121 17085 23155 17119
rect 23305 17085 23339 17119
rect 6745 17017 6779 17051
rect 13829 17017 13863 17051
rect 20545 17017 20579 17051
rect 38209 17017 38243 17051
rect 8769 16949 8803 16983
rect 9689 16949 9723 16983
rect 11161 16949 11195 16983
rect 17969 16949 18003 16983
rect 22661 16949 22695 16983
rect 23489 16949 23523 16983
rect 8401 16745 8435 16779
rect 9689 16745 9723 16779
rect 21465 16745 21499 16779
rect 23305 16745 23339 16779
rect 7757 16677 7791 16711
rect 15209 16677 15243 16711
rect 17417 16677 17451 16711
rect 20821 16677 20855 16711
rect 9321 16609 9355 16643
rect 11161 16609 11195 16643
rect 12357 16609 12391 16643
rect 12725 16609 12759 16643
rect 16129 16609 16163 16643
rect 17233 16609 17267 16643
rect 18245 16609 18279 16643
rect 18613 16609 18647 16643
rect 20269 16609 20303 16643
rect 22661 16609 22695 16643
rect 6469 16541 6503 16575
rect 6561 16541 6595 16575
rect 7113 16541 7147 16575
rect 7941 16541 7975 16575
rect 8585 16541 8619 16575
rect 9137 16541 9171 16575
rect 10609 16541 10643 16575
rect 13737 16541 13771 16575
rect 14841 16541 14875 16575
rect 15025 16541 15059 16575
rect 15945 16541 15979 16575
rect 16589 16541 16623 16575
rect 17049 16541 17083 16575
rect 19533 16541 19567 16575
rect 21373 16541 21407 16575
rect 22017 16541 22051 16575
rect 23489 16541 23523 16575
rect 27077 16541 27111 16575
rect 33793 16541 33827 16575
rect 11253 16473 11287 16507
rect 11805 16473 11839 16507
rect 12449 16473 12483 16507
rect 18337 16473 18371 16507
rect 19625 16473 19659 16507
rect 20361 16473 20395 16507
rect 27169 16473 27203 16507
rect 7205 16405 7239 16439
rect 10425 16405 10459 16439
rect 13553 16405 13587 16439
rect 33609 16405 33643 16439
rect 7113 16201 7147 16235
rect 9689 16201 9723 16235
rect 15209 16201 15243 16235
rect 16313 16201 16347 16235
rect 17509 16201 17543 16235
rect 22661 16201 22695 16235
rect 19165 16133 19199 16167
rect 19257 16133 19291 16167
rect 20913 16133 20947 16167
rect 21465 16133 21499 16167
rect 1593 16065 1627 16099
rect 7297 16065 7331 16099
rect 7757 16065 7791 16099
rect 8585 16065 8619 16099
rect 9873 16065 9907 16099
rect 10333 16065 10367 16099
rect 11161 16065 11195 16099
rect 15853 16065 15887 16099
rect 18153 16065 18187 16099
rect 22845 16065 22879 16099
rect 24133 16065 24167 16099
rect 38301 16065 38335 16099
rect 9045 15997 9079 16031
rect 11897 15997 11931 16031
rect 12081 15997 12115 16031
rect 13001 15997 13035 16031
rect 13185 15997 13219 16031
rect 14565 15997 14599 16031
rect 14749 15997 14783 16031
rect 15669 15997 15703 16031
rect 16865 15997 16899 16031
rect 17049 15997 17083 16031
rect 17969 15997 18003 16031
rect 20821 15997 20855 16031
rect 22017 15997 22051 16031
rect 23305 15997 23339 16031
rect 24593 15997 24627 16031
rect 10425 15929 10459 15963
rect 13369 15929 13403 15963
rect 18337 15929 18371 15963
rect 19717 15929 19751 15963
rect 1777 15861 1811 15895
rect 7849 15861 7883 15895
rect 8401 15861 8435 15895
rect 10977 15861 11011 15895
rect 12541 15861 12575 15895
rect 23949 15861 23983 15895
rect 38117 15861 38151 15895
rect 8401 15657 8435 15691
rect 16681 15657 16715 15691
rect 18705 15657 18739 15691
rect 24593 15657 24627 15691
rect 12081 15589 12115 15623
rect 7389 15521 7423 15555
rect 10609 15521 10643 15555
rect 11897 15521 11931 15555
rect 12909 15521 12943 15555
rect 13185 15521 13219 15555
rect 14657 15521 14691 15555
rect 16037 15521 16071 15555
rect 17325 15521 17359 15555
rect 19993 15521 20027 15555
rect 21649 15521 21683 15555
rect 23121 15521 23155 15555
rect 23305 15521 23339 15555
rect 7297 15453 7331 15487
rect 8585 15453 8619 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 10793 15453 10827 15487
rect 11713 15453 11747 15487
rect 16221 15453 16255 15487
rect 18889 15453 18923 15487
rect 20177 15453 20211 15487
rect 21833 15453 21867 15487
rect 24777 15453 24811 15487
rect 25421 15453 25455 15487
rect 11253 15385 11287 15419
rect 12994 15385 13028 15419
rect 14381 15385 14415 15419
rect 14473 15385 14507 15419
rect 17417 15385 17451 15419
rect 17969 15385 18003 15419
rect 9781 15317 9815 15351
rect 20637 15317 20671 15351
rect 22293 15317 22327 15351
rect 23765 15317 23799 15351
rect 25237 15317 25271 15351
rect 10885 15113 10919 15147
rect 11805 15113 11839 15147
rect 15577 15113 15611 15147
rect 18889 15113 18923 15147
rect 20177 15113 20211 15147
rect 20637 15113 20671 15147
rect 22109 15113 22143 15147
rect 25789 15113 25823 15147
rect 9045 15045 9079 15079
rect 17509 15045 17543 15079
rect 17601 15045 17635 15079
rect 7021 14977 7055 15011
rect 7849 14977 7883 15011
rect 8493 14977 8527 15011
rect 8953 14977 8987 15011
rect 9781 14977 9815 15011
rect 10425 14977 10459 15011
rect 11713 14977 11747 15011
rect 12357 14977 12391 15011
rect 15485 14977 15519 15011
rect 16313 14977 16347 15011
rect 18153 14977 18187 15011
rect 19073 14977 19107 15011
rect 20821 14977 20855 15011
rect 21465 14977 21499 15011
rect 22017 14977 22051 15011
rect 24041 14977 24075 15011
rect 24225 14977 24259 15011
rect 25145 14977 25179 15011
rect 25973 14977 26007 15011
rect 33057 14977 33091 15011
rect 10241 14909 10275 14943
rect 12541 14909 12575 14943
rect 13921 14909 13955 14943
rect 14105 14909 14139 14943
rect 19533 14909 19567 14943
rect 19717 14909 19751 14943
rect 22937 14909 22971 14943
rect 23121 14909 23155 14943
rect 25237 14909 25271 14943
rect 7665 14841 7699 14875
rect 9597 14841 9631 14875
rect 12725 14841 12759 14875
rect 14289 14841 14323 14875
rect 21281 14841 21315 14875
rect 7113 14773 7147 14807
rect 8309 14773 8343 14807
rect 16129 14773 16163 14807
rect 23581 14773 23615 14807
rect 24409 14773 24443 14807
rect 33149 14773 33183 14807
rect 4813 14569 4847 14603
rect 8493 14569 8527 14603
rect 12357 14569 12391 14603
rect 13553 14569 13587 14603
rect 14749 14569 14783 14603
rect 16681 14569 16715 14603
rect 17233 14569 17267 14603
rect 18153 14569 18187 14603
rect 18705 14569 18739 14603
rect 20361 14569 20395 14603
rect 24961 14569 24995 14603
rect 1593 14501 1627 14535
rect 10241 14501 10275 14535
rect 11621 14501 11655 14535
rect 16037 14501 16071 14535
rect 21005 14501 21039 14535
rect 23213 14501 23247 14535
rect 26341 14501 26375 14535
rect 7849 14433 7883 14467
rect 9781 14433 9815 14467
rect 10977 14433 11011 14467
rect 19625 14433 19659 14467
rect 22845 14433 22879 14467
rect 24593 14433 24627 14467
rect 24777 14433 24811 14467
rect 27077 14433 27111 14467
rect 1777 14365 1811 14399
rect 2329 14365 2363 14399
rect 4997 14365 5031 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 9597 14365 9631 14399
rect 11805 14365 11839 14399
rect 12265 14365 12299 14399
rect 13093 14365 13127 14399
rect 13737 14365 13771 14399
rect 14657 14365 14691 14399
rect 15485 14365 15519 14399
rect 15945 14365 15979 14399
rect 16589 14365 16623 14399
rect 17417 14365 17451 14399
rect 18061 14365 18095 14399
rect 18889 14365 18923 14399
rect 20545 14365 20579 14399
rect 21189 14365 21223 14399
rect 22017 14365 22051 14399
rect 23029 14365 23063 14399
rect 25881 14365 25915 14399
rect 26525 14365 26559 14399
rect 26985 14365 27019 14399
rect 38025 14365 38059 14399
rect 2421 14229 2455 14263
rect 12909 14229 12943 14263
rect 15301 14229 15335 14263
rect 21833 14229 21867 14263
rect 25697 14229 25731 14263
rect 38209 14229 38243 14263
rect 7205 14025 7239 14059
rect 7757 14025 7791 14059
rect 9045 14025 9079 14059
rect 9689 14025 9723 14059
rect 10333 14025 10367 14059
rect 11069 14025 11103 14059
rect 13369 14025 13403 14059
rect 14013 14025 14047 14059
rect 14749 14025 14783 14059
rect 18429 14025 18463 14059
rect 19533 14025 19567 14059
rect 20085 14025 20119 14059
rect 21281 14025 21315 14059
rect 25881 14025 25915 14059
rect 8493 13957 8527 13991
rect 12449 13957 12483 13991
rect 24225 13957 24259 13991
rect 1593 13889 1627 13923
rect 2237 13889 2271 13923
rect 2973 13889 3007 13923
rect 3617 13889 3651 13923
rect 7113 13889 7147 13923
rect 7941 13889 7975 13923
rect 8401 13889 8435 13923
rect 9229 13889 9263 13923
rect 9873 13889 9907 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 11989 13889 12023 13923
rect 13553 13889 13587 13923
rect 14197 13889 14231 13923
rect 14657 13889 14691 13923
rect 18613 13889 18647 13923
rect 19441 13889 19475 13923
rect 20269 13889 20303 13923
rect 21465 13889 21499 13923
rect 22201 13889 22235 13923
rect 25421 13889 25455 13923
rect 26065 13889 26099 13923
rect 2329 13821 2363 13855
rect 3065 13821 3099 13855
rect 3709 13821 3743 13855
rect 11805 13821 11839 13855
rect 15301 13821 15335 13855
rect 15485 13821 15519 13855
rect 15945 13821 15979 13855
rect 17049 13821 17083 13855
rect 17233 13821 17267 13855
rect 22017 13821 22051 13855
rect 23121 13821 23155 13855
rect 24133 13821 24167 13855
rect 24777 13821 24811 13855
rect 1685 13685 1719 13719
rect 17417 13685 17451 13719
rect 22661 13685 22695 13719
rect 25237 13685 25271 13719
rect 7113 13481 7147 13515
rect 8401 13481 8435 13515
rect 11437 13481 11471 13515
rect 12265 13481 12299 13515
rect 13001 13481 13035 13515
rect 19533 13481 19567 13515
rect 22477 13481 22511 13515
rect 23581 13481 23615 13515
rect 1593 13413 1627 13447
rect 9505 13413 9539 13447
rect 15853 13413 15887 13447
rect 17969 13413 18003 13447
rect 18705 13413 18739 13447
rect 25881 13413 25915 13447
rect 2697 13345 2731 13379
rect 10241 13345 10275 13379
rect 16497 13345 16531 13379
rect 16681 13345 16715 13379
rect 17601 13345 17635 13379
rect 22017 13345 22051 13379
rect 24961 13345 24995 13379
rect 1777 13277 1811 13311
rect 2605 13277 2639 13311
rect 3249 13277 3283 13311
rect 4169 13277 4203 13311
rect 7297 13277 7331 13311
rect 7941 13277 7975 13311
rect 8585 13277 8619 13311
rect 9689 13277 9723 13311
rect 10149 13277 10183 13311
rect 10793 13277 10827 13311
rect 11621 13277 11655 13311
rect 12449 13277 12483 13311
rect 12909 13277 12943 13311
rect 13737 13277 13771 13311
rect 14841 13277 14875 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 17785 13277 17819 13311
rect 18889 13277 18923 13311
rect 19717 13277 19751 13311
rect 20637 13277 20671 13311
rect 21833 13277 21867 13311
rect 23213 13277 23247 13311
rect 23397 13277 23431 13311
rect 25789 13277 25823 13311
rect 26617 13277 26651 13311
rect 3341 13209 3375 13243
rect 24685 13209 24719 13243
rect 24777 13209 24811 13243
rect 4261 13141 4295 13175
rect 7757 13141 7791 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 14657 13141 14691 13175
rect 17141 13141 17175 13175
rect 20453 13141 20487 13175
rect 21097 13141 21131 13175
rect 26433 13141 26467 13175
rect 5825 12937 5859 12971
rect 11069 12937 11103 12971
rect 12357 12937 12391 12971
rect 13093 12937 13127 12971
rect 16957 12937 16991 12971
rect 18889 12937 18923 12971
rect 20177 12937 20211 12971
rect 26157 12937 26191 12971
rect 32597 12937 32631 12971
rect 7665 12869 7699 12903
rect 22201 12869 22235 12903
rect 23397 12869 23431 12903
rect 25605 12869 25639 12903
rect 1777 12801 1811 12835
rect 2421 12801 2455 12835
rect 3249 12801 3283 12835
rect 4077 12801 4111 12835
rect 4813 12801 4847 12835
rect 6009 12801 6043 12835
rect 6929 12801 6963 12835
rect 7573 12801 7607 12835
rect 8217 12801 8251 12835
rect 8309 12801 8343 12835
rect 10609 12801 10643 12835
rect 12265 12801 12299 12835
rect 13001 12801 13035 12835
rect 13829 12801 13863 12835
rect 14473 12801 14507 12835
rect 15393 12801 15427 12835
rect 17141 12801 17175 12835
rect 18797 12801 18831 12835
rect 19533 12801 19567 12835
rect 20361 12801 20395 12835
rect 20821 12801 20855 12835
rect 21005 12801 21039 12835
rect 24409 12801 24443 12835
rect 25513 12801 25547 12835
rect 26341 12801 26375 12835
rect 32781 12801 32815 12835
rect 38025 12801 38059 12835
rect 4905 12733 4939 12767
rect 8861 12733 8895 12767
rect 9045 12733 9079 12767
rect 10425 12733 10459 12767
rect 14289 12733 14323 12767
rect 15577 12733 15611 12767
rect 17693 12733 17727 12767
rect 17877 12733 17911 12767
rect 22109 12733 22143 12767
rect 23305 12733 23339 12767
rect 23581 12733 23615 12767
rect 24593 12733 24627 12767
rect 1593 12665 1627 12699
rect 3341 12665 3375 12699
rect 7021 12665 7055 12699
rect 13645 12665 13679 12699
rect 18061 12665 18095 12699
rect 22661 12665 22695 12699
rect 2237 12597 2271 12631
rect 3893 12597 3927 12631
rect 9505 12597 9539 12631
rect 14657 12597 14691 12631
rect 16037 12597 16071 12631
rect 19625 12597 19659 12631
rect 21189 12597 21223 12631
rect 24869 12597 24903 12631
rect 38209 12597 38243 12631
rect 6561 12393 6595 12427
rect 15945 12393 15979 12427
rect 17601 12393 17635 12427
rect 18245 12393 18279 12427
rect 21005 12393 21039 12427
rect 37841 12393 37875 12427
rect 9781 12325 9815 12359
rect 11529 12325 11563 12359
rect 23857 12325 23891 12359
rect 24961 12325 24995 12359
rect 5273 12257 5307 12291
rect 7849 12257 7883 12291
rect 9321 12257 9355 12291
rect 11345 12257 11379 12291
rect 14381 12257 14415 12291
rect 16497 12257 16531 12291
rect 16681 12257 16715 12291
rect 20085 12257 20119 12291
rect 20821 12257 20855 12291
rect 23213 12257 23247 12291
rect 24593 12257 24627 12291
rect 1777 12189 1811 12223
rect 2237 12189 2271 12223
rect 2881 12189 2915 12223
rect 3985 12189 4019 12223
rect 5181 12189 5215 12223
rect 5825 12189 5859 12223
rect 6469 12189 6503 12223
rect 7297 12189 7331 12223
rect 7757 12189 7791 12223
rect 8585 12189 8619 12223
rect 9137 12189 9171 12223
rect 10701 12189 10735 12223
rect 11161 12189 11195 12223
rect 13645 12189 13679 12223
rect 15853 12189 15887 12223
rect 17785 12189 17819 12223
rect 18429 12189 18463 12223
rect 19993 12189 20027 12223
rect 20637 12189 20671 12223
rect 22109 12189 22143 12223
rect 22293 12189 22327 12223
rect 23397 12189 23431 12223
rect 24777 12189 24811 12223
rect 36921 12189 36955 12223
rect 37013 12189 37047 12223
rect 38025 12189 38059 12223
rect 4077 12121 4111 12155
rect 12357 12121 12391 12155
rect 12449 12121 12483 12155
rect 13001 12121 13035 12155
rect 14473 12121 14507 12155
rect 15025 12121 15059 12155
rect 25697 12121 25731 12155
rect 1593 12053 1627 12087
rect 2329 12053 2363 12087
rect 2973 12053 3007 12087
rect 5917 12053 5951 12087
rect 7113 12053 7147 12087
rect 8401 12053 8435 12087
rect 10517 12053 10551 12087
rect 13461 12053 13495 12087
rect 17141 12053 17175 12087
rect 22753 12053 22787 12087
rect 7113 11849 7147 11883
rect 9689 11849 9723 11883
rect 17141 11849 17175 11883
rect 18153 11849 18187 11883
rect 21097 11849 21131 11883
rect 22017 11849 22051 11883
rect 25237 11849 25271 11883
rect 25881 11849 25915 11883
rect 12633 11781 12667 11815
rect 14289 11781 14323 11815
rect 23029 11781 23063 11815
rect 24225 11781 24259 11815
rect 1777 11713 1811 11747
rect 2421 11713 2455 11747
rect 5181 11713 5215 11747
rect 5825 11713 5859 11747
rect 7297 11713 7331 11747
rect 7757 11713 7791 11747
rect 8585 11713 8619 11747
rect 9229 11713 9263 11747
rect 10517 11713 10551 11747
rect 10977 11713 11011 11747
rect 11069 11713 11103 11747
rect 14013 11713 14047 11747
rect 17325 11713 17359 11747
rect 18337 11713 18371 11747
rect 18797 11713 18831 11747
rect 19993 11713 20027 11747
rect 20637 11713 20671 11747
rect 22201 11713 22235 11747
rect 25421 11713 25455 11747
rect 26065 11713 26099 11747
rect 2881 11645 2915 11679
rect 3157 11645 3191 11679
rect 11805 11645 11839 11679
rect 12541 11645 12575 11679
rect 12817 11645 12851 11679
rect 20453 11645 20487 11679
rect 22937 11645 22971 11679
rect 23581 11645 23615 11679
rect 24133 11645 24167 11679
rect 1593 11577 1627 11611
rect 5273 11577 5307 11611
rect 5917 11577 5951 11611
rect 8401 11577 8435 11611
rect 9045 11577 9079 11611
rect 10333 11577 10367 11611
rect 24685 11577 24719 11611
rect 2237 11509 2271 11543
rect 4629 11509 4663 11543
rect 7849 11509 7883 11543
rect 15761 11509 15795 11543
rect 18889 11509 18923 11543
rect 19809 11509 19843 11543
rect 1593 11305 1627 11339
rect 4248 11305 4282 11339
rect 9321 11305 9355 11339
rect 16037 11305 16071 11339
rect 21833 11305 21867 11339
rect 24593 11305 24627 11339
rect 25329 11305 25363 11339
rect 25973 11305 26007 11339
rect 2605 11237 2639 11271
rect 5733 11237 5767 11271
rect 10609 11237 10643 11271
rect 13553 11237 13587 11271
rect 19717 11237 19751 11271
rect 38209 11237 38243 11271
rect 6285 11169 6319 11203
rect 9965 11169 9999 11203
rect 11345 11169 11379 11203
rect 12817 11169 12851 11203
rect 16589 11169 16623 11203
rect 16865 11169 16899 11203
rect 20361 11169 20395 11203
rect 22385 11169 22419 11203
rect 1777 11101 1811 11135
rect 2789 11101 2823 11135
rect 3249 11101 3283 11135
rect 3985 11101 4019 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 9505 11101 9539 11135
rect 10149 11101 10183 11135
rect 11069 11101 11103 11135
rect 13737 11101 13771 11135
rect 14289 11101 14323 11135
rect 17693 11101 17727 11135
rect 19901 11101 19935 11135
rect 20545 11101 20579 11135
rect 21741 11101 21775 11135
rect 22569 11101 22603 11135
rect 23673 11101 23707 11135
rect 24777 11101 24811 11135
rect 25237 11101 25271 11135
rect 25881 11101 25915 11135
rect 26985 11101 27019 11135
rect 38025 11101 38059 11135
rect 3341 11033 3375 11067
rect 7113 11033 7147 11067
rect 14565 11033 14599 11067
rect 16681 11033 16715 11067
rect 17785 11033 17819 11067
rect 18337 11033 18371 11067
rect 21005 11033 21039 11067
rect 23029 11033 23063 11067
rect 27077 11033 27111 11067
rect 8585 10965 8619 10999
rect 23489 10965 23523 10999
rect 1593 10761 1627 10795
rect 7021 10761 7055 10795
rect 11069 10761 11103 10795
rect 15945 10761 15979 10795
rect 20177 10761 20211 10795
rect 23765 10761 23799 10795
rect 25053 10761 25087 10795
rect 16957 10693 16991 10727
rect 22661 10693 22695 10727
rect 22753 10693 22787 10727
rect 25605 10693 25639 10727
rect 1777 10625 1811 10659
rect 2605 10625 2639 10659
rect 5825 10625 5859 10659
rect 6929 10625 6963 10659
rect 7573 10625 7607 10659
rect 10241 10625 10275 10659
rect 10977 10625 11011 10659
rect 11989 10625 12023 10659
rect 20361 10625 20395 10659
rect 21005 10625 21039 10659
rect 23305 10625 23339 10659
rect 23949 10625 23983 10659
rect 25513 10625 25547 10659
rect 3065 10557 3099 10591
rect 3341 10557 3375 10591
rect 8217 10557 8251 10591
rect 8493 10557 8527 10591
rect 12265 10557 12299 10591
rect 14197 10557 14231 10591
rect 14473 10557 14507 10591
rect 16865 10557 16899 10591
rect 17141 10557 17175 10591
rect 18613 10557 18647 10591
rect 18797 10557 18831 10591
rect 19533 10557 19567 10591
rect 24409 10557 24443 10591
rect 24593 10557 24627 10591
rect 5917 10489 5951 10523
rect 2421 10421 2455 10455
rect 4813 10421 4847 10455
rect 7665 10421 7699 10455
rect 13737 10421 13771 10455
rect 17785 10421 17819 10455
rect 18337 10421 18371 10455
rect 20821 10421 20855 10455
rect 1948 10217 1982 10251
rect 3433 10217 3467 10251
rect 9400 10217 9434 10251
rect 22753 10217 22787 10251
rect 23397 10217 23431 10251
rect 24685 10217 24719 10251
rect 25329 10217 25363 10251
rect 34897 10217 34931 10251
rect 13369 10149 13403 10183
rect 1685 10081 1719 10115
rect 4537 10081 4571 10115
rect 6837 10081 6871 10115
rect 9137 10081 9171 10115
rect 11621 10081 11655 10115
rect 11897 10081 11931 10115
rect 17693 10081 17727 10115
rect 17969 10081 18003 10115
rect 19533 10081 19567 10115
rect 19809 10081 19843 10115
rect 21005 10081 21039 10115
rect 4261 10013 4295 10047
rect 6561 10013 6595 10047
rect 8585 10013 8619 10047
rect 14289 10013 14323 10047
rect 16957 10013 16991 10047
rect 20821 10013 20855 10047
rect 22293 10013 22327 10047
rect 22937 10013 22971 10047
rect 23581 10013 23615 10047
rect 24593 10013 24627 10047
rect 25237 10013 25271 10047
rect 34345 10013 34379 10047
rect 35081 10013 35115 10047
rect 11161 9945 11195 9979
rect 14565 9945 14599 9979
rect 17785 9945 17819 9979
rect 19618 9945 19652 9979
rect 6009 9877 6043 9911
rect 16037 9877 16071 9911
rect 17049 9877 17083 9911
rect 21465 9877 21499 9911
rect 22109 9877 22143 9911
rect 34161 9877 34195 9911
rect 8677 9673 8711 9707
rect 20913 9673 20947 9707
rect 2421 9605 2455 9639
rect 9413 9605 9447 9639
rect 11161 9605 11195 9639
rect 14013 9605 14047 9639
rect 14749 9605 14783 9639
rect 17049 9605 17083 9639
rect 19257 9605 19291 9639
rect 22477 9605 22511 9639
rect 23949 9605 23983 9639
rect 27537 9605 27571 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 2973 9537 3007 9571
rect 3617 9537 3651 9571
rect 11989 9537 12023 9571
rect 20453 9537 20487 9571
rect 22385 9537 22419 9571
rect 25697 9537 25731 9571
rect 26157 9537 26191 9571
rect 27445 9537 27479 9571
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 6009 9469 6043 9503
rect 6929 9469 6963 9503
rect 7205 9469 7239 9503
rect 9137 9469 9171 9503
rect 12265 9469 12299 9503
rect 14473 9469 14507 9503
rect 16221 9469 16255 9503
rect 16957 9469 16991 9503
rect 18429 9469 18463 9503
rect 19165 9469 19199 9503
rect 19441 9469 19475 9503
rect 23305 9469 23339 9503
rect 23489 9469 23523 9503
rect 24409 9469 24443 9503
rect 24593 9469 24627 9503
rect 1777 9401 1811 9435
rect 17509 9401 17543 9435
rect 3065 9333 3099 9367
rect 3709 9333 3743 9367
rect 20269 9333 20303 9367
rect 24869 9333 24903 9367
rect 25513 9333 25547 9367
rect 26249 9333 26283 9367
rect 5733 9129 5767 9163
rect 9413 9129 9447 9163
rect 11424 9129 11458 9163
rect 16129 9129 16163 9163
rect 18705 9129 18739 9163
rect 19441 9129 19475 9163
rect 20085 9129 20119 9163
rect 22017 9129 22051 9163
rect 22661 9129 22695 9163
rect 25237 9129 25271 9163
rect 18061 9061 18095 9095
rect 7113 8993 7147 9027
rect 11161 8993 11195 9027
rect 14657 8993 14691 9027
rect 21557 8993 21591 9027
rect 1961 8925 1995 8959
rect 2605 8925 2639 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 6193 8925 6227 8959
rect 6837 8925 6871 8959
rect 9597 8925 9631 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 13737 8925 13771 8959
rect 14381 8925 14415 8959
rect 16589 8925 16623 8959
rect 16773 8925 16807 8959
rect 18245 8925 18279 8959
rect 18889 8925 18923 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20729 8925 20763 8959
rect 21373 8925 21407 8959
rect 22845 8925 22879 8959
rect 23305 8925 23339 8959
rect 24593 8925 24627 8959
rect 25421 8925 25455 8959
rect 38025 8925 38059 8959
rect 4261 8857 4295 8891
rect 10701 8857 10735 8891
rect 23397 8857 23431 8891
rect 2053 8789 2087 8823
rect 2697 8789 2731 8823
rect 3341 8789 3375 8823
rect 6285 8789 6319 8823
rect 8585 8789 8619 8823
rect 12909 8789 12943 8823
rect 13553 8789 13587 8823
rect 17233 8789 17267 8823
rect 20821 8789 20855 8823
rect 24685 8789 24719 8823
rect 38209 8789 38243 8823
rect 1777 8585 1811 8619
rect 16129 8585 16163 8619
rect 19257 8585 19291 8619
rect 23213 8585 23247 8619
rect 23673 8585 23707 8619
rect 24317 8585 24351 8619
rect 25053 8585 25087 8619
rect 33701 8585 33735 8619
rect 9321 8517 9355 8551
rect 12725 8517 12759 8551
rect 12817 8517 12851 8551
rect 13369 8517 13403 8551
rect 18245 8517 18279 8551
rect 18797 8517 18831 8551
rect 1685 8449 1719 8483
rect 2513 8449 2547 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 11989 8449 12023 8483
rect 12081 8449 12115 8483
rect 16313 8449 16347 8483
rect 16957 8449 16991 8483
rect 19441 8449 19475 8483
rect 19993 8449 20027 8483
rect 21189 8449 21223 8483
rect 24501 8449 24535 8483
rect 24961 8449 24995 8483
rect 33609 8449 33643 8483
rect 2973 8381 3007 8415
rect 3249 8381 3283 8415
rect 5273 8381 5307 8415
rect 7113 8381 7147 8415
rect 7389 8381 7423 8415
rect 8861 8381 8895 8415
rect 13829 8381 13863 8415
rect 14105 8381 14139 8415
rect 17141 8381 17175 8415
rect 18153 8381 18187 8415
rect 21281 8381 21315 8415
rect 22569 8381 22603 8415
rect 22753 8381 22787 8415
rect 2329 8313 2363 8347
rect 4721 8313 4755 8347
rect 5917 8313 5951 8347
rect 10609 8313 10643 8347
rect 17325 8313 17359 8347
rect 15577 8245 15611 8279
rect 20085 8245 20119 8279
rect 9781 8041 9815 8075
rect 10333 8041 10367 8075
rect 16037 8041 16071 8075
rect 21281 8041 21315 8075
rect 21833 8041 21867 8075
rect 23857 8041 23891 8075
rect 38117 8041 38151 8075
rect 8125 7973 8159 8007
rect 23121 7973 23155 8007
rect 4261 7905 4295 7939
rect 10977 7905 11011 7939
rect 16957 7905 16991 7939
rect 18061 7905 18095 7939
rect 20821 7905 20855 7939
rect 6285 7837 6319 7871
rect 9689 7837 9723 7871
rect 10517 7837 10551 7871
rect 13001 7837 13035 7871
rect 13553 7837 13587 7871
rect 14289 7837 14323 7871
rect 18245 7837 18279 7871
rect 20637 7837 20671 7871
rect 21741 7837 21775 7871
rect 22385 7837 22419 7871
rect 23305 7837 23339 7871
rect 23765 7837 23799 7871
rect 24593 7837 24627 7871
rect 38301 7837 38335 7871
rect 1685 7769 1719 7803
rect 3433 7769 3467 7803
rect 4537 7769 4571 7803
rect 6837 7769 6871 7803
rect 11260 7769 11294 7803
rect 14565 7769 14599 7803
rect 17049 7769 17083 7803
rect 17601 7769 17635 7803
rect 19533 7769 19567 7803
rect 19625 7769 19659 7803
rect 20177 7769 20211 7803
rect 22477 7769 22511 7803
rect 13645 7701 13679 7735
rect 18705 7701 18739 7735
rect 24685 7701 24719 7735
rect 2329 7497 2363 7531
rect 2973 7497 3007 7531
rect 8493 7497 8527 7531
rect 13185 7497 13219 7531
rect 20177 7497 20211 7531
rect 28825 7497 28859 7531
rect 7021 7429 7055 7463
rect 9413 7429 9447 7463
rect 10977 7429 11011 7463
rect 14013 7429 14047 7463
rect 17049 7429 17083 7463
rect 17601 7429 17635 7463
rect 1593 7361 1627 7395
rect 2237 7361 2271 7395
rect 2881 7361 2915 7395
rect 3525 7361 3559 7395
rect 4169 7361 4203 7395
rect 6745 7361 6779 7395
rect 11989 7361 12023 7395
rect 13093 7361 13127 7395
rect 13737 7361 13771 7395
rect 18245 7361 18279 7395
rect 18981 7361 19015 7395
rect 20085 7361 20119 7395
rect 20729 7361 20763 7395
rect 22017 7361 22051 7395
rect 22937 7361 22971 7395
rect 23673 7361 23707 7395
rect 28733 7361 28767 7395
rect 4445 7293 4479 7327
rect 5917 7293 5951 7327
rect 12449 7293 12483 7327
rect 15761 7293 15795 7327
rect 16957 7293 16991 7327
rect 19165 7293 19199 7327
rect 23857 7293 23891 7327
rect 1685 7225 1719 7259
rect 11805 7225 11839 7259
rect 18061 7225 18095 7259
rect 19625 7225 19659 7259
rect 22109 7225 22143 7259
rect 23029 7225 23063 7259
rect 3617 7157 3651 7191
rect 20821 7157 20855 7191
rect 24041 7157 24075 7191
rect 7100 6953 7134 6987
rect 10590 6953 10624 6987
rect 13553 6953 13587 6987
rect 15577 6953 15611 6987
rect 28457 6953 28491 6987
rect 17141 6885 17175 6919
rect 33609 6885 33643 6919
rect 5733 6817 5767 6851
rect 8585 6817 8619 6851
rect 10333 6817 10367 6851
rect 12357 6817 12391 6851
rect 16589 6817 16623 6851
rect 17693 6817 17727 6851
rect 18337 6817 18371 6851
rect 19441 6817 19475 6851
rect 3433 6749 3467 6783
rect 3985 6749 4019 6783
rect 6193 6749 6227 6783
rect 6837 6749 6871 6783
rect 9689 6749 9723 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 13737 6749 13771 6783
rect 17877 6749 17911 6783
rect 20545 6749 20579 6783
rect 21189 6749 21223 6783
rect 22017 6749 22051 6783
rect 22661 6749 22695 6783
rect 23121 6749 23155 6783
rect 23949 6749 23983 6783
rect 28365 6749 28399 6783
rect 33517 6749 33551 6783
rect 36461 6749 36495 6783
rect 1685 6681 1719 6715
rect 4261 6681 4295 6715
rect 14289 6681 14323 6715
rect 16681 6681 16715 6715
rect 6285 6613 6319 6647
rect 9781 6613 9815 6647
rect 20637 6613 20671 6647
rect 21281 6613 21315 6647
rect 21833 6613 21867 6647
rect 22477 6613 22511 6647
rect 23213 6613 23247 6647
rect 23765 6613 23799 6647
rect 36553 6613 36587 6647
rect 2605 6409 2639 6443
rect 4629 6409 4663 6443
rect 14289 6409 14323 6443
rect 18613 6409 18647 6443
rect 21373 6409 21407 6443
rect 22661 6409 22695 6443
rect 9229 6341 9263 6375
rect 15761 6341 15795 6375
rect 17141 6341 17175 6375
rect 19257 6341 19291 6375
rect 19809 6341 19843 6375
rect 1593 6273 1627 6307
rect 5181 6273 5215 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 8953 6273 8987 6307
rect 11713 6273 11747 6307
rect 14933 6273 14967 6307
rect 16313 6273 16347 6307
rect 16854 6273 16888 6307
rect 20637 6273 20671 6307
rect 21281 6273 21315 6307
rect 22201 6273 22235 6307
rect 23305 6273 23339 6307
rect 37749 6273 37783 6307
rect 2881 6205 2915 6239
rect 3157 6205 3191 6239
rect 5273 6205 5307 6239
rect 6837 6205 6871 6239
rect 10977 6205 11011 6239
rect 12541 6205 12575 6239
rect 12817 6205 12851 6239
rect 15669 6205 15703 6239
rect 19165 6205 19199 6239
rect 22017 6205 22051 6239
rect 37473 6205 37507 6239
rect 1777 6137 1811 6171
rect 11805 6137 11839 6171
rect 5917 6069 5951 6103
rect 8309 6069 8343 6103
rect 15025 6069 15059 6103
rect 20729 6069 20763 6103
rect 23121 6069 23155 6103
rect 3341 5865 3375 5899
rect 7941 5865 7975 5899
rect 11713 5865 11747 5899
rect 12909 5865 12943 5899
rect 18245 5865 18279 5899
rect 18705 5865 18739 5899
rect 21925 5865 21959 5899
rect 23857 5865 23891 5899
rect 5733 5797 5767 5831
rect 16037 5797 16071 5831
rect 20085 5797 20119 5831
rect 3985 5729 4019 5763
rect 4261 5729 4295 5763
rect 6193 5729 6227 5763
rect 9413 5729 9447 5763
rect 14289 5729 14323 5763
rect 16497 5729 16531 5763
rect 22569 5729 22603 5763
rect 1593 5661 1627 5695
rect 8401 5661 8435 5695
rect 9137 5661 9171 5695
rect 11161 5661 11195 5695
rect 11621 5661 11655 5695
rect 12449 5661 12483 5695
rect 13093 5661 13127 5695
rect 13737 5661 13771 5695
rect 18889 5661 18923 5695
rect 19441 5661 19475 5695
rect 19625 5661 19659 5695
rect 20545 5661 20579 5695
rect 21189 5661 21223 5695
rect 21833 5661 21867 5695
rect 22477 5661 22511 5695
rect 23121 5661 23155 5695
rect 23765 5661 23799 5695
rect 30665 5661 30699 5695
rect 1869 5593 1903 5627
rect 6469 5593 6503 5627
rect 14565 5593 14599 5627
rect 16773 5593 16807 5627
rect 23213 5593 23247 5627
rect 8493 5525 8527 5559
rect 12265 5525 12299 5559
rect 13553 5525 13587 5559
rect 20637 5525 20671 5559
rect 21281 5525 21315 5559
rect 30481 5525 30515 5559
rect 6745 5321 6779 5355
rect 9045 5321 9079 5355
rect 9781 5321 9815 5355
rect 11069 5321 11103 5355
rect 11897 5321 11931 5355
rect 15117 5321 15151 5355
rect 16221 5321 16255 5355
rect 19073 5321 19107 5355
rect 19809 5321 19843 5355
rect 20545 5321 20579 5355
rect 24041 5321 24075 5355
rect 24685 5321 24719 5355
rect 3893 5253 3927 5287
rect 7560 5253 7594 5287
rect 12817 5253 12851 5287
rect 13645 5253 13679 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 3617 5185 3651 5219
rect 6653 5185 6687 5219
rect 7297 5185 7331 5219
rect 9689 5185 9723 5219
rect 10333 5185 10367 5219
rect 10977 5185 11011 5219
rect 12733 5183 12767 5217
rect 16129 5185 16163 5219
rect 19257 5185 19291 5219
rect 19717 5185 19751 5219
rect 20453 5185 20487 5219
rect 21281 5185 21315 5219
rect 22017 5183 22051 5217
rect 22661 5185 22695 5219
rect 23305 5185 23339 5219
rect 23949 5185 23983 5219
rect 24593 5185 24627 5219
rect 26525 5185 26559 5219
rect 38025 5185 38059 5219
rect 5641 5117 5675 5151
rect 13369 5117 13403 5151
rect 16865 5117 16899 5151
rect 17141 5117 17175 5151
rect 23397 5117 23431 5151
rect 10425 5049 10459 5083
rect 1777 4981 1811 5015
rect 2513 4981 2547 5015
rect 18613 4981 18647 5015
rect 21097 4981 21131 5015
rect 22109 4981 22143 5015
rect 22753 4981 22787 5015
rect 26341 4981 26375 5015
rect 37841 4981 37875 5015
rect 3341 4777 3375 4811
rect 4721 4777 4755 4811
rect 8493 4777 8527 4811
rect 13277 4777 13311 4811
rect 16037 4777 16071 4811
rect 18521 4777 18555 4811
rect 21097 4777 21131 4811
rect 28273 4777 28307 4811
rect 31953 4777 31987 4811
rect 38117 4777 38151 4811
rect 7849 4709 7883 4743
rect 17233 4709 17267 4743
rect 23765 4709 23799 4743
rect 1869 4641 1903 4675
rect 6101 4641 6135 4675
rect 9321 4641 9355 4675
rect 11529 4641 11563 4675
rect 14289 4641 14323 4675
rect 14565 4641 14599 4675
rect 16681 4641 16715 4675
rect 17877 4641 17911 4675
rect 18061 4641 18095 4675
rect 1593 4573 1627 4607
rect 4169 4573 4203 4607
rect 4629 4573 4663 4607
rect 5181 4573 5215 4607
rect 5457 4573 5491 4607
rect 8401 4573 8435 4607
rect 19993 4573 20027 4607
rect 21281 4573 21315 4607
rect 21833 4573 21867 4607
rect 22477 4573 22511 4607
rect 23121 4573 23155 4607
rect 23949 4573 23983 4607
rect 28181 4573 28215 4607
rect 31861 4573 31895 4607
rect 38301 4573 38335 4607
rect 6377 4505 6411 4539
rect 9597 4505 9631 4539
rect 11805 4505 11839 4539
rect 16773 4505 16807 4539
rect 23213 4505 23247 4539
rect 4261 4437 4295 4471
rect 5641 4437 5675 4471
rect 11069 4437 11103 4471
rect 20085 4437 20119 4471
rect 21925 4437 21959 4471
rect 22569 4437 22603 4471
rect 23857 4233 23891 4267
rect 24593 4233 24627 4267
rect 1593 4165 1627 4199
rect 3801 4097 3835 4131
rect 5825 4097 5859 4131
rect 7941 4097 7975 4131
rect 10333 4097 10367 4131
rect 10977 4097 11011 4131
rect 11069 4097 11103 4131
rect 11805 4097 11839 4131
rect 14013 4097 14047 4131
rect 17141 4097 17175 4131
rect 17969 4097 18003 4131
rect 19165 4097 19199 4131
rect 19625 4097 19659 4131
rect 19717 4097 19751 4131
rect 20269 4097 20303 4131
rect 20361 4097 20395 4131
rect 21281 4097 21315 4131
rect 22293 4097 22327 4131
rect 23213 4097 23247 4131
rect 23305 4097 23339 4131
rect 24041 4097 24075 4131
rect 24501 4097 24535 4131
rect 25145 4097 25179 4131
rect 38301 4097 38335 4131
rect 3341 4029 3375 4063
rect 4077 4029 4111 4063
rect 6561 4029 6595 4063
rect 6837 4029 6871 4063
rect 8217 4029 8251 4063
rect 12081 4029 12115 4063
rect 13553 4029 13587 4063
rect 14289 4029 14323 4063
rect 22569 4029 22603 4063
rect 15761 3961 15795 3995
rect 17233 3961 17267 3995
rect 17785 3961 17819 3995
rect 18981 3961 19015 3995
rect 38117 3961 38151 3995
rect 9689 3893 9723 3927
rect 10425 3893 10459 3927
rect 21373 3893 21407 3927
rect 25237 3893 25271 3927
rect 3341 3689 3375 3723
rect 19625 3689 19659 3723
rect 20269 3689 20303 3723
rect 38117 3689 38151 3723
rect 16037 3621 16071 3655
rect 25237 3621 25271 3655
rect 1869 3553 1903 3587
rect 3985 3553 4019 3587
rect 6469 3553 6503 3587
rect 6745 3553 6779 3587
rect 10425 3553 10459 3587
rect 10701 3553 10735 3587
rect 12449 3553 12483 3587
rect 14289 3553 14323 3587
rect 16589 3553 16623 3587
rect 21557 3553 21591 3587
rect 22477 3553 22511 3587
rect 23397 3553 23431 3587
rect 1593 3485 1627 3519
rect 9321 3485 9355 3519
rect 9781 3485 9815 3519
rect 13461 3485 13495 3519
rect 19533 3485 19567 3519
rect 20177 3485 20211 3519
rect 21281 3485 21315 3519
rect 22293 3485 22327 3519
rect 23213 3485 23247 3519
rect 24593 3485 24627 3519
rect 24685 3485 24719 3519
rect 25421 3485 25455 3519
rect 36093 3485 36127 3519
rect 38301 3485 38335 3519
rect 4261 3417 4295 3451
rect 6009 3417 6043 3451
rect 8493 3417 8527 3451
rect 14565 3417 14599 3451
rect 16865 3417 16899 3451
rect 9137 3349 9171 3383
rect 9873 3349 9907 3383
rect 13645 3349 13679 3383
rect 18337 3349 18371 3383
rect 36185 3349 36219 3383
rect 6837 3145 6871 3179
rect 15761 3145 15795 3179
rect 23121 3145 23155 3179
rect 25789 3145 25823 3179
rect 5549 3077 5583 3111
rect 7205 3077 7239 3111
rect 11805 3077 11839 3111
rect 17141 3077 17175 3111
rect 21281 3077 21315 3111
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 6653 3009 6687 3043
rect 9321 3009 9355 3043
rect 9781 3009 9815 3043
rect 10885 3009 10919 3043
rect 13461 3009 13495 3043
rect 14013 3009 14047 3043
rect 16865 3009 16899 3043
rect 19349 3009 19383 3043
rect 19993 3009 20027 3043
rect 21005 3009 21039 3043
rect 22017 3009 22051 3043
rect 22293 3009 22327 3043
rect 23029 3009 23063 3043
rect 23857 3009 23891 3043
rect 24685 3009 24719 3043
rect 25145 3009 25179 3043
rect 25973 3009 26007 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 3801 2941 3835 2975
rect 7297 2941 7331 2975
rect 7573 2941 7607 2975
rect 14289 2941 14323 2975
rect 23949 2941 23983 2975
rect 19441 2873 19475 2907
rect 24501 2873 24535 2907
rect 2973 2805 3007 2839
rect 9965 2805 9999 2839
rect 11069 2805 11103 2839
rect 18613 2805 18647 2839
rect 20085 2805 20119 2839
rect 25237 2805 25271 2839
rect 36737 2805 36771 2839
rect 38209 2805 38243 2839
rect 13553 2601 13587 2635
rect 16037 2601 16071 2635
rect 18245 2601 18279 2635
rect 18705 2601 18739 2635
rect 20269 2601 20303 2635
rect 27169 2601 27203 2635
rect 29745 2601 29779 2635
rect 30389 2601 30423 2635
rect 33609 2601 33643 2635
rect 3341 2533 3375 2567
rect 8493 2533 8527 2567
rect 34897 2533 34931 2567
rect 1593 2465 1627 2499
rect 3985 2465 4019 2499
rect 4261 2465 4295 2499
rect 6009 2465 6043 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 11161 2465 11195 2499
rect 11805 2465 11839 2499
rect 14289 2465 14323 2499
rect 9413 2397 9447 2431
rect 16865 2397 16899 2431
rect 17601 2397 17635 2431
rect 17785 2397 17819 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20177 2397 20211 2431
rect 20821 2397 20855 2431
rect 22017 2397 22051 2431
rect 22937 2397 22971 2431
rect 23673 2397 23707 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 27353 2397 27387 2431
rect 29929 2397 29963 2431
rect 30573 2397 30607 2431
rect 32321 2397 32355 2431
rect 33793 2397 33827 2431
rect 35081 2397 35115 2431
rect 36185 2397 36219 2431
rect 38025 2397 38059 2431
rect 1869 2329 1903 2363
rect 12081 2329 12115 2363
rect 14565 2329 14599 2363
rect 22293 2329 22327 2363
rect 17049 2261 17083 2295
rect 19625 2261 19659 2295
rect 20913 2261 20947 2295
rect 23121 2261 23155 2295
rect 23765 2261 23799 2295
rect 24777 2261 24811 2295
rect 26065 2261 26099 2295
rect 32505 2261 32539 2295
rect 36369 2261 36403 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 14 37272 20 37324
rect 72 37312 78 37324
rect 72 37284 2912 37312
rect 72 37272 78 37284
rect 1302 37204 1308 37256
rect 1360 37244 1366 37256
rect 1765 37247 1823 37253
rect 1765 37244 1777 37247
rect 1360 37216 1777 37244
rect 1360 37204 1366 37216
rect 1765 37213 1777 37216
rect 1811 37213 1823 37247
rect 1765 37207 1823 37213
rect 2409 37247 2467 37253
rect 2409 37213 2421 37247
rect 2455 37244 2467 37247
rect 2774 37244 2780 37256
rect 2455 37216 2780 37244
rect 2455 37213 2467 37216
rect 2409 37207 2467 37213
rect 2774 37204 2780 37216
rect 2832 37204 2838 37256
rect 2884 37244 2912 37284
rect 34716 37284 35204 37312
rect 3053 37247 3111 37253
rect 3053 37244 3065 37247
rect 2884 37216 3065 37244
rect 3053 37213 3065 37216
rect 3099 37213 3111 37247
rect 3053 37207 3111 37213
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37244 4675 37247
rect 5442 37244 5448 37256
rect 4663 37216 5448 37244
rect 4663 37213 4675 37216
rect 4617 37207 4675 37213
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 6546 37244 6552 37256
rect 6507 37216 6552 37244
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 7834 37244 7840 37256
rect 7795 37216 7840 37244
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9030 37204 9036 37256
rect 9088 37244 9094 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 9088 37216 9321 37244
rect 9088 37204 9094 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 10410 37244 10416 37256
rect 10371 37216 10416 37244
rect 9309 37207 9367 37213
rect 10410 37204 10416 37216
rect 10468 37204 10474 37256
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 12492 37216 12541 37244
rect 12492 37204 12498 37216
rect 12529 37213 12541 37216
rect 12575 37213 12587 37247
rect 14274 37244 14280 37256
rect 14235 37216 14280 37244
rect 12529 37207 12587 37213
rect 14274 37204 14280 37216
rect 14332 37204 14338 37256
rect 15565 37247 15623 37253
rect 15565 37213 15577 37247
rect 15611 37244 15623 37247
rect 15746 37244 15752 37256
rect 15611 37216 15752 37244
rect 15611 37213 15623 37216
rect 15565 37207 15623 37213
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 18325 37207 18383 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21324 37216 22201 37244
rect 21324 37204 21330 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22833 37207 22891 37213
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 26053 37207 26111 37213
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 27985 37247 28043 37253
rect 27985 37244 27997 37247
rect 27764 37216 27997 37244
rect 27764 37204 27770 37216
rect 27985 37213 27997 37216
rect 28031 37213 28043 37247
rect 27985 37207 28043 37213
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29052 37216 29929 37244
rect 29052 37204 29058 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30432 37216 30573 37244
rect 30432 37204 30438 37216
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 30561 37207 30619 37213
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32272 37216 32505 37244
rect 32272 37204 32278 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 33962 37204 33968 37256
rect 34020 37244 34026 37256
rect 34716 37244 34744 37284
rect 34020 37216 34744 37244
rect 34020 37204 34026 37216
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 5350 37176 5356 37188
rect 2240 37148 5356 37176
rect 1578 37108 1584 37120
rect 1539 37080 1584 37108
rect 1578 37068 1584 37080
rect 1636 37068 1642 37120
rect 2240 37117 2268 37148
rect 5350 37136 5356 37148
rect 5408 37136 5414 37188
rect 20346 37136 20352 37188
rect 20404 37176 20410 37188
rect 20404 37148 22692 37176
rect 20404 37136 20410 37148
rect 2225 37111 2283 37117
rect 2225 37077 2237 37111
rect 2271 37077 2283 37111
rect 2866 37108 2872 37120
rect 2827 37080 2872 37108
rect 2225 37071 2283 37077
rect 2866 37068 2872 37080
rect 2924 37068 2930 37120
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4801 37111 4859 37117
rect 4801 37108 4813 37111
rect 4672 37080 4813 37108
rect 4672 37068 4678 37080
rect 4801 37077 4813 37080
rect 4847 37077 4859 37111
rect 4801 37071 4859 37077
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 6733 37111 6791 37117
rect 6733 37108 6745 37111
rect 5868 37080 6745 37108
rect 5868 37068 5874 37080
rect 6733 37077 6745 37080
rect 6779 37077 6791 37111
rect 6733 37071 6791 37077
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 9125 37111 9183 37117
rect 9125 37077 9137 37111
rect 9171 37108 9183 37111
rect 9306 37108 9312 37120
rect 9171 37080 9312 37108
rect 9171 37077 9183 37080
rect 9125 37071 9183 37077
rect 9306 37068 9312 37080
rect 9364 37068 9370 37120
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 12342 37108 12348 37120
rect 12303 37080 12348 37108
rect 10597 37071 10655 37077
rect 12342 37068 12348 37080
rect 12400 37068 12406 37120
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13596 37080 14473 37108
rect 13596 37068 13602 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 17126 37068 17132 37120
rect 17184 37108 17190 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 17184 37080 18153 37108
rect 17184 37068 17190 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 20438 37068 20444 37120
rect 20496 37108 20502 37120
rect 22664 37117 22692 37148
rect 23382 37136 23388 37188
rect 23440 37176 23446 37188
rect 23440 37148 25912 37176
rect 23440 37136 23446 37148
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 20496 37080 22017 37108
rect 20496 37068 20502 37080
rect 22005 37077 22017 37080
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 22649 37111 22707 37117
rect 22649 37077 22661 37111
rect 22695 37077 22707 37111
rect 22649 37071 22707 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 25884 37117 25912 37148
rect 29638 37136 29644 37188
rect 29696 37176 29702 37188
rect 29696 37148 32352 37176
rect 29696 37136 29702 37148
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25869 37111 25927 37117
rect 25869 37077 25881 37111
rect 25915 37077 25927 37111
rect 25869 37071 25927 37077
rect 27614 37068 27620 37120
rect 27672 37108 27678 37120
rect 27801 37111 27859 37117
rect 27801 37108 27813 37111
rect 27672 37080 27813 37108
rect 27672 37068 27678 37080
rect 27801 37077 27813 37080
rect 27847 37077 27859 37111
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 27801 37071 27859 37077
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 32324 37117 32352 37148
rect 32582 37136 32588 37188
rect 32640 37176 32646 37188
rect 35176 37176 35204 37284
rect 36722 37204 36728 37256
rect 36780 37244 36786 37256
rect 36909 37247 36967 37253
rect 36909 37244 36921 37247
rect 36780 37216 36921 37244
rect 36780 37204 36786 37216
rect 36909 37213 36921 37216
rect 36955 37213 36967 37247
rect 36909 37207 36967 37213
rect 38013 37247 38071 37253
rect 38013 37213 38025 37247
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 38028 37176 38056 37207
rect 32640 37148 34928 37176
rect 35176 37148 38056 37176
rect 32640 37136 32646 37148
rect 30377 37111 30435 37117
rect 30377 37108 30389 37111
rect 29880 37080 30389 37108
rect 29880 37068 29886 37080
rect 30377 37077 30389 37080
rect 30423 37077 30435 37111
rect 30377 37071 30435 37077
rect 32309 37111 32367 37117
rect 32309 37077 32321 37111
rect 32355 37077 32367 37111
rect 32309 37071 32367 37077
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 34900 37117 34928 37148
rect 33597 37111 33655 37117
rect 33597 37108 33609 37111
rect 32456 37080 33609 37108
rect 32456 37068 32462 37080
rect 33597 37077 33609 37080
rect 33643 37077 33655 37111
rect 33597 37071 33655 37077
rect 34885 37111 34943 37117
rect 34885 37077 34897 37111
rect 34931 37077 34943 37111
rect 34885 37071 34943 37077
rect 35342 37068 35348 37120
rect 35400 37108 35406 37120
rect 36725 37111 36783 37117
rect 36725 37108 36737 37111
rect 35400 37080 36737 37108
rect 35400 37068 35406 37080
rect 36725 37077 36737 37080
rect 36771 37077 36783 37111
rect 38194 37108 38200 37120
rect 38155 37080 38200 37108
rect 36725 37071 36783 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1578 36864 1584 36916
rect 1636 36904 1642 36916
rect 6454 36904 6460 36916
rect 1636 36876 6460 36904
rect 1636 36864 1642 36876
rect 6454 36864 6460 36876
rect 6512 36864 6518 36916
rect 6546 36864 6552 36916
rect 6604 36904 6610 36916
rect 9125 36907 9183 36913
rect 9125 36904 9137 36907
rect 6604 36876 9137 36904
rect 6604 36864 6610 36876
rect 9125 36873 9137 36876
rect 9171 36873 9183 36907
rect 9125 36867 9183 36873
rect 3970 36796 3976 36848
rect 4028 36836 4034 36848
rect 9398 36836 9404 36848
rect 4028 36808 9404 36836
rect 4028 36796 4034 36808
rect 9398 36796 9404 36808
rect 9456 36796 9462 36848
rect 24854 36796 24860 36848
rect 24912 36836 24918 36848
rect 29730 36836 29736 36848
rect 24912 36808 29736 36836
rect 24912 36796 24918 36808
rect 29730 36796 29736 36808
rect 29788 36796 29794 36848
rect 39298 36836 39304 36848
rect 37660 36808 39304 36836
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 9309 36771 9367 36777
rect 9309 36737 9321 36771
rect 9355 36768 9367 36771
rect 10686 36768 10692 36780
rect 9355 36740 10692 36768
rect 9355 36737 9367 36740
rect 9309 36731 9367 36737
rect 10686 36728 10692 36740
rect 10744 36728 10750 36780
rect 37660 36777 37688 36808
rect 39298 36796 39304 36808
rect 39356 36796 39362 36848
rect 37645 36771 37703 36777
rect 37645 36737 37657 36771
rect 37691 36737 37703 36771
rect 37645 36731 37703 36737
rect 38010 36728 38016 36780
rect 38068 36768 38074 36780
rect 38289 36771 38347 36777
rect 38289 36768 38301 36771
rect 38068 36740 38301 36768
rect 38068 36728 38074 36740
rect 38289 36737 38301 36740
rect 38335 36737 38347 36771
rect 38289 36731 38347 36737
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 2682 36564 2688 36576
rect 1627 36536 2688 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 2682 36524 2688 36536
rect 2740 36524 2746 36576
rect 29270 36524 29276 36576
rect 29328 36564 29334 36576
rect 37461 36567 37519 36573
rect 37461 36564 37473 36567
rect 29328 36536 37473 36564
rect 29328 36524 29334 36536
rect 37461 36533 37473 36536
rect 37507 36533 37519 36567
rect 38102 36564 38108 36576
rect 38063 36536 38108 36564
rect 37461 36527 37519 36533
rect 38102 36524 38108 36536
rect 38160 36524 38166 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 15746 36360 15752 36372
rect 15707 36332 15752 36360
rect 15746 36320 15752 36332
rect 15804 36320 15810 36372
rect 15930 36156 15936 36168
rect 15891 36128 15936 36156
rect 15930 36116 15936 36128
rect 15988 36116 15994 36168
rect 37182 36116 37188 36168
rect 37240 36156 37246 36168
rect 38289 36159 38347 36165
rect 38289 36156 38301 36159
rect 37240 36128 38301 36156
rect 37240 36116 37246 36128
rect 38289 36125 38301 36128
rect 38335 36125 38347 36159
rect 38289 36119 38347 36125
rect 35894 35980 35900 36032
rect 35952 36020 35958 36032
rect 38105 36023 38163 36029
rect 38105 36020 38117 36023
rect 35952 35992 38117 36020
rect 35952 35980 35958 35992
rect 38105 35989 38117 35992
rect 38151 35989 38163 36023
rect 38105 35983 38163 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 10686 35272 10692 35284
rect 10647 35244 10692 35272
rect 10686 35232 10692 35244
rect 10744 35232 10750 35284
rect 10597 35071 10655 35077
rect 10597 35037 10609 35071
rect 10643 35068 10655 35071
rect 12250 35068 12256 35080
rect 10643 35040 12256 35068
rect 10643 35037 10655 35040
rect 10597 35031 10655 35037
rect 12250 35028 12256 35040
rect 12308 35028 12314 35080
rect 33870 35028 33876 35080
rect 33928 35068 33934 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 33928 35040 38025 35068
rect 33928 35028 33934 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 16850 34728 16856 34740
rect 16811 34700 16856 34728
rect 16850 34688 16856 34700
rect 16908 34688 16914 34740
rect 22833 34731 22891 34737
rect 22833 34697 22845 34731
rect 22879 34728 22891 34731
rect 24578 34728 24584 34740
rect 22879 34700 24584 34728
rect 22879 34697 22891 34700
rect 22833 34691 22891 34697
rect 24578 34688 24584 34700
rect 24636 34688 24642 34740
rect 17034 34592 17040 34604
rect 16995 34564 17040 34592
rect 17034 34552 17040 34564
rect 17092 34552 17098 34604
rect 23014 34592 23020 34604
rect 22975 34564 23020 34592
rect 23014 34552 23020 34564
rect 23072 34552 23078 34604
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 5442 34144 5448 34196
rect 5500 34184 5506 34196
rect 7285 34187 7343 34193
rect 7285 34184 7297 34187
rect 5500 34156 7297 34184
rect 5500 34144 5506 34156
rect 7285 34153 7297 34156
rect 7331 34153 7343 34187
rect 7285 34147 7343 34153
rect 10410 34144 10416 34196
rect 10468 34184 10474 34196
rect 13265 34187 13323 34193
rect 13265 34184 13277 34187
rect 10468 34156 13277 34184
rect 10468 34144 10474 34156
rect 13265 34153 13277 34156
rect 13311 34153 13323 34187
rect 14274 34184 14280 34196
rect 14235 34156 14280 34184
rect 13265 34147 13323 34153
rect 14274 34144 14280 34156
rect 14332 34144 14338 34196
rect 7469 33983 7527 33989
rect 7469 33949 7481 33983
rect 7515 33980 7527 33983
rect 8754 33980 8760 33992
rect 7515 33952 8760 33980
rect 7515 33949 7527 33952
rect 7469 33943 7527 33949
rect 8754 33940 8760 33952
rect 8812 33940 8818 33992
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 13464 33912 13492 33943
rect 13630 33940 13636 33992
rect 13688 33980 13694 33992
rect 14461 33983 14519 33989
rect 14461 33980 14473 33983
rect 13688 33952 14473 33980
rect 13688 33940 13694 33952
rect 14461 33949 14473 33952
rect 14507 33949 14519 33983
rect 14461 33943 14519 33949
rect 14550 33912 14556 33924
rect 13464 33884 14556 33912
rect 14550 33872 14556 33884
rect 14608 33872 14614 33924
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 19429 33643 19487 33649
rect 19429 33609 19441 33643
rect 19475 33640 19487 33643
rect 20070 33640 20076 33652
rect 19475 33612 20076 33640
rect 19475 33609 19487 33612
rect 19429 33603 19487 33609
rect 20070 33600 20076 33612
rect 20128 33600 20134 33652
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33504 1639 33507
rect 3418 33504 3424 33516
rect 1627 33476 3424 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 3418 33464 3424 33476
rect 3476 33464 3482 33516
rect 12342 33464 12348 33516
rect 12400 33504 12406 33516
rect 14185 33507 14243 33513
rect 14185 33504 14197 33507
rect 12400 33476 14197 33504
rect 12400 33464 12406 33476
rect 14185 33473 14197 33476
rect 14231 33473 14243 33507
rect 14185 33467 14243 33473
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19484 33476 19625 33504
rect 19484 33464 19490 33476
rect 19613 33473 19625 33476
rect 19659 33473 19671 33507
rect 23382 33504 23388 33516
rect 23343 33476 23388 33504
rect 19613 33467 19671 33473
rect 23382 33464 23388 33476
rect 23440 33464 23446 33516
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 37826 33464 37832 33516
rect 37884 33504 37890 33516
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 37884 33476 38025 33504
rect 37884 33464 37890 33476
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 1762 33368 1768 33380
rect 1723 33340 1768 33368
rect 1762 33328 1768 33340
rect 1820 33328 1826 33380
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 14277 33303 14335 33309
rect 14277 33269 14289 33303
rect 14323 33300 14335 33303
rect 15654 33300 15660 33312
rect 14323 33272 15660 33300
rect 14323 33269 14335 33272
rect 14277 33263 14335 33269
rect 15654 33260 15660 33272
rect 15712 33260 15718 33312
rect 22186 33260 22192 33312
rect 22244 33300 22250 33312
rect 23477 33303 23535 33309
rect 23477 33300 23489 33303
rect 22244 33272 23489 33300
rect 22244 33260 22250 33272
rect 23477 33269 23489 33272
rect 23523 33269 23535 33303
rect 24946 33300 24952 33312
rect 24907 33272 24952 33300
rect 23477 33263 23535 33269
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 7834 33056 7840 33108
rect 7892 33096 7898 33108
rect 9769 33099 9827 33105
rect 9769 33096 9781 33099
rect 7892 33068 9781 33096
rect 7892 33056 7898 33068
rect 9769 33065 9781 33068
rect 9815 33065 9827 33099
rect 9769 33059 9827 33065
rect 32398 33028 32404 33040
rect 28184 33000 32404 33028
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32892 10011 32895
rect 11790 32892 11796 32904
rect 9999 32864 11796 32892
rect 9999 32861 10011 32864
rect 9953 32855 10011 32861
rect 11790 32852 11796 32864
rect 11848 32852 11854 32904
rect 16853 32895 16911 32901
rect 16853 32861 16865 32895
rect 16899 32892 16911 32895
rect 17126 32892 17132 32904
rect 16899 32864 17132 32892
rect 16899 32861 16911 32864
rect 16853 32855 16911 32861
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 28184 32901 28212 33000
rect 32398 32988 32404 33000
rect 32456 32988 32462 33040
rect 35342 32960 35348 32972
rect 31036 32932 35348 32960
rect 31036 32901 31064 32932
rect 35342 32920 35348 32932
rect 35400 32920 35406 32972
rect 28169 32895 28227 32901
rect 28169 32861 28181 32895
rect 28215 32861 28227 32895
rect 28169 32855 28227 32861
rect 31021 32895 31079 32901
rect 31021 32861 31033 32895
rect 31067 32861 31079 32895
rect 31021 32855 31079 32861
rect 31665 32895 31723 32901
rect 31665 32861 31677 32895
rect 31711 32892 31723 32895
rect 38102 32892 38108 32904
rect 31711 32864 38108 32892
rect 31711 32861 31723 32864
rect 31665 32855 31723 32861
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 15102 32716 15108 32768
rect 15160 32756 15166 32768
rect 16945 32759 17003 32765
rect 16945 32756 16957 32759
rect 15160 32728 16957 32756
rect 15160 32716 15166 32728
rect 16945 32725 16957 32728
rect 16991 32725 17003 32759
rect 28258 32756 28264 32768
rect 28219 32728 28264 32756
rect 16945 32719 17003 32725
rect 28258 32716 28264 32728
rect 28316 32716 28322 32768
rect 31110 32756 31116 32768
rect 31071 32728 31116 32756
rect 31110 32716 31116 32728
rect 31168 32716 31174 32768
rect 31757 32759 31815 32765
rect 31757 32725 31769 32759
rect 31803 32756 31815 32759
rect 31846 32756 31852 32768
rect 31803 32728 31852 32756
rect 31803 32725 31815 32728
rect 31757 32719 31815 32725
rect 31846 32716 31852 32728
rect 31904 32716 31910 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 15930 32512 15936 32564
rect 15988 32552 15994 32564
rect 16945 32555 17003 32561
rect 16945 32552 16957 32555
rect 15988 32524 16957 32552
rect 15988 32512 15994 32524
rect 16945 32521 16957 32524
rect 16991 32521 17003 32555
rect 16945 32515 17003 32521
rect 20438 32484 20444 32496
rect 19628 32456 20444 32484
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 5350 32376 5356 32428
rect 5408 32416 5414 32428
rect 7377 32419 7435 32425
rect 7377 32416 7389 32419
rect 5408 32388 7389 32416
rect 5408 32376 5414 32388
rect 7377 32385 7389 32388
rect 7423 32385 7435 32419
rect 7377 32379 7435 32385
rect 16853 32419 16911 32425
rect 16853 32385 16865 32419
rect 16899 32416 16911 32419
rect 16942 32416 16948 32428
rect 16899 32388 16948 32416
rect 16899 32385 16911 32388
rect 16853 32379 16911 32385
rect 16942 32376 16948 32388
rect 17000 32376 17006 32428
rect 19628 32425 19656 32456
rect 20438 32444 20444 32456
rect 20496 32444 20502 32496
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 20346 32416 20352 32428
rect 20307 32388 20352 32416
rect 19613 32379 19671 32385
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 38286 32416 38292 32428
rect 38247 32388 38292 32416
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 6730 32212 6736 32224
rect 1627 32184 6736 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 6730 32172 6736 32184
rect 6788 32172 6794 32224
rect 7466 32212 7472 32224
rect 7427 32184 7472 32212
rect 7466 32172 7472 32184
rect 7524 32172 7530 32224
rect 18046 32172 18052 32224
rect 18104 32212 18110 32224
rect 19705 32215 19763 32221
rect 19705 32212 19717 32215
rect 18104 32184 19717 32212
rect 18104 32172 18110 32184
rect 19705 32181 19717 32184
rect 19751 32181 19763 32215
rect 20438 32212 20444 32224
rect 20399 32184 20444 32212
rect 19705 32175 19763 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 33226 32172 33232 32224
rect 33284 32212 33290 32224
rect 38105 32215 38163 32221
rect 38105 32212 38117 32215
rect 33284 32184 38117 32212
rect 33284 32172 33290 32184
rect 38105 32181 38117 32184
rect 38151 32181 38163 32215
rect 38105 32175 38163 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 33873 32011 33931 32017
rect 33873 31977 33885 32011
rect 33919 32008 33931 32011
rect 33962 32008 33968 32020
rect 33919 31980 33968 32008
rect 33919 31977 33931 31980
rect 33873 31971 33931 31977
rect 33962 31968 33968 31980
rect 34020 31968 34026 32020
rect 35894 31872 35900 31884
rect 32140 31844 35900 31872
rect 12250 31764 12256 31816
rect 12308 31804 12314 31816
rect 12802 31804 12808 31816
rect 12308 31776 12808 31804
rect 12308 31764 12314 31776
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 28994 31764 29000 31816
rect 29052 31804 29058 31816
rect 32140 31813 32168 31844
rect 35894 31832 35900 31844
rect 35952 31832 35958 31884
rect 32125 31807 32183 31813
rect 29052 31776 32076 31804
rect 29052 31764 29058 31776
rect 32048 31736 32076 31776
rect 32125 31773 32137 31807
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32214 31764 32220 31816
rect 32272 31804 32278 31816
rect 34057 31807 34115 31813
rect 34057 31804 34069 31807
rect 32272 31776 32317 31804
rect 32416 31776 34069 31804
rect 32272 31764 32278 31776
rect 32416 31736 32444 31776
rect 34057 31773 34069 31776
rect 34103 31773 34115 31807
rect 34057 31767 34115 31773
rect 32048 31708 32444 31736
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 27614 30920 27620 30932
rect 25700 30892 27620 30920
rect 1581 30855 1639 30861
rect 1581 30821 1593 30855
rect 1627 30852 1639 30855
rect 5534 30852 5540 30864
rect 1627 30824 5540 30852
rect 1627 30821 1639 30824
rect 1581 30815 1639 30821
rect 5534 30812 5540 30824
rect 5592 30812 5598 30864
rect 9401 30855 9459 30861
rect 9401 30821 9413 30855
rect 9447 30852 9459 30855
rect 11330 30852 11336 30864
rect 9447 30824 11336 30852
rect 9447 30821 9459 30824
rect 9401 30815 9459 30821
rect 11330 30812 11336 30824
rect 11388 30812 11394 30864
rect 19242 30812 19248 30864
rect 19300 30852 19306 30864
rect 25041 30855 25099 30861
rect 25041 30852 25053 30855
rect 19300 30824 25053 30852
rect 19300 30812 19306 30824
rect 25041 30821 25053 30824
rect 25087 30821 25099 30855
rect 25041 30815 25099 30821
rect 25700 30784 25728 30892
rect 27614 30880 27620 30892
rect 27672 30880 27678 30932
rect 33870 30920 33876 30932
rect 33831 30892 33876 30920
rect 33870 30880 33876 30892
rect 33928 30880 33934 30932
rect 29822 30852 29828 30864
rect 23492 30756 25728 30784
rect 25792 30824 29828 30852
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 2682 30676 2688 30728
rect 2740 30716 2746 30728
rect 5997 30719 6055 30725
rect 5997 30716 6009 30719
rect 2740 30688 6009 30716
rect 2740 30676 2746 30688
rect 5997 30685 6009 30688
rect 6043 30685 6055 30719
rect 9306 30716 9312 30728
rect 9267 30688 9312 30716
rect 5997 30679 6055 30685
rect 9306 30676 9312 30688
rect 9364 30676 9370 30728
rect 9398 30676 9404 30728
rect 9456 30716 9462 30728
rect 23492 30725 23520 30756
rect 9953 30719 10011 30725
rect 9953 30716 9965 30719
rect 9456 30688 9965 30716
rect 9456 30676 9462 30688
rect 9953 30685 9965 30688
rect 9999 30685 10011 30719
rect 9953 30679 10011 30685
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30685 23535 30719
rect 23477 30679 23535 30685
rect 24949 30719 25007 30725
rect 24949 30685 24961 30719
rect 24995 30716 25007 30719
rect 25792 30716 25820 30824
rect 29822 30812 29828 30824
rect 29880 30812 29886 30864
rect 32582 30784 32588 30796
rect 27724 30756 32588 30784
rect 27724 30725 27752 30756
rect 32582 30744 32588 30756
rect 32640 30744 32646 30796
rect 24995 30688 25820 30716
rect 25869 30719 25927 30725
rect 24995 30685 25007 30688
rect 24949 30679 25007 30685
rect 25869 30685 25881 30719
rect 25915 30685 25927 30719
rect 25869 30679 25927 30685
rect 27709 30719 27767 30725
rect 27709 30685 27721 30719
rect 27755 30685 27767 30719
rect 27709 30679 27767 30685
rect 25884 30648 25912 30679
rect 31754 30676 31760 30728
rect 31812 30716 31818 30728
rect 34057 30719 34115 30725
rect 34057 30716 34069 30719
rect 31812 30688 34069 30716
rect 31812 30676 31818 30688
rect 34057 30685 34069 30688
rect 34103 30685 34115 30719
rect 34057 30679 34115 30685
rect 29638 30648 29644 30660
rect 25884 30620 29644 30648
rect 29638 30608 29644 30620
rect 29696 30608 29702 30660
rect 6086 30580 6092 30592
rect 6047 30552 6092 30580
rect 6086 30540 6092 30552
rect 6144 30540 6150 30592
rect 10045 30583 10103 30589
rect 10045 30549 10057 30583
rect 10091 30580 10103 30583
rect 11974 30580 11980 30592
rect 10091 30552 11980 30580
rect 10091 30549 10103 30552
rect 10045 30543 10103 30549
rect 11974 30540 11980 30552
rect 12032 30540 12038 30592
rect 19978 30540 19984 30592
rect 20036 30580 20042 30592
rect 23569 30583 23627 30589
rect 23569 30580 23581 30583
rect 20036 30552 23581 30580
rect 20036 30540 20042 30552
rect 23569 30549 23581 30552
rect 23615 30549 23627 30583
rect 25958 30580 25964 30592
rect 25919 30552 25964 30580
rect 23569 30543 23627 30549
rect 25958 30540 25964 30552
rect 26016 30540 26022 30592
rect 27798 30580 27804 30592
rect 27759 30552 27804 30580
rect 27798 30540 27804 30552
rect 27856 30540 27862 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 6454 30200 6460 30252
rect 6512 30240 6518 30252
rect 8113 30243 8171 30249
rect 8113 30240 8125 30243
rect 6512 30212 8125 30240
rect 6512 30200 6518 30212
rect 8113 30209 8125 30212
rect 8159 30209 8171 30243
rect 29270 30240 29276 30252
rect 29231 30212 29276 30240
rect 8113 30203 8171 30209
rect 29270 30200 29276 30212
rect 29328 30200 29334 30252
rect 38286 30240 38292 30252
rect 38247 30212 38292 30240
rect 38286 30200 38292 30212
rect 38344 30200 38350 30252
rect 8205 30039 8263 30045
rect 8205 30005 8217 30039
rect 8251 30036 8263 30039
rect 11606 30036 11612 30048
rect 8251 30008 11612 30036
rect 8251 30005 8263 30008
rect 8205 29999 8263 30005
rect 11606 29996 11612 30008
rect 11664 29996 11670 30048
rect 29362 30036 29368 30048
rect 29323 30008 29368 30036
rect 29362 29996 29368 30008
rect 29420 29996 29426 30048
rect 36538 29996 36544 30048
rect 36596 30036 36602 30048
rect 38105 30039 38163 30045
rect 38105 30036 38117 30039
rect 36596 30008 38117 30036
rect 36596 29996 36602 30008
rect 38105 30005 38117 30008
rect 38151 30005 38163 30039
rect 38105 29999 38163 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 1627 29260 2774 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 2746 29220 2774 29260
rect 3418 29248 3424 29300
rect 3476 29288 3482 29300
rect 5261 29291 5319 29297
rect 5261 29288 5273 29291
rect 3476 29260 5273 29288
rect 3476 29248 3482 29260
rect 5261 29257 5273 29260
rect 5307 29257 5319 29291
rect 5261 29251 5319 29257
rect 22649 29291 22707 29297
rect 22649 29257 22661 29291
rect 22695 29288 22707 29291
rect 23014 29288 23020 29300
rect 22695 29260 23020 29288
rect 22695 29257 22707 29260
rect 22649 29251 22707 29257
rect 23014 29248 23020 29260
rect 23072 29248 23078 29300
rect 9306 29220 9312 29232
rect 2746 29192 9312 29220
rect 9306 29180 9312 29192
rect 9364 29180 9370 29232
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 5445 29155 5503 29161
rect 5445 29121 5457 29155
rect 5491 29152 5503 29155
rect 10134 29152 10140 29164
rect 5491 29124 10140 29152
rect 5491 29121 5503 29124
rect 5445 29115 5503 29121
rect 10134 29112 10140 29124
rect 10192 29112 10198 29164
rect 11701 29155 11759 29161
rect 11701 29121 11713 29155
rect 11747 29121 11759 29155
rect 22554 29152 22560 29164
rect 22515 29124 22560 29152
rect 11701 29115 11759 29121
rect 2866 29044 2872 29096
rect 2924 29084 2930 29096
rect 11716 29084 11744 29115
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 2924 29056 11744 29084
rect 2924 29044 2930 29056
rect 11793 29019 11851 29025
rect 11793 28985 11805 29019
rect 11839 29016 11851 29019
rect 16850 29016 16856 29028
rect 11839 28988 16856 29016
rect 11839 28985 11851 28988
rect 11793 28979 11851 28985
rect 16850 28976 16856 28988
rect 16908 28976 16914 29028
rect 38102 29016 38108 29028
rect 38063 28988 38108 29016
rect 38102 28976 38108 28988
rect 38160 28976 38166 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 14550 28704 14556 28756
rect 14608 28744 14614 28756
rect 15565 28747 15623 28753
rect 15565 28744 15577 28747
rect 14608 28716 15577 28744
rect 14608 28704 14614 28716
rect 15565 28713 15577 28716
rect 15611 28713 15623 28747
rect 15565 28707 15623 28713
rect 16853 28747 16911 28753
rect 16853 28713 16865 28747
rect 16899 28744 16911 28747
rect 17034 28744 17040 28756
rect 16899 28716 17040 28744
rect 16899 28713 16911 28716
rect 16853 28707 16911 28713
rect 17034 28704 17040 28716
rect 17092 28704 17098 28756
rect 15473 28543 15531 28549
rect 15473 28509 15485 28543
rect 15519 28509 15531 28543
rect 16758 28540 16764 28552
rect 16719 28512 16764 28540
rect 15473 28503 15531 28509
rect 15488 28472 15516 28503
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 17402 28472 17408 28484
rect 15488 28444 17408 28472
rect 17402 28432 17408 28444
rect 17460 28432 17466 28484
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 8754 28200 8760 28212
rect 8715 28172 8760 28200
rect 8754 28160 8760 28172
rect 8812 28160 8818 28212
rect 11790 28200 11796 28212
rect 11751 28172 11796 28200
rect 11790 28160 11796 28172
rect 11848 28160 11854 28212
rect 13630 28200 13636 28212
rect 13591 28172 13636 28200
rect 13630 28160 13636 28172
rect 13688 28160 13694 28212
rect 28994 28200 29000 28212
rect 28955 28172 29000 28200
rect 28994 28160 29000 28172
rect 29052 28160 29058 28212
rect 8665 28067 8723 28073
rect 8665 28033 8677 28067
rect 8711 28064 8723 28067
rect 11054 28064 11060 28076
rect 8711 28036 11060 28064
rect 8711 28033 8723 28036
rect 8665 28027 8723 28033
rect 11054 28024 11060 28036
rect 11112 28024 11118 28076
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28064 11759 28067
rect 12710 28064 12716 28076
rect 11747 28036 12716 28064
rect 11747 28033 11759 28036
rect 11701 28027 11759 28033
rect 12710 28024 12716 28036
rect 12768 28024 12774 28076
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28064 13599 28067
rect 13814 28064 13820 28076
rect 13587 28036 13820 28064
rect 13587 28033 13599 28036
rect 13541 28027 13599 28033
rect 13814 28024 13820 28036
rect 13872 28024 13878 28076
rect 28902 28064 28908 28076
rect 28863 28036 28908 28064
rect 28902 28024 28908 28036
rect 28960 28024 28966 28076
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 19521 27591 19579 27597
rect 19521 27588 19533 27591
rect 19484 27560 19533 27588
rect 19484 27548 19490 27560
rect 19521 27557 19533 27560
rect 19567 27557 19579 27591
rect 19521 27551 19579 27557
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27452 1639 27455
rect 3970 27452 3976 27464
rect 1627 27424 3976 27452
rect 1627 27421 1639 27424
rect 1581 27415 1639 27421
rect 3970 27412 3976 27424
rect 4028 27412 4034 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27452 19487 27455
rect 20070 27452 20076 27464
rect 19475 27424 20076 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 20070 27412 20076 27424
rect 20128 27412 20134 27464
rect 33226 27452 33232 27464
rect 33187 27424 33232 27452
rect 33226 27412 33232 27424
rect 33284 27412 33290 27464
rect 33502 27412 33508 27464
rect 33560 27452 33566 27464
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 33560 27424 38025 27452
rect 33560 27412 33566 27424
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 33318 27316 33324 27328
rect 33279 27288 33324 27316
rect 33318 27276 33324 27288
rect 33376 27276 33382 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 28077 27115 28135 27121
rect 28077 27081 28089 27115
rect 28123 27112 28135 27115
rect 31754 27112 31760 27124
rect 28123 27084 31760 27112
rect 28123 27081 28135 27084
rect 28077 27075 28135 27081
rect 31754 27072 31760 27084
rect 31812 27072 31818 27124
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 6788 26948 8033 26976
rect 6788 26936 6794 26948
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 27985 26979 28043 26985
rect 27985 26976 27997 26979
rect 24820 26948 27997 26976
rect 24820 26936 24826 26948
rect 27985 26945 27997 26948
rect 28031 26945 28043 26979
rect 27985 26939 28043 26945
rect 8113 26775 8171 26781
rect 8113 26741 8125 26775
rect 8159 26772 8171 26775
rect 8938 26772 8944 26784
rect 8159 26744 8944 26772
rect 8159 26741 8171 26744
rect 8113 26735 8171 26741
rect 8938 26732 8944 26744
rect 8996 26732 9002 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 5534 25848 5540 25900
rect 5592 25888 5598 25900
rect 7653 25891 7711 25897
rect 7653 25888 7665 25891
rect 5592 25860 7665 25888
rect 5592 25848 5598 25860
rect 7653 25857 7665 25860
rect 7699 25857 7711 25891
rect 7653 25851 7711 25857
rect 15562 25848 15568 25900
rect 15620 25888 15626 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 15620 25860 17601 25888
rect 15620 25848 15626 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18509 25891 18567 25897
rect 18509 25888 18521 25891
rect 18012 25860 18521 25888
rect 18012 25848 18018 25860
rect 18509 25857 18521 25860
rect 18555 25857 18567 25891
rect 18509 25851 18567 25857
rect 7745 25687 7803 25693
rect 7745 25653 7757 25687
rect 7791 25684 7803 25687
rect 9582 25684 9588 25696
rect 7791 25656 9588 25684
rect 7791 25653 7803 25656
rect 7745 25647 7803 25653
rect 9582 25644 9588 25656
rect 9640 25644 9646 25696
rect 17678 25684 17684 25696
rect 17639 25656 17684 25684
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 18325 25687 18383 25693
rect 18325 25653 18337 25687
rect 18371 25684 18383 25687
rect 18966 25684 18972 25696
rect 18371 25656 18972 25684
rect 18371 25653 18383 25656
rect 18325 25647 18383 25653
rect 18966 25644 18972 25656
rect 19024 25644 19030 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 10134 25480 10140 25492
rect 10095 25452 10140 25480
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 38102 25412 38108 25424
rect 31680 25384 38108 25412
rect 1762 25276 1768 25288
rect 1723 25248 1768 25276
rect 1762 25236 1768 25248
rect 1820 25236 1826 25288
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 12342 25276 12348 25288
rect 10091 25248 12348 25276
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 12342 25236 12348 25248
rect 12400 25236 12406 25288
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 15841 25279 15899 25285
rect 15841 25276 15853 25279
rect 15344 25248 15853 25276
rect 15344 25236 15350 25248
rect 15841 25245 15853 25248
rect 15887 25245 15899 25279
rect 17586 25276 17592 25288
rect 17547 25248 17592 25276
rect 15841 25239 15899 25245
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 19426 25276 19432 25288
rect 19387 25248 19432 25276
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 31680 25285 31708 25384
rect 38102 25372 38108 25384
rect 38160 25372 38166 25424
rect 36538 25344 36544 25356
rect 35866 25316 36544 25344
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25245 31723 25279
rect 31665 25239 31723 25245
rect 32309 25279 32367 25285
rect 32309 25245 32321 25279
rect 32355 25276 32367 25279
rect 35866 25276 35894 25316
rect 36538 25304 36544 25316
rect 36596 25304 36602 25356
rect 32355 25248 35894 25276
rect 32355 25245 32367 25248
rect 32309 25239 32367 25245
rect 36906 25236 36912 25288
rect 36964 25276 36970 25288
rect 38013 25279 38071 25285
rect 38013 25276 38025 25279
rect 36964 25248 38025 25276
rect 36964 25236 36970 25248
rect 38013 25245 38025 25248
rect 38059 25245 38071 25279
rect 38013 25239 38071 25245
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 4062 25140 4068 25152
rect 1627 25112 4068 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 4062 25100 4068 25112
rect 4120 25100 4126 25152
rect 15930 25140 15936 25152
rect 15891 25112 15936 25140
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 17681 25143 17739 25149
rect 17681 25109 17693 25143
rect 17727 25140 17739 25143
rect 18230 25140 18236 25152
rect 17727 25112 18236 25140
rect 17727 25109 17739 25112
rect 17681 25103 17739 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 18598 25140 18604 25152
rect 18559 25112 18604 25140
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 19521 25143 19579 25149
rect 19521 25140 19533 25143
rect 19392 25112 19533 25140
rect 19392 25100 19398 25112
rect 19521 25109 19533 25112
rect 19567 25109 19579 25143
rect 31754 25140 31760 25152
rect 31715 25112 31760 25140
rect 19521 25103 19579 25109
rect 31754 25100 31760 25112
rect 31812 25100 31818 25152
rect 32398 25140 32404 25152
rect 32359 25112 32404 25140
rect 32398 25100 32404 25112
rect 32456 25100 32462 25152
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 18800 24840 19104 24868
rect 6086 24760 6092 24812
rect 6144 24800 6150 24812
rect 9766 24800 9772 24812
rect 6144 24772 9772 24800
rect 6144 24760 6150 24772
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 15470 24800 15476 24812
rect 15431 24772 15476 24800
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 16298 24800 16304 24812
rect 16259 24772 16304 24800
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 17037 24803 17095 24809
rect 17037 24800 17049 24803
rect 16408 24772 17049 24800
rect 15488 24732 15516 24760
rect 16408 24732 16436 24772
rect 17037 24769 17049 24772
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24769 17739 24803
rect 18322 24800 18328 24812
rect 18283 24772 18328 24800
rect 17681 24763 17739 24769
rect 15488 24704 16436 24732
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 17696 24732 17724 24763
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 18800 24800 18828 24840
rect 18966 24800 18972 24812
rect 18708 24772 18828 24800
rect 18927 24772 18972 24800
rect 16632 24704 17724 24732
rect 16632 24692 16638 24704
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18708 24732 18736 24772
rect 18966 24760 18972 24772
rect 19024 24760 19030 24812
rect 19076 24800 19104 24840
rect 20732 24840 21128 24868
rect 20533 24803 20591 24809
rect 20533 24800 20545 24803
rect 19076 24772 20545 24800
rect 20533 24769 20545 24772
rect 20579 24800 20591 24803
rect 20732 24800 20760 24840
rect 20579 24772 20760 24800
rect 20579 24769 20591 24772
rect 20533 24763 20591 24769
rect 20806 24760 20812 24812
rect 20864 24800 20870 24812
rect 20993 24803 21051 24809
rect 20993 24800 21005 24803
rect 20864 24772 21005 24800
rect 20864 24760 20870 24772
rect 20993 24769 21005 24772
rect 21039 24769 21051 24803
rect 21100 24800 21128 24840
rect 22002 24800 22008 24812
rect 21100 24772 22008 24800
rect 20993 24763 21051 24769
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 17828 24704 18736 24732
rect 18785 24735 18843 24741
rect 17828 24692 17834 24704
rect 18785 24701 18797 24735
rect 18831 24732 18843 24735
rect 20622 24732 20628 24744
rect 18831 24704 20628 24732
rect 18831 24701 18843 24704
rect 18785 24695 18843 24701
rect 20622 24692 20628 24704
rect 20680 24732 20686 24744
rect 27798 24732 27804 24744
rect 20680 24704 27804 24732
rect 20680 24692 20686 24704
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 16853 24667 16911 24673
rect 16853 24633 16865 24667
rect 16899 24664 16911 24667
rect 17954 24664 17960 24676
rect 16899 24636 17960 24664
rect 16899 24633 16911 24636
rect 16853 24627 16911 24633
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 18141 24667 18199 24673
rect 18141 24633 18153 24667
rect 18187 24664 18199 24667
rect 19610 24664 19616 24676
rect 18187 24636 19616 24664
rect 18187 24633 18199 24636
rect 18141 24627 18199 24633
rect 19610 24624 19616 24636
rect 19668 24624 19674 24676
rect 15565 24599 15623 24605
rect 15565 24565 15577 24599
rect 15611 24596 15623 24599
rect 15838 24596 15844 24608
rect 15611 24568 15844 24596
rect 15611 24565 15623 24568
rect 15565 24559 15623 24565
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 17494 24596 17500 24608
rect 17455 24568 17500 24596
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 19150 24596 19156 24608
rect 19111 24568 19156 24596
rect 19150 24556 19156 24568
rect 19208 24556 19214 24608
rect 20346 24596 20352 24608
rect 20307 24568 20352 24596
rect 20346 24556 20352 24568
rect 20404 24556 20410 24608
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 15381 24395 15439 24401
rect 15381 24361 15393 24395
rect 15427 24392 15439 24395
rect 16298 24392 16304 24404
rect 15427 24364 16304 24392
rect 15427 24361 15439 24364
rect 15381 24355 15439 24361
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 16669 24395 16727 24401
rect 16669 24361 16681 24395
rect 16715 24392 16727 24395
rect 16758 24392 16764 24404
rect 16715 24364 16764 24392
rect 16715 24361 16727 24364
rect 16669 24355 16727 24361
rect 16758 24352 16764 24364
rect 16816 24352 16822 24404
rect 19150 24392 19156 24404
rect 17052 24364 19156 24392
rect 15930 24216 15936 24268
rect 15988 24256 15994 24268
rect 16209 24259 16267 24265
rect 16209 24256 16221 24259
rect 15988 24228 16221 24256
rect 15988 24216 15994 24228
rect 16209 24225 16221 24228
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 6178 24188 6184 24200
rect 1627 24160 6184 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 15562 24188 15568 24200
rect 15523 24160 15568 24188
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24188 16083 24191
rect 16298 24188 16304 24200
rect 16071 24160 16304 24188
rect 16071 24157 16083 24160
rect 16025 24151 16083 24157
rect 16298 24148 16304 24160
rect 16356 24188 16362 24200
rect 17052 24188 17080 24364
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 33502 24392 33508 24404
rect 33463 24364 33508 24392
rect 33502 24352 33508 24364
rect 33560 24352 33566 24404
rect 31110 24324 31116 24336
rect 17144 24296 31116 24324
rect 17144 24265 17172 24296
rect 31110 24284 31116 24296
rect 31168 24284 31174 24336
rect 17129 24259 17187 24265
rect 17129 24225 17141 24259
rect 17175 24225 17187 24259
rect 17129 24219 17187 24225
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 17678 24256 17684 24268
rect 17359 24228 17684 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24256 18291 24259
rect 18598 24256 18604 24268
rect 18279 24228 18604 24256
rect 18279 24225 18291 24228
rect 18233 24219 18291 24225
rect 18598 24216 18604 24228
rect 18656 24216 18662 24268
rect 20346 24216 20352 24268
rect 20404 24256 20410 24268
rect 20404 24228 21864 24256
rect 20404 24216 20410 24228
rect 16356 24160 17080 24188
rect 16356 24148 16362 24160
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 18417 24191 18475 24197
rect 18417 24188 18429 24191
rect 17552 24160 18429 24188
rect 17552 24148 17558 24160
rect 18417 24157 18429 24160
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 21836 24197 21864 24228
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20772 24160 21005 24188
rect 20772 24148 20778 24160
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 20993 24151 21051 24157
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24157 21879 24191
rect 21821 24151 21879 24157
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 33689 24191 33747 24197
rect 33689 24188 33701 24191
rect 30432 24160 33701 24188
rect 30432 24148 30438 24160
rect 33689 24157 33701 24160
rect 33735 24157 33747 24191
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 33689 24151 33747 24157
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 18690 24080 18696 24132
rect 18748 24120 18754 24132
rect 18877 24123 18935 24129
rect 18877 24120 18889 24123
rect 18748 24092 18889 24120
rect 18748 24080 18754 24092
rect 18877 24089 18889 24092
rect 18923 24120 18935 24123
rect 19521 24123 19579 24129
rect 19521 24120 19533 24123
rect 18923 24092 19533 24120
rect 18923 24089 18935 24092
rect 18877 24083 18935 24089
rect 19521 24089 19533 24092
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 19610 24080 19616 24132
rect 19668 24120 19674 24132
rect 20162 24120 20168 24132
rect 19668 24092 19713 24120
rect 20123 24092 20168 24120
rect 19668 24080 19674 24092
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 21085 24123 21143 24129
rect 21085 24089 21097 24123
rect 21131 24120 21143 24123
rect 22370 24120 22376 24132
rect 21131 24092 22376 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 16482 24012 16488 24064
rect 16540 24052 16546 24064
rect 17773 24055 17831 24061
rect 17773 24052 17785 24055
rect 16540 24024 17785 24052
rect 16540 24012 16546 24024
rect 17773 24021 17785 24024
rect 17819 24021 17831 24055
rect 17773 24015 17831 24021
rect 20898 24012 20904 24064
rect 20956 24052 20962 24064
rect 21637 24055 21695 24061
rect 21637 24052 21649 24055
rect 20956 24024 21649 24052
rect 20956 24012 20962 24024
rect 21637 24021 21649 24024
rect 21683 24021 21695 24055
rect 21637 24015 21695 24021
rect 36998 24012 37004 24064
rect 37056 24052 37062 24064
rect 38105 24055 38163 24061
rect 38105 24052 38117 24055
rect 37056 24024 38117 24052
rect 37056 24012 37062 24024
rect 38105 24021 38117 24024
rect 38151 24021 38163 24055
rect 38105 24015 38163 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3970 23848 3976 23860
rect 3931 23820 3976 23848
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 14369 23851 14427 23857
rect 14369 23817 14381 23851
rect 14415 23817 14427 23851
rect 16298 23848 16304 23860
rect 16259 23820 16304 23848
rect 14369 23811 14427 23817
rect 14384 23780 14412 23811
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 20162 23848 20168 23860
rect 19904 23820 20168 23848
rect 19334 23780 19340 23792
rect 14384 23752 15240 23780
rect 19295 23752 19340 23780
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23712 4215 23715
rect 5534 23712 5540 23724
rect 4203 23684 5540 23712
rect 4203 23681 4215 23684
rect 4157 23675 4215 23681
rect 5534 23672 5540 23684
rect 5592 23672 5598 23724
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13998 23712 14004 23724
rect 13679 23684 14004 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 15212 23721 15240 23752
rect 19334 23740 19340 23752
rect 19392 23740 19398 23792
rect 19904 23789 19932 23820
rect 20162 23808 20168 23820
rect 20220 23848 20226 23860
rect 24762 23848 24768 23860
rect 20220 23820 24768 23848
rect 20220 23808 20226 23820
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 19889 23783 19947 23789
rect 19889 23749 19901 23783
rect 19935 23749 19947 23783
rect 20898 23780 20904 23792
rect 20859 23752 20904 23780
rect 19889 23743 19947 23749
rect 20898 23740 20904 23752
rect 20956 23740 20962 23792
rect 21453 23783 21511 23789
rect 21453 23749 21465 23783
rect 21499 23780 21511 23783
rect 22554 23780 22560 23792
rect 21499 23752 22560 23780
rect 21499 23749 21511 23752
rect 21453 23743 21511 23749
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15654 23712 15660 23724
rect 15615 23684 15660 23712
rect 15197 23675 15255 23681
rect 12986 23644 12992 23656
rect 12947 23616 12992 23644
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 14090 23604 14096 23656
rect 14148 23644 14154 23656
rect 14568 23644 14596 23675
rect 15654 23672 15660 23684
rect 15712 23672 15718 23724
rect 15838 23712 15844 23724
rect 15799 23684 15844 23712
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 16172 23684 17049 23712
rect 16172 23672 16178 23684
rect 17037 23681 17049 23684
rect 17083 23681 17095 23715
rect 18046 23712 18052 23724
rect 18007 23684 18052 23712
rect 17037 23675 17095 23681
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 22002 23712 22008 23724
rect 21963 23684 22008 23712
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 15286 23644 15292 23656
rect 14148 23616 15292 23644
rect 14148 23604 14154 23616
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 16022 23604 16028 23656
rect 16080 23644 16086 23656
rect 16080 23616 16804 23644
rect 16080 23604 16086 23616
rect 15013 23579 15071 23585
rect 15013 23545 15025 23579
rect 15059 23576 15071 23579
rect 16666 23576 16672 23588
rect 15059 23548 16672 23576
rect 15059 23545 15071 23548
rect 15013 23539 15071 23545
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 16776 23576 16804 23616
rect 16850 23604 16856 23656
rect 16908 23644 16914 23656
rect 16908 23616 16953 23644
rect 16908 23604 16914 23616
rect 17126 23604 17132 23656
rect 17184 23644 17190 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 17184 23616 18245 23644
rect 17184 23604 17190 23616
rect 18233 23613 18245 23616
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 19245 23647 19303 23653
rect 19245 23613 19257 23647
rect 19291 23613 19303 23647
rect 19245 23607 19303 23613
rect 20809 23647 20867 23653
rect 20809 23613 20821 23647
rect 20855 23644 20867 23647
rect 22649 23647 22707 23653
rect 22649 23644 22661 23647
rect 20855 23616 22661 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 22649 23613 22661 23616
rect 22695 23613 22707 23647
rect 22649 23607 22707 23613
rect 18417 23579 18475 23585
rect 18417 23576 18429 23579
rect 16776 23548 18429 23576
rect 18417 23545 18429 23548
rect 18463 23576 18475 23579
rect 19260 23576 19288 23607
rect 18463 23548 19288 23576
rect 18463 23545 18475 23548
rect 18417 23539 18475 23545
rect 13722 23508 13728 23520
rect 13683 23480 13728 23508
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 15562 23468 15568 23520
rect 15620 23508 15626 23520
rect 16482 23508 16488 23520
rect 15620 23480 16488 23508
rect 15620 23468 15626 23480
rect 16482 23468 16488 23480
rect 16540 23508 16546 23520
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 16540 23480 17233 23508
rect 16540 23468 16546 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 17221 23471 17279 23477
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22152 23480 22197 23508
rect 22152 23468 22158 23480
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 9214 23264 9220 23316
rect 9272 23304 9278 23316
rect 15197 23307 15255 23313
rect 9272 23276 12434 23304
rect 9272 23264 9278 23276
rect 11977 23239 12035 23245
rect 11977 23205 11989 23239
rect 12023 23205 12035 23239
rect 12406 23236 12434 23276
rect 15197 23273 15209 23307
rect 15243 23304 15255 23307
rect 16574 23304 16580 23316
rect 15243 23276 16580 23304
rect 15243 23273 15255 23276
rect 15197 23267 15255 23273
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 16853 23307 16911 23313
rect 16853 23304 16865 23307
rect 16816 23276 16865 23304
rect 16816 23264 16822 23276
rect 16853 23273 16865 23276
rect 16899 23273 16911 23307
rect 18690 23304 18696 23316
rect 18651 23276 18696 23304
rect 16853 23267 16911 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 24946 23304 24952 23316
rect 19904 23276 24952 23304
rect 15933 23239 15991 23245
rect 12406 23208 15424 23236
rect 11977 23199 12035 23205
rect 11992 23168 12020 23199
rect 11992 23140 12434 23168
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23069 12219 23103
rect 12406 23100 12434 23140
rect 12805 23103 12863 23109
rect 12805 23100 12817 23103
rect 12406 23072 12817 23100
rect 12161 23063 12219 23069
rect 12805 23069 12817 23072
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 12176 23032 12204 23063
rect 14458 23060 14464 23112
rect 14516 23100 14522 23112
rect 15396 23109 15424 23208
rect 15933 23205 15945 23239
rect 15979 23236 15991 23239
rect 17126 23236 17132 23248
rect 15979 23208 17132 23236
rect 15979 23205 15991 23208
rect 15933 23199 15991 23205
rect 17126 23196 17132 23208
rect 17184 23196 17190 23248
rect 17862 23196 17868 23248
rect 17920 23236 17926 23248
rect 19426 23236 19432 23248
rect 17920 23208 19432 23236
rect 17920 23196 17926 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 16666 23168 16672 23180
rect 16627 23140 16672 23168
rect 16666 23128 16672 23140
rect 16724 23128 16730 23180
rect 16850 23128 16856 23180
rect 16908 23168 16914 23180
rect 17678 23168 17684 23180
rect 16908 23140 17684 23168
rect 16908 23128 16914 23140
rect 17678 23128 17684 23140
rect 17736 23168 17742 23180
rect 18049 23171 18107 23177
rect 18049 23168 18061 23171
rect 17736 23140 18061 23168
rect 17736 23128 17742 23140
rect 18049 23137 18061 23140
rect 18095 23137 18107 23171
rect 18230 23168 18236 23180
rect 18191 23140 18236 23168
rect 18049 23131 18107 23137
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 19904 23177 19932 23276
rect 24946 23264 24952 23276
rect 25004 23264 25010 23316
rect 21266 23196 21272 23248
rect 21324 23236 21330 23248
rect 22557 23239 22615 23245
rect 22557 23236 22569 23239
rect 21324 23208 22569 23236
rect 21324 23196 21330 23208
rect 22557 23205 22569 23208
rect 22603 23205 22615 23239
rect 22557 23199 22615 23205
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 20073 23171 20131 23177
rect 20073 23137 20085 23171
rect 20119 23168 20131 23171
rect 21082 23168 21088 23180
rect 20119 23140 21088 23168
rect 20119 23137 20131 23140
rect 20073 23131 20131 23137
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 22186 23168 22192 23180
rect 22147 23140 22192 23168
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 22370 23168 22376 23180
rect 22331 23140 22376 23168
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 14553 23103 14611 23109
rect 14553 23100 14565 23103
rect 14516 23072 14565 23100
rect 14516 23060 14522 23072
rect 14553 23069 14565 23072
rect 14599 23069 14611 23103
rect 14553 23063 14611 23069
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 15841 23103 15899 23109
rect 15841 23100 15853 23103
rect 15427 23072 15853 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 15841 23069 15853 23072
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23100 16543 23103
rect 17310 23100 17316 23112
rect 16531 23072 17316 23100
rect 16531 23069 16543 23072
rect 16485 23063 16543 23069
rect 13446 23032 13452 23044
rect 12176 23004 13452 23032
rect 13446 22992 13452 23004
rect 13504 22992 13510 23044
rect 14645 23035 14703 23041
rect 14645 23001 14657 23035
rect 14691 23032 14703 23035
rect 15746 23032 15752 23044
rect 14691 23004 15752 23032
rect 14691 23001 14703 23004
rect 14645 22995 14703 23001
rect 15746 22992 15752 23004
rect 15804 22992 15810 23044
rect 15856 23032 15884 23063
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22554 23100 22560 23112
rect 21775 23072 22560 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 22554 23060 22560 23072
rect 22612 23060 22618 23112
rect 17586 23032 17592 23044
rect 15856 23004 17592 23032
rect 17586 22992 17592 23004
rect 17644 22992 17650 23044
rect 21085 23035 21143 23041
rect 21085 23001 21097 23035
rect 21131 23001 21143 23035
rect 21085 22995 21143 23001
rect 21177 23035 21235 23041
rect 21177 23001 21189 23035
rect 21223 23032 21235 23035
rect 22094 23032 22100 23044
rect 21223 23004 22100 23032
rect 21223 23001 21235 23004
rect 21177 22995 21235 23001
rect 12621 22967 12679 22973
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 13170 22964 13176 22976
rect 12667 22936 13176 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 13541 22967 13599 22973
rect 13541 22933 13553 22967
rect 13587 22964 13599 22967
rect 14274 22964 14280 22976
rect 13587 22936 14280 22964
rect 13587 22933 13599 22936
rect 13541 22927 13599 22933
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 20533 22967 20591 22973
rect 20533 22964 20545 22967
rect 19300 22936 20545 22964
rect 19300 22924 19306 22936
rect 20533 22933 20545 22936
rect 20579 22933 20591 22967
rect 21100 22964 21128 22995
rect 22094 22992 22100 23004
rect 22152 22992 22158 23044
rect 21266 22964 21272 22976
rect 21100 22936 21272 22964
rect 20533 22927 20591 22933
rect 21266 22924 21272 22936
rect 21324 22924 21330 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 5534 22760 5540 22772
rect 5495 22732 5540 22760
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 18322 22760 18328 22772
rect 17267 22732 18328 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 21266 22760 21272 22772
rect 21227 22732 21272 22760
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 32953 22763 33011 22769
rect 32953 22729 32965 22763
rect 32999 22760 33011 22763
rect 36906 22760 36912 22772
rect 32999 22732 36912 22760
rect 32999 22729 33011 22732
rect 32953 22723 33011 22729
rect 36906 22720 36912 22732
rect 36964 22720 36970 22772
rect 10410 22692 10416 22704
rect 5460 22664 10416 22692
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 5460 22633 5488 22664
rect 10410 22652 10416 22664
rect 10468 22652 10474 22704
rect 16758 22652 16764 22704
rect 16816 22692 16822 22704
rect 18049 22695 18107 22701
rect 18049 22692 18061 22695
rect 16816 22664 18061 22692
rect 16816 22652 16822 22664
rect 18049 22661 18061 22664
rect 18095 22661 18107 22695
rect 18049 22655 18107 22661
rect 18601 22695 18659 22701
rect 18601 22661 18613 22695
rect 18647 22692 18659 22695
rect 21358 22692 21364 22704
rect 18647 22664 21364 22692
rect 18647 22661 18659 22664
rect 18601 22655 18659 22661
rect 21358 22652 21364 22664
rect 21416 22652 21422 22704
rect 5445 22627 5503 22633
rect 5445 22593 5457 22627
rect 5491 22593 5503 22627
rect 9306 22624 9312 22636
rect 9267 22596 9312 22624
rect 5445 22587 5503 22593
rect 9306 22584 9312 22596
rect 9364 22584 9370 22636
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 9732 22596 9965 22624
rect 9732 22584 9738 22596
rect 9953 22593 9965 22596
rect 9999 22593 10011 22627
rect 13078 22624 13084 22636
rect 13039 22596 13084 22624
rect 9953 22587 10011 22593
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 13538 22624 13544 22636
rect 13499 22596 13544 22624
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22624 14430 22636
rect 14829 22627 14887 22633
rect 14829 22624 14841 22627
rect 14424 22596 14841 22624
rect 14424 22584 14430 22596
rect 14829 22593 14841 22596
rect 14875 22593 14887 22627
rect 14829 22587 14887 22593
rect 14918 22584 14924 22636
rect 14976 22624 14982 22636
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 14976 22596 15669 22624
rect 14976 22584 14982 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 16298 22624 16304 22636
rect 16259 22596 16304 22624
rect 15657 22587 15715 22593
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 17402 22624 17408 22636
rect 17363 22596 17408 22624
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 21818 22624 21824 22636
rect 19751 22596 21824 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22189 22627 22247 22633
rect 22189 22624 22201 22627
rect 21968 22596 22201 22624
rect 21968 22584 21974 22596
rect 22189 22593 22201 22596
rect 22235 22593 22247 22627
rect 33134 22624 33140 22636
rect 33095 22596 33140 22624
rect 22189 22587 22247 22593
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 10226 22516 10232 22568
rect 10284 22556 10290 22568
rect 10689 22559 10747 22565
rect 10689 22556 10701 22559
rect 10284 22528 10701 22556
rect 10284 22516 10290 22528
rect 10689 22525 10701 22528
rect 10735 22525 10747 22559
rect 10689 22519 10747 22525
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 12894 22556 12900 22568
rect 12299 22528 12900 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 17678 22516 17684 22568
rect 17736 22556 17742 22568
rect 17957 22559 18015 22565
rect 17957 22556 17969 22559
rect 17736 22528 17969 22556
rect 17736 22516 17742 22528
rect 17957 22525 17969 22528
rect 18003 22525 18015 22559
rect 19518 22556 19524 22568
rect 19431 22528 19524 22556
rect 17957 22519 18015 22525
rect 19518 22516 19524 22528
rect 19576 22556 19582 22568
rect 19978 22556 19984 22568
rect 19576 22528 19984 22556
rect 19576 22516 19582 22528
rect 19978 22516 19984 22528
rect 20036 22516 20042 22568
rect 20622 22556 20628 22568
rect 20583 22528 20628 22556
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 20809 22559 20867 22565
rect 20809 22525 20821 22559
rect 20855 22525 20867 22559
rect 20809 22519 20867 22525
rect 9401 22491 9459 22497
rect 9401 22457 9413 22491
rect 9447 22488 9459 22491
rect 10870 22488 10876 22500
rect 9447 22460 10876 22488
rect 9447 22457 9459 22460
rect 9401 22451 9459 22457
rect 10870 22448 10876 22460
rect 10928 22448 10934 22500
rect 14550 22488 14556 22500
rect 12912 22460 14556 22488
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 5534 22420 5540 22432
rect 1627 22392 5540 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 10045 22423 10103 22429
rect 10045 22389 10057 22423
rect 10091 22420 10103 22423
rect 10318 22420 10324 22432
rect 10091 22392 10324 22420
rect 10091 22389 10103 22392
rect 10045 22383 10103 22389
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 12912 22429 12940 22460
rect 14550 22448 14556 22460
rect 14608 22448 14614 22500
rect 14921 22491 14979 22497
rect 14921 22457 14933 22491
rect 14967 22488 14979 22491
rect 16117 22491 16175 22497
rect 14967 22460 16068 22488
rect 14967 22457 14979 22460
rect 14921 22451 14979 22457
rect 12897 22423 12955 22429
rect 12897 22389 12909 22423
rect 12943 22389 12955 22423
rect 12897 22383 12955 22389
rect 13633 22423 13691 22429
rect 13633 22389 13645 22423
rect 13679 22420 13691 22423
rect 13906 22420 13912 22432
rect 13679 22392 13912 22420
rect 13679 22389 13691 22392
rect 13633 22383 13691 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 14182 22420 14188 22432
rect 14143 22392 14188 22420
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 15473 22423 15531 22429
rect 15473 22389 15485 22423
rect 15519 22420 15531 22423
rect 15654 22420 15660 22432
rect 15519 22392 15660 22420
rect 15519 22389 15531 22392
rect 15473 22383 15531 22389
rect 15654 22380 15660 22392
rect 15712 22380 15718 22432
rect 16040 22420 16068 22460
rect 16117 22457 16129 22491
rect 16163 22488 16175 22491
rect 18230 22488 18236 22500
rect 16163 22460 18236 22488
rect 16163 22457 16175 22460
rect 16117 22451 16175 22457
rect 18230 22448 18236 22460
rect 18288 22448 18294 22500
rect 17034 22420 17040 22432
rect 16040 22392 17040 22420
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17402 22380 17408 22432
rect 17460 22420 17466 22432
rect 17770 22420 17776 22432
rect 17460 22392 17776 22420
rect 17460 22380 17466 22392
rect 17770 22380 17776 22392
rect 17828 22380 17834 22432
rect 18414 22380 18420 22432
rect 18472 22420 18478 22432
rect 19242 22420 19248 22432
rect 18472 22392 19248 22420
rect 18472 22380 18478 22392
rect 19242 22380 19248 22392
rect 19300 22420 19306 22432
rect 19889 22423 19947 22429
rect 19889 22420 19901 22423
rect 19300 22392 19901 22420
rect 19300 22380 19306 22392
rect 19889 22389 19901 22392
rect 19935 22389 19947 22423
rect 20640 22420 20668 22516
rect 20824 22488 20852 22519
rect 22005 22491 22063 22497
rect 22005 22488 22017 22491
rect 20824 22460 22017 22488
rect 22005 22457 22017 22460
rect 22051 22457 22063 22491
rect 22005 22451 22063 22457
rect 21634 22420 21640 22432
rect 20640 22392 21640 22420
rect 19889 22383 19947 22389
rect 21634 22380 21640 22392
rect 21692 22380 21698 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 12345 22219 12403 22225
rect 12345 22185 12357 22219
rect 12391 22216 12403 22219
rect 13078 22216 13084 22228
rect 12391 22188 13084 22216
rect 12391 22185 12403 22188
rect 12345 22179 12403 22185
rect 13078 22176 13084 22188
rect 13136 22176 13142 22228
rect 17310 22216 17316 22228
rect 17271 22188 17316 22216
rect 17310 22176 17316 22188
rect 17368 22216 17374 22228
rect 18417 22219 18475 22225
rect 18417 22216 18429 22219
rect 17368 22188 18429 22216
rect 17368 22176 17374 22188
rect 18417 22185 18429 22188
rect 18463 22185 18475 22219
rect 18417 22179 18475 22185
rect 20714 22176 20720 22228
rect 20772 22176 20778 22228
rect 21818 22216 21824 22228
rect 21779 22188 21824 22216
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 10042 22148 10048 22160
rect 9784 22120 10048 22148
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 22012 9367 22015
rect 9674 22012 9680 22024
rect 9355 21984 9680 22012
rect 9355 21981 9367 21984
rect 9309 21975 9367 21981
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 9784 22021 9812 22120
rect 10042 22108 10048 22120
rect 10100 22148 10106 22160
rect 15930 22148 15936 22160
rect 10100 22120 15936 22148
rect 10100 22108 10106 22120
rect 15930 22108 15936 22120
rect 15988 22108 15994 22160
rect 16666 22108 16672 22160
rect 16724 22148 16730 22160
rect 19518 22148 19524 22160
rect 16724 22120 19524 22148
rect 16724 22108 16730 22120
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22080 9919 22083
rect 11790 22080 11796 22092
rect 9907 22052 11796 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12894 22040 12900 22092
rect 12952 22080 12958 22092
rect 13081 22083 13139 22089
rect 13081 22080 13093 22083
rect 12952 22052 13093 22080
rect 12952 22040 12958 22052
rect 13081 22049 13093 22052
rect 13127 22049 13139 22083
rect 13081 22043 13139 22049
rect 13262 22040 13268 22092
rect 13320 22080 13326 22092
rect 14458 22080 14464 22092
rect 13320 22052 14464 22080
rect 13320 22040 13326 22052
rect 14458 22040 14464 22052
rect 14516 22040 14522 22092
rect 15562 22080 15568 22092
rect 15523 22052 15568 22080
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 16960 22089 16988 22120
rect 19518 22108 19524 22120
rect 19576 22108 19582 22160
rect 20732 22148 20760 22176
rect 20640 22120 20760 22148
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22049 17003 22083
rect 18230 22080 18236 22092
rect 18191 22052 18236 22080
rect 16945 22043 17003 22049
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 20640 22080 20668 22120
rect 20180 22052 20668 22080
rect 20717 22083 20775 22089
rect 9769 22015 9827 22021
rect 9769 21981 9781 22015
rect 9815 21981 9827 22015
rect 10597 22015 10655 22021
rect 10597 22012 10609 22015
rect 9769 21975 9827 21981
rect 9876 21984 10609 22012
rect 8478 21904 8484 21956
rect 8536 21944 8542 21956
rect 9876 21944 9904 21984
rect 10597 21981 10609 21984
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 10778 21972 10784 22024
rect 10836 22012 10842 22024
rect 11057 22015 11115 22021
rect 11057 22012 11069 22015
rect 10836 21984 11069 22012
rect 10836 21972 10842 21984
rect 11057 21981 11069 21984
rect 11103 22012 11115 22015
rect 11885 22015 11943 22021
rect 11103 21984 11836 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 11238 21944 11244 21956
rect 8536 21916 9904 21944
rect 10428 21916 11244 21944
rect 8536 21904 8542 21916
rect 9122 21876 9128 21888
rect 9083 21848 9128 21876
rect 9122 21836 9128 21848
rect 9180 21836 9186 21888
rect 10428 21885 10456 21916
rect 11238 21904 11244 21916
rect 11296 21904 11302 21956
rect 11808 21944 11836 21984
rect 11885 21981 11897 22015
rect 11931 22012 11943 22015
rect 12066 22012 12072 22024
rect 11931 21984 12072 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12406 21984 12541 22012
rect 12406 21944 12434 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 14274 22012 14280 22024
rect 14056 21984 14280 22012
rect 14056 21972 14062 21984
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 15378 22012 15384 22024
rect 15059 21984 15384 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 16209 22015 16267 22021
rect 16209 21981 16221 22015
rect 16255 22012 16267 22015
rect 16850 22012 16856 22024
rect 16255 21984 16856 22012
rect 16255 21981 16267 21984
rect 16209 21975 16267 21981
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 17126 22012 17132 22024
rect 17087 21984 17132 22012
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 18046 22012 18052 22024
rect 18007 21984 18052 22012
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 20180 22021 20208 22052
rect 20717 22049 20729 22083
rect 20763 22080 20775 22083
rect 28258 22080 28264 22092
rect 20763 22052 28264 22080
rect 20763 22049 20775 22052
rect 20717 22043 20775 22049
rect 28258 22040 28264 22052
rect 28316 22040 28322 22092
rect 20165 22015 20223 22021
rect 20165 22012 20177 22015
rect 20036 21984 20177 22012
rect 20036 21972 20042 21984
rect 20165 21981 20177 21984
rect 20211 21981 20223 22015
rect 20165 21975 20223 21981
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21508 21984 22017 22012
rect 21508 21972 21514 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 27433 22015 27491 22021
rect 27433 21981 27445 22015
rect 27479 21981 27491 22015
rect 27433 21975 27491 21981
rect 27525 22015 27583 22021
rect 27525 21981 27537 22015
rect 27571 22012 27583 22015
rect 30374 22012 30380 22024
rect 27571 21984 30380 22012
rect 27571 21981 27583 21984
rect 27525 21975 27583 21981
rect 11808 21916 12434 21944
rect 13170 21904 13176 21956
rect 13228 21944 13234 21956
rect 13725 21947 13783 21953
rect 13228 21916 13273 21944
rect 13228 21904 13234 21916
rect 13725 21913 13737 21947
rect 13771 21913 13783 21947
rect 13725 21907 13783 21913
rect 15657 21947 15715 21953
rect 15657 21913 15669 21947
rect 15703 21944 15715 21947
rect 15746 21944 15752 21956
rect 15703 21916 15752 21944
rect 15703 21913 15715 21916
rect 15657 21907 15715 21913
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21845 10471 21879
rect 11146 21876 11152 21888
rect 11107 21848 11152 21876
rect 10413 21839 10471 21845
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11422 21836 11428 21888
rect 11480 21876 11486 21888
rect 11701 21879 11759 21885
rect 11701 21876 11713 21879
rect 11480 21848 11713 21876
rect 11480 21836 11486 21848
rect 11701 21845 11713 21848
rect 11747 21845 11759 21879
rect 11701 21839 11759 21845
rect 12342 21836 12348 21888
rect 12400 21876 12406 21888
rect 13740 21876 13768 21907
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 18138 21944 18144 21956
rect 15988 21916 18144 21944
rect 15988 21904 15994 21916
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 20070 21904 20076 21956
rect 20128 21944 20134 21956
rect 20809 21947 20867 21953
rect 20809 21944 20821 21947
rect 20128 21916 20821 21944
rect 20128 21904 20134 21916
rect 20809 21913 20821 21916
rect 20855 21913 20867 21947
rect 21358 21944 21364 21956
rect 21319 21916 21364 21944
rect 20809 21907 20867 21913
rect 21358 21904 21364 21916
rect 21416 21904 21422 21956
rect 21542 21904 21548 21956
rect 21600 21944 21606 21956
rect 27448 21944 27476 21975
rect 30374 21972 30380 21984
rect 30432 21972 30438 22024
rect 38102 21944 38108 21956
rect 21600 21916 27476 21944
rect 38063 21916 38108 21944
rect 21600 21904 21606 21916
rect 38102 21904 38108 21916
rect 38160 21904 38166 21956
rect 13998 21876 14004 21888
rect 12400 21848 14004 21876
rect 12400 21836 12406 21848
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 14829 21879 14887 21885
rect 14829 21845 14841 21879
rect 14875 21876 14887 21879
rect 16298 21876 16304 21888
rect 14875 21848 16304 21876
rect 14875 21845 14887 21848
rect 14829 21839 14887 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 19981 21879 20039 21885
rect 19981 21845 19993 21879
rect 20027 21876 20039 21879
rect 21910 21876 21916 21888
rect 20027 21848 21916 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 37918 21836 37924 21888
rect 37976 21876 37982 21888
rect 38197 21879 38255 21885
rect 38197 21876 38209 21879
rect 37976 21848 38209 21876
rect 37976 21836 37982 21848
rect 38197 21845 38209 21848
rect 38243 21845 38255 21879
rect 38197 21839 38255 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 8481 21675 8539 21681
rect 8481 21641 8493 21675
rect 8527 21672 8539 21675
rect 13170 21672 13176 21684
rect 8527 21644 10640 21672
rect 8527 21641 8539 21644
rect 8481 21635 8539 21641
rect 7929 21607 7987 21613
rect 7929 21573 7941 21607
rect 7975 21604 7987 21607
rect 7975 21576 10180 21604
rect 7975 21573 7987 21576
rect 7929 21567 7987 21573
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 4120 21508 7849 21536
rect 4120 21496 4126 21508
rect 7837 21505 7849 21508
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21536 8723 21539
rect 9122 21536 9128 21548
rect 8711 21508 9128 21536
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 9306 21536 9312 21548
rect 9267 21508 9312 21536
rect 9306 21496 9312 21508
rect 9364 21496 9370 21548
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 9968 21468 9996 21499
rect 9140 21440 9996 21468
rect 10152 21468 10180 21576
rect 10226 21564 10232 21616
rect 10284 21604 10290 21616
rect 10612 21613 10640 21644
rect 11992 21644 13176 21672
rect 10505 21607 10563 21613
rect 10505 21604 10517 21607
rect 10284 21576 10517 21604
rect 10284 21564 10290 21576
rect 10505 21573 10517 21576
rect 10551 21573 10563 21607
rect 10505 21567 10563 21573
rect 10597 21607 10655 21613
rect 10597 21573 10609 21607
rect 10643 21573 10655 21607
rect 10597 21567 10655 21573
rect 10686 21564 10692 21616
rect 10744 21604 10750 21616
rect 10744 21576 11192 21604
rect 10744 21564 10750 21576
rect 11164 21536 11192 21576
rect 11992 21545 12020 21644
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 14182 21672 14188 21684
rect 13280 21644 14188 21672
rect 13078 21604 13084 21616
rect 12084 21576 13084 21604
rect 11977 21539 12035 21545
rect 11977 21536 11989 21539
rect 11164 21508 11989 21536
rect 11977 21505 11989 21508
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12084 21468 12112 21576
rect 13078 21564 13084 21576
rect 13136 21564 13142 21616
rect 13280 21545 13308 21644
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21641 15531 21675
rect 15473 21635 15531 21641
rect 16117 21675 16175 21681
rect 16117 21641 16129 21675
rect 16163 21672 16175 21675
rect 18046 21672 18052 21684
rect 16163 21644 18052 21672
rect 16163 21641 16175 21644
rect 16117 21635 16175 21641
rect 13906 21604 13912 21616
rect 13867 21576 13912 21604
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 15488 21604 15516 21635
rect 18046 21632 18052 21644
rect 18104 21632 18110 21684
rect 18138 21632 18144 21684
rect 18196 21672 18202 21684
rect 23106 21672 23112 21684
rect 18196 21644 23112 21672
rect 18196 21632 18202 21644
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 16758 21604 16764 21616
rect 15488 21576 16764 21604
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 17034 21604 17040 21616
rect 16995 21576 17040 21604
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 17586 21604 17592 21616
rect 17547 21576 17592 21604
rect 17586 21564 17592 21576
rect 17644 21564 17650 21616
rect 31754 21604 31760 21616
rect 20456 21576 31760 21604
rect 12621 21539 12679 21545
rect 12621 21536 12633 21539
rect 10152 21440 12112 21468
rect 12406 21508 12633 21536
rect 9140 21409 9168 21440
rect 9125 21403 9183 21409
rect 9125 21369 9137 21403
rect 9171 21369 9183 21403
rect 9125 21363 9183 21369
rect 10226 21360 10232 21412
rect 10284 21400 10290 21412
rect 10778 21400 10784 21412
rect 10284 21372 10784 21400
rect 10284 21360 10290 21372
rect 10778 21360 10784 21372
rect 10836 21360 10842 21412
rect 11054 21400 11060 21412
rect 11015 21372 11060 21400
rect 11054 21360 11060 21372
rect 11112 21360 11118 21412
rect 11793 21403 11851 21409
rect 11793 21369 11805 21403
rect 11839 21400 11851 21403
rect 12406 21400 12434 21508
rect 12621 21505 12633 21508
rect 12667 21505 12679 21539
rect 12621 21499 12679 21505
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 15654 21536 15660 21548
rect 15615 21508 15660 21536
rect 13265 21499 13323 21505
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 18782 21536 18788 21548
rect 18743 21508 18788 21536
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 19242 21536 19248 21548
rect 19203 21508 19248 21536
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 20456 21545 20484 21576
rect 31754 21564 31760 21576
rect 31812 21564 31818 21616
rect 20441 21539 20499 21545
rect 20441 21505 20453 21539
rect 20487 21505 20499 21539
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 20441 21499 20499 21505
rect 20548 21508 22201 21536
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 11839 21372 12434 21400
rect 13832 21400 13860 21431
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 14093 21471 14151 21477
rect 14093 21468 14105 21471
rect 14056 21440 14105 21468
rect 14056 21428 14062 21440
rect 14093 21437 14105 21440
rect 14139 21437 14151 21471
rect 16945 21471 17003 21477
rect 14093 21431 14151 21437
rect 15304 21440 16896 21468
rect 15304 21400 15332 21440
rect 13832 21372 15332 21400
rect 11839 21369 11851 21372
rect 11793 21363 11851 21369
rect 4706 21292 4712 21344
rect 4764 21332 4770 21344
rect 9674 21332 9680 21344
rect 4764 21304 9680 21332
rect 4764 21292 4770 21304
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9769 21335 9827 21341
rect 9769 21301 9781 21335
rect 9815 21332 9827 21335
rect 12158 21332 12164 21344
rect 9815 21304 12164 21332
rect 9815 21301 9827 21304
rect 9769 21295 9827 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 13081 21335 13139 21341
rect 12492 21304 12537 21332
rect 12492 21292 12498 21304
rect 13081 21301 13093 21335
rect 13127 21332 13139 21335
rect 16758 21332 16764 21344
rect 13127 21304 16764 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 16868 21332 16896 21440
rect 16945 21437 16957 21471
rect 16991 21468 17003 21471
rect 18414 21468 18420 21480
rect 16991 21440 18420 21468
rect 16991 21437 17003 21440
rect 16945 21431 17003 21437
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 19426 21468 19432 21480
rect 19387 21440 19432 21468
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 18601 21403 18659 21409
rect 18601 21369 18613 21403
rect 18647 21400 18659 21403
rect 20548 21400 20576 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 20625 21471 20683 21477
rect 20625 21437 20637 21471
rect 20671 21437 20683 21471
rect 20625 21431 20683 21437
rect 18647 21372 20576 21400
rect 20640 21400 20668 21431
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20640 21372 22017 21400
rect 18647 21369 18659 21372
rect 18601 21363 18659 21369
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 16868 21304 19625 21332
rect 19613 21301 19625 21304
rect 19659 21332 19671 21335
rect 20809 21335 20867 21341
rect 20809 21332 20821 21335
rect 19659 21304 20821 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 20809 21301 20821 21304
rect 20855 21301 20867 21335
rect 20809 21295 20867 21301
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 22646 21332 22652 21344
rect 20956 21304 22652 21332
rect 20956 21292 20962 21304
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6178 21088 6184 21140
rect 6236 21128 6242 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6236 21100 6929 21128
rect 6236 21088 6242 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 9582 21088 9588 21140
rect 9640 21128 9646 21140
rect 13725 21131 13783 21137
rect 9640 21100 12434 21128
rect 9640 21088 9646 21100
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21029 7803 21063
rect 10686 21060 10692 21072
rect 10647 21032 10692 21060
rect 7745 21023 7803 21029
rect 7760 20992 7788 21023
rect 10686 21020 10692 21032
rect 10744 21020 10750 21072
rect 10505 20995 10563 21001
rect 10505 20992 10517 20995
rect 7760 20964 10517 20992
rect 10505 20961 10517 20964
rect 10551 20961 10563 20995
rect 10505 20955 10563 20961
rect 11146 20952 11152 21004
rect 11204 20992 11210 21004
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 11204 20964 12173 20992
rect 11204 20952 11210 20964
rect 12161 20961 12173 20964
rect 12207 20961 12219 20995
rect 12406 20992 12434 21100
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 13771 21100 16313 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 16301 21097 16313 21100
rect 16347 21097 16359 21131
rect 16301 21091 16359 21097
rect 12621 21063 12679 21069
rect 12621 21029 12633 21063
rect 12667 21060 12679 21063
rect 14734 21060 14740 21072
rect 12667 21032 14740 21060
rect 12667 21029 12679 21032
rect 12621 21023 12679 21029
rect 14734 21020 14740 21032
rect 14792 21020 14798 21072
rect 16316 21060 16344 21091
rect 17034 21088 17040 21140
rect 17092 21128 17098 21140
rect 18322 21128 18328 21140
rect 17092 21100 18328 21128
rect 17092 21088 17098 21100
rect 18322 21088 18328 21100
rect 18380 21088 18386 21140
rect 18785 21131 18843 21137
rect 18785 21097 18797 21131
rect 18831 21128 18843 21131
rect 19426 21128 19432 21140
rect 18831 21100 19432 21128
rect 18831 21097 18843 21100
rect 18785 21091 18843 21097
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 19613 21131 19671 21137
rect 19613 21097 19625 21131
rect 19659 21128 19671 21131
rect 21450 21128 21456 21140
rect 19659 21100 21456 21128
rect 19659 21097 19671 21100
rect 19613 21091 19671 21097
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 21726 21088 21732 21140
rect 21784 21128 21790 21140
rect 21784 21100 25912 21128
rect 21784 21088 21790 21100
rect 19978 21060 19984 21072
rect 16316 21032 19984 21060
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 20990 21020 20996 21072
rect 21048 21060 21054 21072
rect 21085 21063 21143 21069
rect 21085 21060 21097 21063
rect 21048 21032 21097 21060
rect 21048 21020 21054 21032
rect 21085 21029 21097 21032
rect 21131 21029 21143 21063
rect 22465 21063 22523 21069
rect 22465 21060 22477 21063
rect 21085 21023 21143 21029
rect 22066 21032 22477 21060
rect 13081 20995 13139 21001
rect 13081 20992 13093 20995
rect 12406 20964 13093 20992
rect 12161 20955 12219 20961
rect 13081 20961 13093 20964
rect 13127 20961 13139 20995
rect 13081 20955 13139 20961
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 13722 20992 13728 21004
rect 13311 20964 13728 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 14366 20992 14372 21004
rect 14327 20964 14372 20992
rect 14366 20952 14372 20964
rect 14424 20952 14430 21004
rect 14550 20992 14556 21004
rect 14511 20964 14556 20992
rect 14550 20952 14556 20964
rect 14608 20952 14614 21004
rect 17586 20992 17592 21004
rect 17547 20964 17592 20992
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 20806 20992 20812 21004
rect 19812 20964 20812 20992
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20893 7159 20927
rect 7926 20924 7932 20936
rect 7887 20896 7932 20924
rect 7101 20887 7159 20893
rect 7116 20856 7144 20887
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 8435 20896 10333 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 11977 20927 12035 20933
rect 11977 20893 11989 20927
rect 12023 20893 12035 20927
rect 15930 20924 15936 20936
rect 15891 20896 15936 20924
rect 11977 20887 12035 20893
rect 8662 20856 8668 20868
rect 7116 20828 8668 20856
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 9677 20859 9735 20865
rect 9677 20825 9689 20859
rect 9723 20856 9735 20859
rect 11698 20856 11704 20868
rect 9723 20828 11704 20856
rect 9723 20825 9735 20828
rect 9677 20819 9735 20825
rect 11698 20816 11704 20828
rect 11756 20816 11762 20868
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 5810 20788 5816 20800
rect 1627 20760 5816 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 5810 20748 5816 20760
rect 5868 20748 5874 20800
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 11992 20788 12020 20887
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16114 20924 16120 20936
rect 16075 20896 16120 20924
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18564 20896 18705 20924
rect 18564 20884 18570 20896
rect 18693 20893 18705 20896
rect 18739 20924 18751 20927
rect 18782 20924 18788 20936
rect 18739 20896 18788 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 18782 20884 18788 20896
rect 18840 20884 18846 20936
rect 19812 20933 19840 20964
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 22066 20992 22094 21032
rect 22465 21029 22477 21032
rect 22511 21029 22523 21063
rect 22465 21023 22523 21029
rect 20947 20964 22094 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 19797 20887 19855 20893
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21140 20896 22017 20924
rect 21140 20884 21146 20896
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 23106 20924 23112 20936
rect 23019 20896 23112 20924
rect 22649 20887 22707 20893
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 16482 20856 16488 20868
rect 12492 20828 16488 20856
rect 12492 20816 12498 20828
rect 16482 20816 16488 20828
rect 16540 20816 16546 20868
rect 17129 20859 17187 20865
rect 17129 20825 17141 20859
rect 17175 20825 17187 20859
rect 17129 20819 17187 20825
rect 7524 20760 12020 20788
rect 7524 20748 7530 20760
rect 12066 20748 12072 20800
rect 12124 20788 12130 20800
rect 17034 20788 17040 20800
rect 12124 20760 17040 20788
rect 12124 20748 12130 20760
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17145 20788 17173 20819
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 17276 20828 17321 20856
rect 17276 20816 17282 20828
rect 17586 20816 17592 20868
rect 17644 20856 17650 20868
rect 21726 20856 21732 20868
rect 17644 20828 21732 20856
rect 17644 20816 17650 20828
rect 21726 20816 21732 20828
rect 21784 20816 21790 20868
rect 22664 20856 22692 20887
rect 23106 20884 23112 20896
rect 23164 20924 23170 20936
rect 25498 20924 25504 20936
rect 23164 20896 25504 20924
rect 23164 20884 23170 20896
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 25884 20933 25912 21100
rect 25869 20927 25927 20933
rect 25869 20893 25881 20927
rect 25915 20893 25927 20927
rect 25869 20887 25927 20893
rect 33594 20884 33600 20936
rect 33652 20924 33658 20936
rect 38013 20927 38071 20933
rect 38013 20924 38025 20927
rect 33652 20896 38025 20924
rect 33652 20884 33658 20896
rect 38013 20893 38025 20896
rect 38059 20893 38071 20927
rect 38013 20887 38071 20893
rect 21836 20828 22692 20856
rect 19426 20788 19432 20800
rect 17145 20760 19432 20788
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 21836 20797 21864 20828
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20757 21879 20791
rect 21821 20751 21879 20757
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 23201 20791 23259 20797
rect 23201 20788 23213 20791
rect 22152 20760 23213 20788
rect 22152 20748 22158 20760
rect 23201 20757 23213 20760
rect 23247 20757 23259 20791
rect 23201 20751 23259 20757
rect 25961 20791 26019 20797
rect 25961 20757 25973 20791
rect 26007 20788 26019 20791
rect 33134 20788 33140 20800
rect 26007 20760 33140 20788
rect 26007 20757 26019 20760
rect 25961 20751 26019 20757
rect 33134 20748 33140 20760
rect 33192 20748 33198 20800
rect 38194 20788 38200 20800
rect 38155 20760 38200 20788
rect 38194 20748 38200 20760
rect 38252 20748 38258 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 7561 20587 7619 20593
rect 7561 20553 7573 20587
rect 7607 20584 7619 20587
rect 7926 20584 7932 20596
rect 7607 20556 7932 20584
rect 7607 20553 7619 20556
rect 7561 20547 7619 20553
rect 7926 20544 7932 20556
rect 7984 20544 7990 20596
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 14461 20587 14519 20593
rect 11296 20556 13400 20584
rect 11296 20544 11302 20556
rect 10318 20516 10324 20528
rect 10279 20488 10324 20516
rect 10318 20476 10324 20488
rect 10376 20476 10382 20528
rect 10873 20519 10931 20525
rect 10873 20485 10885 20519
rect 10919 20516 10931 20519
rect 11054 20516 11060 20528
rect 10919 20488 11060 20516
rect 10919 20485 10931 20488
rect 10873 20479 10931 20485
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 12158 20516 12164 20528
rect 12119 20488 12164 20516
rect 12158 20476 12164 20488
rect 12216 20476 12222 20528
rect 12250 20476 12256 20528
rect 12308 20516 12314 20528
rect 13372 20525 13400 20556
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 18598 20584 18604 20596
rect 14507 20556 18604 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 18800 20556 20116 20584
rect 13265 20519 13323 20525
rect 13265 20516 13277 20519
rect 12308 20488 13277 20516
rect 12308 20476 12314 20488
rect 13265 20485 13277 20488
rect 13311 20485 13323 20519
rect 13265 20479 13323 20485
rect 13357 20519 13415 20525
rect 13357 20485 13369 20519
rect 13403 20485 13415 20519
rect 13357 20479 13415 20485
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 17037 20519 17095 20525
rect 17037 20516 17049 20519
rect 16540 20488 17049 20516
rect 16540 20476 16546 20488
rect 17037 20485 17049 20488
rect 17083 20485 17095 20519
rect 17037 20479 17095 20485
rect 17310 20476 17316 20528
rect 17368 20516 17374 20528
rect 18800 20516 18828 20556
rect 17368 20488 18828 20516
rect 17368 20476 17374 20488
rect 18874 20476 18880 20528
rect 18932 20516 18938 20528
rect 19978 20516 19984 20528
rect 18932 20488 18977 20516
rect 19939 20488 19984 20516
rect 18932 20476 18938 20488
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 20088 20525 20116 20556
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 20772 20556 22017 20584
rect 20772 20544 20778 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 20073 20519 20131 20525
rect 20073 20485 20085 20519
rect 20119 20485 20131 20519
rect 20073 20479 20131 20485
rect 20625 20519 20683 20525
rect 20625 20485 20637 20519
rect 20671 20516 20683 20519
rect 21266 20516 21272 20528
rect 20671 20488 21272 20516
rect 20671 20485 20683 20488
rect 20625 20479 20683 20485
rect 21266 20476 21272 20488
rect 21324 20516 21330 20528
rect 21542 20516 21548 20528
rect 21324 20488 21548 20516
rect 21324 20476 21330 20488
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 6914 20448 6920 20460
rect 6875 20420 6920 20448
rect 6914 20408 6920 20420
rect 6972 20448 6978 20460
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 6972 20420 7757 20448
rect 6972 20408 6978 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 8220 20380 8248 20411
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 8444 20420 9045 20448
rect 8444 20408 8450 20420
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9674 20448 9680 20460
rect 9635 20420 9680 20448
rect 9033 20411 9091 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15102 20448 15108 20460
rect 15063 20420 15108 20448
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 18049 20411 18107 20417
rect 9306 20380 9312 20392
rect 3384 20352 9312 20380
rect 3384 20340 3390 20352
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10318 20380 10324 20392
rect 10275 20352 10324 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 12069 20383 12127 20389
rect 10468 20352 10732 20380
rect 10468 20340 10474 20352
rect 8849 20315 8907 20321
rect 8849 20281 8861 20315
rect 8895 20312 8907 20315
rect 10594 20312 10600 20324
rect 8895 20284 10600 20312
rect 8895 20281 8907 20284
rect 8849 20275 8907 20281
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 10704 20312 10732 20352
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 12342 20380 12348 20392
rect 12115 20352 12348 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 15286 20380 15292 20392
rect 15247 20352 15292 20380
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 12526 20312 12532 20324
rect 10704 20284 12532 20312
rect 12526 20272 12532 20284
rect 12584 20312 12590 20324
rect 12621 20315 12679 20321
rect 12621 20312 12633 20315
rect 12584 20284 12633 20312
rect 12584 20272 12590 20284
rect 12621 20281 12633 20284
rect 12667 20281 12679 20315
rect 13814 20312 13820 20324
rect 13775 20284 13820 20312
rect 12621 20275 12679 20281
rect 13814 20272 13820 20284
rect 13872 20272 13878 20324
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 16960 20312 16988 20343
rect 17034 20340 17040 20392
rect 17092 20380 17098 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 17092 20352 17233 20380
rect 17092 20340 17098 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 17678 20312 17684 20324
rect 14976 20284 16896 20312
rect 16960 20284 17684 20312
rect 14976 20272 14982 20284
rect 7006 20244 7012 20256
rect 6967 20216 7012 20244
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 8297 20247 8355 20253
rect 8297 20213 8309 20247
rect 8343 20244 8355 20247
rect 9398 20244 9404 20256
rect 8343 20216 9404 20244
rect 8343 20213 8355 20216
rect 8297 20207 8355 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 9493 20247 9551 20253
rect 9493 20213 9505 20247
rect 9539 20244 9551 20247
rect 11514 20244 11520 20256
rect 9539 20216 11520 20244
rect 9539 20213 9551 20216
rect 9493 20207 9551 20213
rect 11514 20204 11520 20216
rect 11572 20204 11578 20256
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 12250 20244 12256 20256
rect 11756 20216 12256 20244
rect 11756 20204 11762 20216
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 15654 20244 15660 20256
rect 12492 20216 15660 20244
rect 12492 20204 12498 20216
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 15746 20204 15752 20256
rect 15804 20244 15810 20256
rect 16868 20244 16896 20284
rect 17678 20272 17684 20284
rect 17736 20272 17742 20324
rect 18064 20244 18092 20411
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20448 22891 20451
rect 23014 20448 23020 20460
rect 22879 20420 23020 20448
rect 22879 20417 22891 20420
rect 22833 20411 22891 20417
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 18785 20383 18843 20389
rect 18785 20349 18797 20383
rect 18831 20380 18843 20383
rect 20990 20380 20996 20392
rect 18831 20352 20996 20380
rect 18831 20349 18843 20352
rect 18785 20343 18843 20349
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 22646 20340 22652 20392
rect 22704 20380 22710 20392
rect 23492 20380 23520 20411
rect 22704 20352 23520 20380
rect 22704 20340 22710 20352
rect 19334 20312 19340 20324
rect 19295 20284 19340 20312
rect 19334 20272 19340 20284
rect 19392 20312 19398 20324
rect 20162 20312 20168 20324
rect 19392 20284 20168 20312
rect 19392 20272 19398 20284
rect 20162 20272 20168 20284
rect 20220 20272 20226 20324
rect 15804 20216 15849 20244
rect 16868 20216 18092 20244
rect 18141 20247 18199 20253
rect 15804 20204 15810 20216
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 20070 20244 20076 20256
rect 18187 20216 20076 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20898 20204 20904 20256
rect 20956 20244 20962 20256
rect 21177 20247 21235 20253
rect 21177 20244 21189 20247
rect 20956 20216 21189 20244
rect 20956 20204 20962 20216
rect 21177 20213 21189 20216
rect 21223 20213 21235 20247
rect 21177 20207 21235 20213
rect 22649 20247 22707 20253
rect 22649 20213 22661 20247
rect 22695 20244 22707 20247
rect 23198 20244 23204 20256
rect 22695 20216 23204 20244
rect 22695 20213 22707 20216
rect 22649 20207 22707 20213
rect 23198 20204 23204 20216
rect 23256 20204 23262 20256
rect 23290 20204 23296 20256
rect 23348 20244 23354 20256
rect 23348 20216 23393 20244
rect 23348 20204 23354 20216
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 8386 20040 8392 20052
rect 8347 20012 8392 20040
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10008 20012 10333 20040
rect 10008 20000 10014 20012
rect 10321 20009 10333 20012
rect 10367 20040 10379 20043
rect 10686 20040 10692 20052
rect 10367 20012 10692 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 15286 20040 15292 20052
rect 11379 20012 15292 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 15654 20000 15660 20052
rect 15712 20040 15718 20052
rect 15712 20012 16528 20040
rect 15712 20000 15718 20012
rect 7006 19932 7012 19984
rect 7064 19972 7070 19984
rect 16500 19972 16528 20012
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17589 20043 17647 20049
rect 17589 20040 17601 20043
rect 17184 20012 17601 20040
rect 17184 20000 17190 20012
rect 17589 20009 17601 20012
rect 17635 20009 17647 20043
rect 17589 20003 17647 20009
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19484 20012 19901 20040
rect 19484 20000 19490 20012
rect 19889 20009 19901 20012
rect 19935 20040 19947 20043
rect 19978 20040 19984 20052
rect 19935 20012 19984 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20990 20000 20996 20052
rect 21048 20040 21054 20052
rect 21085 20043 21143 20049
rect 21085 20040 21097 20043
rect 21048 20012 21097 20040
rect 21048 20000 21054 20012
rect 21085 20009 21097 20012
rect 21131 20009 21143 20043
rect 21085 20003 21143 20009
rect 32214 19972 32220 19984
rect 7064 19944 9904 19972
rect 7064 19932 7070 19944
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 9766 19904 9772 19916
rect 9723 19876 9772 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 9876 19913 9904 19944
rect 9968 19944 16436 19972
rect 16500 19944 20300 19972
rect 9861 19907 9919 19913
rect 9861 19873 9873 19907
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 5592 19808 7113 19836
rect 5592 19796 5598 19808
rect 7101 19805 7113 19808
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 8386 19836 8392 19848
rect 7975 19808 8392 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8619 19808 9260 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 7193 19771 7251 19777
rect 7193 19737 7205 19771
rect 7239 19768 7251 19771
rect 9030 19768 9036 19780
rect 7239 19740 9036 19768
rect 7239 19737 7251 19740
rect 7193 19731 7251 19737
rect 9030 19728 9036 19740
rect 9088 19728 9094 19780
rect 7745 19703 7803 19709
rect 7745 19669 7757 19703
rect 7791 19700 7803 19703
rect 8478 19700 8484 19712
rect 7791 19672 8484 19700
rect 7791 19669 7803 19672
rect 7745 19663 7803 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 9122 19700 9128 19712
rect 8628 19672 9128 19700
rect 8628 19660 8634 19672
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 9232 19700 9260 19808
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 9968 19836 9996 19944
rect 12069 19907 12127 19913
rect 12069 19873 12081 19907
rect 12115 19904 12127 19907
rect 12434 19904 12440 19916
rect 12115 19876 12440 19904
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 12584 19876 12629 19904
rect 12584 19864 12590 19876
rect 14734 19864 14740 19916
rect 14792 19904 14798 19916
rect 15105 19907 15163 19913
rect 15105 19904 15117 19907
rect 14792 19876 15117 19904
rect 14792 19864 14798 19876
rect 15105 19873 15117 19876
rect 15151 19873 15163 19907
rect 16206 19904 16212 19916
rect 16167 19876 16212 19904
rect 15105 19867 15163 19873
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16408 19913 16436 19944
rect 16393 19907 16451 19913
rect 16393 19873 16405 19907
rect 16439 19873 16451 19907
rect 17586 19904 17592 19916
rect 16393 19867 16451 19873
rect 16546 19876 17592 19904
rect 11514 19836 11520 19848
rect 9364 19808 9996 19836
rect 11475 19808 11520 19836
rect 9364 19796 9370 19808
rect 11514 19796 11520 19808
rect 11572 19796 11578 19848
rect 14274 19796 14280 19848
rect 14332 19836 14338 19848
rect 14550 19836 14556 19848
rect 14332 19808 14556 19836
rect 14332 19796 14338 19808
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19836 15807 19839
rect 16298 19836 16304 19848
rect 15795 19808 16304 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 16298 19796 16304 19808
rect 16356 19836 16362 19848
rect 16546 19836 16574 19876
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 19242 19904 19248 19916
rect 18279 19876 19248 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 16356 19808 16574 19836
rect 17497 19839 17555 19845
rect 16356 19796 16362 19808
rect 17497 19805 17509 19839
rect 17543 19805 17555 19839
rect 18414 19836 18420 19848
rect 18375 19808 18420 19836
rect 17497 19799 17555 19805
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 12161 19771 12219 19777
rect 12161 19768 12173 19771
rect 9456 19740 12173 19768
rect 9456 19728 9462 19740
rect 12161 19737 12173 19740
rect 12207 19737 12219 19771
rect 15194 19768 15200 19780
rect 15155 19740 15200 19768
rect 12161 19731 12219 19737
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 15470 19728 15476 19780
rect 15528 19768 15534 19780
rect 17512 19768 17540 19799
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 19426 19796 19432 19848
rect 19484 19836 19490 19848
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 19484 19808 19533 19836
rect 19484 19796 19490 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 15528 19740 17540 19768
rect 15528 19728 15534 19740
rect 18690 19728 18696 19780
rect 18748 19768 18754 19780
rect 19720 19768 19748 19799
rect 18748 19740 19748 19768
rect 18748 19728 18754 19740
rect 10042 19700 10048 19712
rect 9232 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 13538 19700 13544 19712
rect 13499 19672 13544 19700
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 15838 19700 15844 19712
rect 14415 19672 15844 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19700 16911 19703
rect 18230 19700 18236 19712
rect 16899 19672 18236 19700
rect 16899 19669 16911 19672
rect 16853 19663 16911 19669
rect 18230 19660 18236 19672
rect 18288 19700 18294 19712
rect 18877 19703 18935 19709
rect 18877 19700 18889 19703
rect 18288 19672 18889 19700
rect 18288 19660 18294 19672
rect 18877 19669 18889 19672
rect 18923 19669 18935 19703
rect 20272 19700 20300 19944
rect 20732 19944 32220 19972
rect 20732 19913 20760 19944
rect 32214 19932 32220 19944
rect 32272 19932 32278 19984
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19873 20775 19907
rect 20898 19904 20904 19916
rect 20859 19876 20904 19904
rect 20717 19867 20775 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 32398 19904 32404 19916
rect 21959 19876 32404 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 32398 19864 32404 19876
rect 32456 19864 32462 19916
rect 23014 19836 23020 19848
rect 22975 19808 23020 19836
rect 23014 19796 23020 19808
rect 23072 19796 23078 19848
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 36998 19836 37004 19848
rect 29779 19808 37004 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 36998 19796 37004 19808
rect 37056 19796 37062 19848
rect 22002 19768 22008 19780
rect 21963 19740 22008 19768
rect 22002 19728 22008 19740
rect 22060 19728 22066 19780
rect 22557 19771 22615 19777
rect 22557 19768 22569 19771
rect 22112 19740 22569 19768
rect 22112 19700 22140 19740
rect 22557 19737 22569 19740
rect 22603 19768 22615 19771
rect 24946 19768 24952 19780
rect 22603 19740 24952 19768
rect 22603 19737 22615 19740
rect 22557 19731 22615 19737
rect 24946 19728 24952 19740
rect 25004 19728 25010 19780
rect 20272 19672 22140 19700
rect 18877 19663 18935 19669
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 23109 19703 23167 19709
rect 23109 19700 23121 19703
rect 22244 19672 23121 19700
rect 22244 19660 22250 19672
rect 23109 19669 23121 19672
rect 23155 19669 23167 19703
rect 23109 19663 23167 19669
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 29825 19703 29883 19709
rect 29825 19700 29837 19703
rect 27672 19672 29837 19700
rect 27672 19660 27678 19672
rect 29825 19669 29837 19672
rect 29871 19669 29883 19703
rect 29825 19663 29883 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 5166 19496 5172 19508
rect 1627 19468 5172 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 6733 19499 6791 19505
rect 6733 19465 6745 19499
rect 6779 19465 6791 19499
rect 6733 19459 6791 19465
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 9582 19496 9588 19508
rect 7423 19468 9588 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 6748 19428 6776 19459
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 12342 19496 12348 19508
rect 12303 19468 12348 19496
rect 12342 19456 12348 19468
rect 12400 19496 12406 19508
rect 13633 19499 13691 19505
rect 13633 19496 13645 19499
rect 12400 19468 13645 19496
rect 12400 19456 12406 19468
rect 13633 19465 13645 19468
rect 13679 19465 13691 19499
rect 13633 19459 13691 19465
rect 14645 19499 14703 19505
rect 14645 19465 14657 19499
rect 14691 19496 14703 19499
rect 15930 19496 15936 19508
rect 14691 19468 15936 19496
rect 14691 19465 14703 19468
rect 14645 19459 14703 19465
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 18690 19496 18696 19508
rect 18651 19468 18696 19496
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 23290 19496 23296 19508
rect 18892 19468 23296 19496
rect 8478 19428 8484 19440
rect 6748 19400 7604 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 5810 19360 5816 19372
rect 5771 19332 5816 19360
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 5951 19332 6868 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 6840 19292 6868 19332
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7576 19369 7604 19400
rect 8036 19400 8484 19428
rect 8036 19369 8064 19400
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 9766 19428 9772 19440
rect 8680 19400 9772 19428
rect 7561 19363 7619 19369
rect 6972 19332 7017 19360
rect 6972 19320 6978 19332
rect 7561 19329 7573 19363
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8570 19360 8576 19372
rect 8159 19332 8576 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 8202 19292 8208 19304
rect 6840 19264 8208 19292
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8680 19233 8708 19400
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 17954 19428 17960 19440
rect 15396 19400 17960 19428
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19360 9551 19363
rect 9858 19360 9864 19372
rect 9539 19332 9864 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 11330 19360 11336 19372
rect 9968 19332 11336 19360
rect 9968 19301 9996 19332
rect 11330 19320 11336 19332
rect 11388 19360 11394 19372
rect 12986 19360 12992 19372
rect 11388 19332 12434 19360
rect 12947 19332 12992 19360
rect 11388 19320 11394 19332
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10138 19295 10196 19301
rect 10138 19261 10150 19295
rect 10184 19261 10196 19295
rect 10138 19255 10196 19261
rect 8665 19227 8723 19233
rect 8665 19193 8677 19227
rect 8711 19193 8723 19227
rect 8665 19187 8723 19193
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 10152 19224 10180 19255
rect 11606 19252 11612 19304
rect 11664 19292 11670 19304
rect 11701 19295 11759 19301
rect 11701 19292 11713 19295
rect 11664 19264 11713 19292
rect 11664 19252 11670 19264
rect 11701 19261 11713 19264
rect 11747 19261 11759 19295
rect 11701 19255 11759 19261
rect 11790 19252 11796 19304
rect 11848 19292 11854 19304
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11848 19264 11897 19292
rect 11848 19252 11854 19264
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 12406 19292 12434 19332
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 13096 19332 13308 19360
rect 13096 19292 13124 19332
rect 12406 19264 13124 19292
rect 13173 19295 13231 19301
rect 11885 19255 11943 19261
rect 13173 19261 13185 19295
rect 13219 19261 13231 19295
rect 13280 19292 13308 19332
rect 15194 19292 15200 19304
rect 13280 19264 15200 19292
rect 13173 19255 13231 19261
rect 10318 19224 10324 19236
rect 8812 19196 10180 19224
rect 10279 19196 10324 19224
rect 8812 19184 8818 19196
rect 10318 19184 10324 19196
rect 10376 19184 10382 19236
rect 10594 19184 10600 19236
rect 10652 19224 10658 19236
rect 13188 19224 13216 19255
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15396 19292 15424 19400
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16908 19332 17049 19360
rect 16908 19320 16914 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17678 19360 17684 19372
rect 17639 19332 17684 19360
rect 17037 19323 17095 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 18892 19369 18920 19468
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 31846 19428 31852 19440
rect 20732 19400 31852 19428
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19024 19332 19993 19360
rect 19024 19320 19030 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20732 19369 20760 19400
rect 31846 19388 31852 19400
rect 31904 19388 31910 19440
rect 20717 19363 20775 19369
rect 20496 19332 20668 19360
rect 20496 19320 20502 19332
rect 15335 19264 15424 19292
rect 15473 19295 15531 19301
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15473 19261 15485 19295
rect 15519 19261 15531 19295
rect 17218 19292 17224 19304
rect 17179 19264 17224 19292
rect 15473 19255 15531 19261
rect 10652 19196 13216 19224
rect 10652 19184 10658 19196
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 15488 19224 15516 19255
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19300 19264 19349 19292
rect 19300 19252 19306 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19518 19292 19524 19304
rect 19479 19264 19524 19292
rect 19337 19255 19395 19261
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 20640 19292 20668 19332
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 21361 19363 21419 19369
rect 21361 19360 21373 19363
rect 20717 19323 20775 19329
rect 20824 19332 21373 19360
rect 20824 19292 20852 19332
rect 21361 19329 21373 19332
rect 21407 19360 21419 19363
rect 22649 19363 22707 19369
rect 22649 19360 22661 19363
rect 21407 19332 22661 19360
rect 21407 19329 21419 19332
rect 21361 19323 21419 19329
rect 22649 19329 22661 19332
rect 22695 19329 22707 19363
rect 22649 19323 22707 19329
rect 23198 19320 23204 19372
rect 23256 19360 23262 19372
rect 23293 19363 23351 19369
rect 23293 19360 23305 19363
rect 23256 19332 23305 19360
rect 23256 19320 23262 19332
rect 23293 19329 23305 19332
rect 23339 19329 23351 19363
rect 23293 19323 23351 19329
rect 20640 19264 20852 19292
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19261 20959 19295
rect 22002 19292 22008 19304
rect 21963 19264 22008 19292
rect 20901 19255 20959 19261
rect 17586 19224 17592 19236
rect 13964 19196 15516 19224
rect 15580 19196 17592 19224
rect 13964 19184 13970 19196
rect 9306 19156 9312 19168
rect 9267 19128 9312 19156
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 13262 19156 13268 19168
rect 9732 19128 13268 19156
rect 9732 19116 9738 19128
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 15580 19156 15608 19196
rect 17586 19184 17592 19196
rect 17644 19184 17650 19236
rect 20916 19224 20944 19255
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 22189 19295 22247 19301
rect 22189 19261 22201 19295
rect 22235 19261 22247 19295
rect 22189 19255 22247 19261
rect 22094 19224 22100 19236
rect 20916 19196 22100 19224
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 22204 19224 22232 19255
rect 23109 19227 23167 19233
rect 23109 19224 23121 19227
rect 22204 19196 23121 19224
rect 23109 19193 23121 19196
rect 23155 19193 23167 19227
rect 23109 19187 23167 19193
rect 13504 19128 15608 19156
rect 13504 19116 13510 19128
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 15930 19156 15936 19168
rect 15804 19128 15936 19156
rect 15804 19116 15810 19128
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 23014 19156 23020 19168
rect 18380 19128 23020 19156
rect 18380 19116 18386 19128
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 8754 18952 8760 18964
rect 7239 18924 8760 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 10318 18952 10324 18964
rect 9999 18924 10324 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 13906 18952 13912 18964
rect 10551 18924 13912 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14642 18912 14648 18964
rect 14700 18952 14706 18964
rect 15013 18955 15071 18961
rect 15013 18952 15025 18955
rect 14700 18924 15025 18952
rect 14700 18912 14706 18924
rect 15013 18921 15025 18924
rect 15059 18921 15071 18955
rect 15013 18915 15071 18921
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 16114 18952 16120 18964
rect 15703 18924 16120 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16301 18955 16359 18961
rect 16301 18921 16313 18955
rect 16347 18952 16359 18955
rect 17310 18952 17316 18964
rect 16347 18924 17316 18952
rect 16347 18921 16359 18924
rect 16301 18915 16359 18921
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 18877 18955 18935 18961
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 18966 18952 18972 18964
rect 18923 18924 18972 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 13446 18884 13452 18896
rect 8404 18856 13452 18884
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 6972 18788 7788 18816
rect 6972 18776 6978 18788
rect 6638 18748 6644 18760
rect 6599 18720 6644 18748
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7282 18748 7288 18760
rect 7147 18720 7288 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7760 18757 7788 18788
rect 8404 18757 8432 18856
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 13541 18887 13599 18893
rect 13541 18853 13553 18887
rect 13587 18884 13599 18887
rect 13814 18884 13820 18896
rect 13587 18856 13820 18884
rect 13587 18853 13599 18856
rect 13541 18847 13599 18853
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 15194 18844 15200 18896
rect 15252 18884 15258 18896
rect 15252 18856 15332 18884
rect 15252 18844 15258 18856
rect 8478 18776 8484 18828
rect 8536 18816 8542 18828
rect 9309 18819 9367 18825
rect 9309 18816 9321 18819
rect 8536 18788 9321 18816
rect 8536 18776 8542 18788
rect 9309 18785 9321 18788
rect 9355 18785 9367 18819
rect 9309 18779 9367 18785
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 11241 18819 11299 18825
rect 11241 18816 11253 18819
rect 9640 18788 11253 18816
rect 9640 18776 9646 18788
rect 11241 18785 11253 18788
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 11848 18788 12572 18816
rect 11848 18776 11854 18788
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9508 18680 9536 18711
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9732 18720 10425 18748
rect 9732 18708 9738 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11330 18748 11336 18760
rect 11103 18720 11336 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 12250 18748 12256 18760
rect 12211 18720 12256 18748
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12544 18748 12572 18788
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 15304 18816 15332 18856
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15746 18884 15752 18896
rect 15528 18856 15752 18884
rect 15528 18844 15534 18856
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 17586 18884 17592 18896
rect 17547 18856 17592 18884
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 16390 18816 16396 18828
rect 12676 18788 15240 18816
rect 15304 18788 16396 18816
rect 12676 18776 12682 18788
rect 14553 18751 14611 18757
rect 12544 18720 12848 18748
rect 12820 18680 12848 18720
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 15102 18748 15108 18760
rect 14599 18720 15108 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15212 18757 15240 18788
rect 16390 18776 16396 18788
rect 16448 18776 16454 18828
rect 17037 18819 17095 18825
rect 17037 18785 17049 18819
rect 17083 18816 17095 18819
rect 18892 18816 18920 18915
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 23017 18955 23075 18961
rect 23017 18952 23029 18955
rect 20312 18924 23029 18952
rect 20312 18912 20318 18924
rect 23017 18921 23029 18924
rect 23063 18921 23075 18955
rect 33594 18952 33600 18964
rect 33555 18924 33600 18952
rect 23017 18915 23075 18921
rect 33594 18912 33600 18924
rect 33652 18912 33658 18964
rect 25958 18884 25964 18896
rect 19628 18856 25964 18884
rect 17083 18788 18920 18816
rect 17083 18785 17095 18788
rect 17037 18779 17095 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19484 18788 19533 18816
rect 19484 18776 19490 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 15197 18751 15255 18757
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15838 18748 15844 18760
rect 15799 18720 15844 18748
rect 15197 18711 15255 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18748 16543 18751
rect 16850 18748 16856 18760
rect 16531 18720 16856 18748
rect 16531 18717 16543 18720
rect 16485 18711 16543 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 19334 18748 19340 18760
rect 18463 18720 19340 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 6472 18652 9536 18680
rect 10152 18652 12756 18680
rect 12820 18652 13001 18680
rect 6472 18621 6500 18652
rect 6457 18615 6515 18621
rect 6457 18581 6469 18615
rect 6503 18581 6515 18615
rect 6457 18575 6515 18581
rect 7837 18615 7895 18621
rect 7837 18581 7849 18615
rect 7883 18612 7895 18615
rect 8294 18612 8300 18624
rect 7883 18584 8300 18612
rect 7883 18581 7895 18584
rect 7837 18575 7895 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 8478 18612 8484 18624
rect 8439 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 10152 18612 10180 18652
rect 11698 18612 11704 18624
rect 8628 18584 10180 18612
rect 11659 18584 11704 18612
rect 8628 18572 8634 18584
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12618 18612 12624 18624
rect 12391 18584 12624 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12728 18612 12756 18652
rect 12989 18649 13001 18652
rect 13035 18649 13047 18683
rect 12989 18643 13047 18649
rect 13081 18683 13139 18689
rect 13081 18649 13093 18683
rect 13127 18649 13139 18683
rect 13081 18643 13139 18649
rect 13096 18612 13124 18643
rect 13354 18640 13360 18692
rect 13412 18680 13418 18692
rect 16666 18680 16672 18692
rect 13412 18652 16672 18680
rect 13412 18640 13418 18652
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 17126 18680 17132 18692
rect 17087 18652 17132 18680
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17954 18640 17960 18692
rect 18012 18680 18018 18692
rect 18248 18680 18276 18711
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19628 18680 19656 18856
rect 25958 18844 25964 18856
rect 26016 18844 26022 18896
rect 20806 18816 20812 18828
rect 20767 18788 20812 18816
rect 20806 18776 20812 18788
rect 20864 18816 20870 18828
rect 21637 18819 21695 18825
rect 20864 18788 21404 18816
rect 20864 18776 20870 18788
rect 21376 18748 21404 18788
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 22002 18816 22008 18828
rect 21683 18788 22008 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 22002 18776 22008 18788
rect 22060 18776 22066 18828
rect 28902 18816 28908 18828
rect 22112 18788 28908 18816
rect 22112 18748 22140 18788
rect 28902 18776 28908 18788
rect 28960 18776 28966 18828
rect 21376 18720 22140 18748
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22244 18720 22937 18748
rect 22244 18708 22250 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 33410 18708 33416 18760
rect 33468 18748 33474 18760
rect 33781 18751 33839 18757
rect 33781 18748 33793 18751
rect 33468 18720 33793 18748
rect 33468 18708 33474 18720
rect 33781 18717 33793 18720
rect 33827 18717 33839 18751
rect 33781 18711 33839 18717
rect 18012 18652 19656 18680
rect 20533 18683 20591 18689
rect 18012 18640 18018 18652
rect 20533 18649 20545 18683
rect 20579 18649 20591 18683
rect 20533 18643 20591 18649
rect 12728 18584 13124 18612
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 14274 18612 14280 18624
rect 13320 18584 14280 18612
rect 13320 18572 13326 18584
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 14369 18615 14427 18621
rect 14369 18581 14381 18615
rect 14415 18612 14427 18615
rect 16206 18612 16212 18624
rect 14415 18584 16212 18612
rect 14415 18581 14427 18584
rect 14369 18575 14427 18581
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 20548 18612 20576 18643
rect 20622 18640 20628 18692
rect 20680 18680 20686 18692
rect 20680 18652 20725 18680
rect 20680 18640 20686 18652
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 20548 18584 22293 18612
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 7193 18411 7251 18417
rect 7193 18408 7205 18411
rect 6696 18380 7205 18408
rect 6696 18368 6702 18380
rect 7193 18377 7205 18380
rect 7239 18377 7251 18411
rect 7193 18371 7251 18377
rect 9125 18411 9183 18417
rect 9125 18377 9137 18411
rect 9171 18377 9183 18411
rect 15105 18411 15163 18417
rect 9125 18371 9183 18377
rect 10244 18380 12296 18408
rect 9140 18340 9168 18371
rect 9140 18312 9996 18340
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7340 18244 7389 18272
rect 7340 18232 7346 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18272 8079 18275
rect 8386 18272 8392 18284
rect 8067 18244 8392 18272
rect 8067 18241 8079 18244
rect 8021 18235 8079 18241
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 8662 18272 8668 18284
rect 8623 18244 8668 18272
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9306 18272 9312 18284
rect 9267 18244 9312 18272
rect 9306 18232 9312 18244
rect 9364 18232 9370 18284
rect 9968 18281 9996 18312
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 10244 18204 10272 18380
rect 10594 18300 10600 18352
rect 10652 18340 10658 18352
rect 10652 18312 10697 18340
rect 10652 18300 10658 18312
rect 12268 18281 12296 18380
rect 15105 18377 15117 18411
rect 15151 18408 15163 18411
rect 16022 18408 16028 18420
rect 15151 18380 16028 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 18414 18408 18420 18420
rect 18375 18380 18420 18408
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 19978 18408 19984 18420
rect 19659 18380 19984 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 21269 18411 21327 18417
rect 21269 18408 21281 18411
rect 20680 18380 21281 18408
rect 20680 18368 20686 18380
rect 21269 18377 21281 18380
rect 21315 18377 21327 18411
rect 21269 18371 21327 18377
rect 22005 18411 22063 18417
rect 22005 18377 22017 18411
rect 22051 18377 22063 18411
rect 33410 18408 33416 18420
rect 33371 18380 33416 18408
rect 22005 18371 22063 18377
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 12676 18312 17141 18340
rect 12676 18300 12682 18312
rect 17129 18309 17141 18312
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 17681 18343 17739 18349
rect 17681 18309 17693 18343
rect 17727 18340 17739 18343
rect 19242 18340 19248 18352
rect 17727 18312 19248 18340
rect 17727 18309 17739 18312
rect 17681 18303 17739 18309
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 20254 18340 20260 18352
rect 20215 18312 20260 18340
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 20806 18340 20812 18352
rect 20767 18312 20812 18340
rect 20806 18300 20812 18312
rect 20864 18300 20870 18352
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 16114 18272 16120 18284
rect 12943 18244 15976 18272
rect 16075 18244 16120 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 9088 18176 10272 18204
rect 10505 18207 10563 18213
rect 9088 18164 9094 18176
rect 10505 18173 10517 18207
rect 10551 18204 10563 18207
rect 11698 18204 11704 18216
rect 10551 18176 11704 18204
rect 10551 18173 10563 18176
rect 10505 18167 10563 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 12342 18164 12348 18216
rect 12400 18204 12406 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12400 18176 12449 18204
rect 12400 18164 12406 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 13354 18204 13360 18216
rect 13315 18176 13360 18204
rect 12437 18167 12495 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 13504 18176 13553 18204
rect 13504 18164 13510 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 13541 18167 13599 18173
rect 13924 18176 14473 18204
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 9582 18136 9588 18148
rect 7883 18108 9588 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 9766 18136 9772 18148
rect 9727 18108 9772 18136
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 11057 18139 11115 18145
rect 11057 18136 11069 18139
rect 10100 18108 11069 18136
rect 10100 18096 10106 18108
rect 11057 18105 11069 18108
rect 11103 18105 11115 18139
rect 11057 18099 11115 18105
rect 11790 18096 11796 18148
rect 11848 18136 11854 18148
rect 13725 18139 13783 18145
rect 13725 18136 13737 18139
rect 11848 18108 13737 18136
rect 11848 18096 11854 18108
rect 13725 18105 13737 18108
rect 13771 18105 13783 18139
rect 13725 18099 13783 18105
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 5534 18068 5540 18080
rect 1627 18040 5540 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 8481 18071 8539 18077
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 11146 18068 11152 18080
rect 8527 18040 11152 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 13924 18068 13952 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14642 18204 14648 18216
rect 14603 18176 14648 18204
rect 14461 18167 14519 18173
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 15948 18204 15976 18244
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 18322 18272 18328 18284
rect 18283 18244 18328 18272
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 21453 18275 21511 18281
rect 19076 18244 19334 18272
rect 17034 18204 17040 18216
rect 15948 18176 16896 18204
rect 16995 18176 17040 18204
rect 14274 18096 14280 18148
rect 14332 18136 14338 18148
rect 16390 18136 16396 18148
rect 14332 18108 16396 18136
rect 14332 18096 14338 18108
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 16868 18136 16896 18176
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 18969 18207 19027 18213
rect 18969 18204 18981 18207
rect 18932 18176 18981 18204
rect 18932 18164 18938 18176
rect 18969 18173 18981 18176
rect 19015 18173 19027 18207
rect 18969 18167 19027 18173
rect 17402 18136 17408 18148
rect 16868 18108 17408 18136
rect 17402 18096 17408 18108
rect 17460 18136 17466 18148
rect 19076 18136 19104 18244
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19306 18204 19334 18244
rect 21453 18241 21465 18275
rect 21499 18272 21511 18275
rect 22020 18272 22048 18371
rect 33410 18368 33416 18380
rect 33468 18368 33474 18420
rect 22186 18272 22192 18284
rect 21499 18244 22048 18272
rect 22147 18244 22192 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 22646 18272 22652 18284
rect 22607 18244 22652 18272
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 23290 18272 23296 18284
rect 23251 18244 23296 18272
rect 23290 18232 23296 18244
rect 23348 18232 23354 18284
rect 33321 18275 33379 18281
rect 33321 18272 33333 18275
rect 31726 18244 33333 18272
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 19306 18176 20177 18204
rect 19153 18167 19211 18173
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 17460 18108 19104 18136
rect 19168 18136 19196 18167
rect 19168 18108 20024 18136
rect 17460 18096 17466 18108
rect 12492 18040 13952 18068
rect 16209 18071 16267 18077
rect 12492 18028 12498 18040
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 17862 18068 17868 18080
rect 16255 18040 17868 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 19702 18068 19708 18080
rect 18472 18040 19708 18068
rect 18472 18028 18478 18040
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 19996 18068 20024 18108
rect 22094 18096 22100 18148
rect 22152 18136 22158 18148
rect 31726 18136 31754 18244
rect 33321 18241 33333 18244
rect 33367 18241 33379 18275
rect 33321 18235 33379 18241
rect 22152 18108 31754 18136
rect 22152 18096 22158 18108
rect 22741 18071 22799 18077
rect 22741 18068 22753 18071
rect 19996 18040 22753 18068
rect 22741 18037 22753 18040
rect 22787 18037 22799 18071
rect 23382 18068 23388 18080
rect 23343 18040 23388 18068
rect 22741 18031 22799 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 8662 17864 8668 17876
rect 8435 17836 8668 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 9217 17867 9275 17873
rect 9217 17864 9229 17867
rect 8904 17836 9229 17864
rect 8904 17824 8910 17836
rect 9217 17833 9229 17836
rect 9263 17833 9275 17867
rect 9217 17827 9275 17833
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 10962 17864 10968 17876
rect 9640 17836 10968 17864
rect 9640 17824 9646 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11698 17864 11704 17876
rect 11659 17836 11704 17864
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12434 17864 12440 17876
rect 12124 17836 12440 17864
rect 12124 17824 12130 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 16209 17867 16267 17873
rect 16209 17833 16221 17867
rect 16255 17864 16267 17867
rect 17218 17864 17224 17876
rect 16255 17836 17224 17864
rect 16255 17833 16267 17836
rect 16209 17827 16267 17833
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19484 17836 19717 17864
rect 19484 17824 19490 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 23382 17864 23388 17876
rect 19705 17827 19763 17833
rect 20180 17836 23388 17864
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 17313 17799 17371 17805
rect 17313 17796 17325 17799
rect 8352 17768 11284 17796
rect 8352 17756 8358 17768
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 9582 17728 9588 17740
rect 8996 17700 9588 17728
rect 8996 17688 9002 17700
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9950 17728 9956 17740
rect 9911 17700 9956 17728
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 11256 17737 11284 17768
rect 12728 17768 17325 17796
rect 12728 17737 12756 17768
rect 17313 17765 17325 17768
rect 17359 17796 17371 17799
rect 18046 17796 18052 17808
rect 17359 17768 18052 17796
rect 17359 17765 17371 17768
rect 17313 17759 17371 17765
rect 18046 17756 18052 17768
rect 18104 17756 18110 17808
rect 20180 17796 20208 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 18340 17768 20208 17796
rect 20993 17799 21051 17805
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 10100 17700 10241 17728
rect 10100 17688 10106 17700
rect 10229 17697 10241 17700
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17697 11299 17731
rect 11241 17691 11299 17697
rect 12713 17731 12771 17737
rect 12713 17697 12725 17731
rect 12759 17697 12771 17731
rect 12713 17691 12771 17697
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 12989 17731 13047 17737
rect 12989 17728 13001 17731
rect 12860 17700 13001 17728
rect 12860 17688 12866 17700
rect 12989 17697 13001 17700
rect 13035 17697 13047 17731
rect 12989 17691 13047 17697
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13136 17700 13400 17728
rect 13136 17688 13142 17700
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17660 7343 17663
rect 7650 17660 7656 17672
rect 7331 17632 7656 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8662 17660 8668 17672
rect 8619 17632 8668 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9088 17632 9413 17660
rect 9088 17620 9094 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17660 11115 17663
rect 11974 17660 11980 17672
rect 11103 17632 11980 17660
rect 11103 17629 11115 17632
rect 11057 17623 11115 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 13372 17660 13400 17700
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 18340 17737 18368 17768
rect 20993 17765 21005 17799
rect 21039 17796 21051 17799
rect 21266 17796 21272 17808
rect 21039 17768 21272 17796
rect 21039 17765 21051 17768
rect 20993 17759 21051 17765
rect 21266 17756 21272 17768
rect 21324 17756 21330 17808
rect 27614 17796 27620 17808
rect 21560 17768 27620 17796
rect 17037 17731 17095 17737
rect 17037 17728 17049 17731
rect 13872 17700 17049 17728
rect 13872 17688 13878 17700
rect 17037 17697 17049 17700
rect 17083 17697 17095 17731
rect 17037 17691 17095 17697
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 19484 17700 20453 17728
rect 19484 17688 19490 17700
rect 20441 17697 20453 17700
rect 20487 17728 20499 17731
rect 20487 17700 21128 17728
rect 20487 17697 20499 17700
rect 20441 17691 20499 17697
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13372 17632 14289 17660
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 5261 17595 5319 17601
rect 5261 17561 5273 17595
rect 5307 17592 5319 17595
rect 9122 17592 9128 17604
rect 5307 17564 9128 17592
rect 5307 17561 5319 17564
rect 5261 17555 5319 17561
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 9272 17564 10057 17592
rect 9272 17552 9278 17564
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 10318 17552 10324 17604
rect 10376 17592 10382 17604
rect 11606 17592 11612 17604
rect 10376 17564 11612 17592
rect 10376 17552 10382 17564
rect 11606 17552 11612 17564
rect 11664 17552 11670 17604
rect 12805 17595 12863 17601
rect 12805 17561 12817 17595
rect 12851 17592 12863 17595
rect 12894 17592 12900 17604
rect 12851 17564 12900 17592
rect 12851 17561 12863 17564
rect 12805 17555 12863 17561
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 6972 17496 7113 17524
rect 6972 17484 6978 17496
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7101 17487 7159 17493
rect 7745 17527 7803 17533
rect 7745 17493 7757 17527
rect 7791 17524 7803 17527
rect 11054 17524 11060 17536
rect 7791 17496 11060 17524
rect 7791 17493 7803 17496
rect 7745 17487 7803 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 14476 17524 14504 17623
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16264 17632 16405 17660
rect 16264 17620 16270 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17660 16911 17663
rect 17954 17660 17960 17672
rect 16899 17632 17960 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 19794 17660 19800 17672
rect 18187 17632 19800 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 20254 17660 20260 17672
rect 19935 17632 20260 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 14921 17595 14979 17601
rect 14921 17561 14933 17595
rect 14967 17592 14979 17595
rect 16574 17592 16580 17604
rect 14967 17564 16580 17592
rect 14967 17561 14979 17564
rect 14921 17555 14979 17561
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 17862 17552 17868 17604
rect 17920 17592 17926 17604
rect 20533 17595 20591 17601
rect 17920 17564 20392 17592
rect 17920 17552 17926 17564
rect 15562 17524 15568 17536
rect 11204 17496 14504 17524
rect 15523 17496 15568 17524
rect 11204 17484 11210 17496
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18785 17527 18843 17533
rect 18785 17524 18797 17527
rect 18012 17496 18797 17524
rect 18012 17484 18018 17496
rect 18785 17493 18797 17496
rect 18831 17493 18843 17527
rect 20364 17524 20392 17564
rect 20533 17561 20545 17595
rect 20579 17561 20591 17595
rect 20533 17555 20591 17561
rect 20548 17524 20576 17555
rect 20364 17496 20576 17524
rect 21100 17524 21128 17700
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21560 17669 21588 17768
rect 27614 17756 27620 17768
rect 27672 17756 27678 17808
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21324 17632 21557 17660
rect 21324 17620 21330 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21726 17660 21732 17672
rect 21687 17632 21732 17660
rect 21545 17623 21603 17629
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 21818 17620 21824 17672
rect 21876 17660 21882 17672
rect 22649 17663 22707 17669
rect 22649 17660 22661 17663
rect 21876 17632 22661 17660
rect 21876 17620 21882 17632
rect 22649 17629 22661 17632
rect 22695 17660 22707 17663
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 22695 17632 23489 17660
rect 22695 17629 22707 17632
rect 22649 17623 22707 17629
rect 23477 17629 23489 17632
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 22189 17527 22247 17533
rect 22189 17524 22201 17527
rect 21100 17496 22201 17524
rect 18785 17487 18843 17493
rect 22189 17493 22201 17496
rect 22235 17493 22247 17527
rect 22738 17524 22744 17536
rect 22699 17496 22744 17524
rect 22189 17487 22247 17493
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 23474 17524 23480 17536
rect 23339 17496 23480 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 7377 17323 7435 17329
rect 7377 17289 7389 17323
rect 7423 17289 7435 17323
rect 7377 17283 7435 17289
rect 8021 17323 8079 17329
rect 8021 17289 8033 17323
rect 8067 17320 8079 17323
rect 8067 17292 13676 17320
rect 8067 17289 8079 17292
rect 8021 17283 8079 17289
rect 7392 17252 7420 17283
rect 7392 17224 10732 17252
rect 6914 17184 6920 17196
rect 6875 17156 6920 17184
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8570 17184 8576 17196
rect 8251 17156 8576 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 7576 17116 7604 17147
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9766 17184 9772 17196
rect 8720 17156 9772 17184
rect 8720 17144 8726 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10704 17193 10732 17224
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 12437 17255 12495 17261
rect 12437 17252 12449 17255
rect 11020 17224 12449 17252
rect 11020 17212 11026 17224
rect 12437 17221 12449 17224
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 12989 17255 13047 17261
rect 12989 17252 13001 17255
rect 12860 17224 13001 17252
rect 12860 17212 12866 17224
rect 12989 17221 13001 17224
rect 13035 17221 13047 17255
rect 12989 17215 13047 17221
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17153 10747 17187
rect 13446 17184 13452 17196
rect 13407 17156 13452 17184
rect 10689 17147 10747 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 13648 17193 13676 17292
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16908 17292 16957 17320
rect 16908 17280 16914 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 19426 17320 19432 17332
rect 19387 17292 19432 17320
rect 16945 17283 17003 17289
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20312 17292 21097 17320
rect 20312 17280 20318 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 21085 17283 21143 17289
rect 15286 17252 15292 17264
rect 15247 17224 15292 17252
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 15562 17212 15568 17264
rect 15620 17252 15626 17264
rect 20070 17252 20076 17264
rect 15620 17224 17632 17252
rect 20031 17224 20076 17252
rect 15620 17212 15626 17224
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 16298 17184 16304 17196
rect 15887 17156 16304 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 17604 17193 17632 17224
rect 20070 17212 20076 17224
rect 20128 17212 20134 17264
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 8294 17116 8300 17128
rect 7576 17088 8300 17116
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 9398 17116 9404 17128
rect 9355 17088 9404 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 6733 17051 6791 17057
rect 6733 17017 6745 17051
rect 6779 17048 6791 17051
rect 9508 17048 9536 17079
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 9640 17088 10517 17116
rect 9640 17076 9646 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12345 17119 12403 17125
rect 12345 17116 12357 17119
rect 11940 17088 12357 17116
rect 11940 17076 11946 17088
rect 12345 17085 12357 17088
rect 12391 17116 12403 17119
rect 15194 17116 15200 17128
rect 12391 17088 13860 17116
rect 15155 17088 15200 17116
rect 12391 17085 12403 17088
rect 12345 17079 12403 17085
rect 13832 17057 13860 17088
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 16114 17116 16120 17128
rect 15672 17088 16120 17116
rect 6779 17020 9536 17048
rect 13817 17051 13875 17057
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 13817 17017 13829 17051
rect 13863 17017 13875 17051
rect 13817 17011 13875 17017
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 15672 17048 15700 17088
rect 16114 17076 16120 17088
rect 16172 17116 16178 17128
rect 17144 17116 17172 17147
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 20680 17156 21281 17184
rect 20680 17144 20686 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21692 17156 22017 17184
rect 21692 17144 21698 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17184 22247 17187
rect 22738 17184 22744 17196
rect 22235 17156 22744 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 38013 17187 38071 17193
rect 38013 17184 38025 17187
rect 34572 17156 38025 17184
rect 34572 17144 34578 17156
rect 38013 17153 38025 17156
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 17770 17116 17776 17128
rect 16172 17088 17172 17116
rect 17731 17088 17776 17116
rect 16172 17076 16178 17088
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 18782 17116 18788 17128
rect 18743 17088 18788 17116
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 18966 17116 18972 17128
rect 18927 17088 18972 17116
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 20438 17116 20444 17128
rect 20027 17088 20444 17116
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 23106 17116 23112 17128
rect 23067 17088 23112 17116
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 23290 17116 23296 17128
rect 23251 17088 23296 17116
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 14884 17020 15700 17048
rect 14884 17008 14890 17020
rect 18598 17008 18604 17060
rect 18656 17048 18662 17060
rect 20533 17051 20591 17057
rect 20533 17048 20545 17051
rect 18656 17020 20545 17048
rect 18656 17008 18662 17020
rect 20533 17017 20545 17020
rect 20579 17017 20591 17051
rect 38194 17048 38200 17060
rect 38155 17020 38200 17048
rect 20533 17011 20591 17017
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 8754 16980 8760 16992
rect 8715 16952 8760 16980
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 11149 16983 11207 16989
rect 11149 16949 11161 16983
rect 11195 16980 11207 16983
rect 12526 16980 12532 16992
rect 11195 16952 12532 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 17954 16980 17960 16992
rect 16172 16952 17960 16980
rect 16172 16940 16178 16952
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 22649 16983 22707 16989
rect 22649 16949 22661 16983
rect 22695 16980 22707 16983
rect 23382 16980 23388 16992
rect 22695 16952 23388 16980
rect 22695 16949 22707 16952
rect 22649 16943 22707 16949
rect 23382 16940 23388 16952
rect 23440 16980 23446 16992
rect 23477 16983 23535 16989
rect 23477 16980 23489 16983
rect 23440 16952 23489 16980
rect 23440 16940 23446 16952
rect 23477 16949 23489 16952
rect 23523 16949 23535 16983
rect 23477 16943 23535 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 8386 16776 8392 16788
rect 8347 16748 8392 16776
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 9214 16776 9220 16788
rect 8680 16748 9220 16776
rect 7745 16711 7803 16717
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 8680 16708 8708 16748
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 16298 16776 16304 16788
rect 9824 16748 16304 16776
rect 9824 16736 9830 16748
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 17218 16736 17224 16788
rect 17276 16776 17282 16788
rect 21266 16776 21272 16788
rect 17276 16748 21272 16776
rect 17276 16736 17282 16748
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 21453 16779 21511 16785
rect 21453 16745 21465 16779
rect 21499 16776 21511 16779
rect 21726 16776 21732 16788
rect 21499 16748 21732 16776
rect 21499 16745 21511 16748
rect 21453 16739 21511 16745
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 23290 16776 23296 16788
rect 23251 16748 23296 16776
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 7791 16680 8708 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 8754 16668 8760 16720
rect 8812 16708 8818 16720
rect 15194 16708 15200 16720
rect 8812 16680 14320 16708
rect 15155 16680 15200 16708
rect 8812 16668 8818 16680
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 7024 16612 9321 16640
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16572 6607 16575
rect 7024 16572 7052 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 10318 16640 10324 16652
rect 9456 16612 10324 16640
rect 9456 16600 9462 16612
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10686 16640 10692 16652
rect 10428 16612 10692 16640
rect 6595 16544 7052 16572
rect 6595 16541 6607 16544
rect 6549 16535 6607 16541
rect 6472 16504 6500 16535
rect 7098 16532 7104 16584
rect 7156 16572 7162 16584
rect 7926 16572 7932 16584
rect 7156 16544 7201 16572
rect 7887 16544 7932 16572
rect 7156 16532 7162 16544
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8938 16572 8944 16584
rect 8619 16544 8944 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 10428 16572 10456 16612
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 10928 16612 11161 16640
rect 10928 16600 10934 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 12345 16643 12403 16649
rect 12345 16640 12357 16643
rect 11664 16612 12357 16640
rect 11664 16600 11670 16612
rect 12345 16609 12357 16612
rect 12391 16640 12403 16643
rect 12618 16640 12624 16652
rect 12391 16612 12624 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 13078 16640 13084 16652
rect 12768 16612 13084 16640
rect 12768 16600 12774 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 14292 16640 14320 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 17236 16708 17264 16736
rect 17402 16708 17408 16720
rect 16684 16680 17264 16708
rect 17363 16680 17408 16708
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 14292 16612 16129 16640
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16684 16640 16712 16680
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 18874 16708 18880 16720
rect 17972 16680 18880 16708
rect 17972 16652 18000 16680
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 20622 16708 20628 16720
rect 19536 16680 20628 16708
rect 16117 16603 16175 16609
rect 16224 16612 16712 16640
rect 9646 16544 10456 16572
rect 10597 16575 10655 16581
rect 7650 16504 7656 16516
rect 6472 16476 7656 16504
rect 7650 16464 7656 16476
rect 7708 16464 7714 16516
rect 7193 16439 7251 16445
rect 7193 16405 7205 16439
rect 7239 16436 7251 16439
rect 9646 16436 9674 16544
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 14734 16572 14740 16584
rect 13771 16544 14740 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 10410 16436 10416 16448
rect 7239 16408 9674 16436
rect 10371 16408 10416 16436
rect 7239 16405 7251 16408
rect 7193 16399 7251 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10612 16436 10640 16535
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16541 14887 16575
rect 15010 16572 15016 16584
rect 14971 16544 15016 16572
rect 14829 16535 14887 16541
rect 11238 16504 11244 16516
rect 11199 16476 11244 16504
rect 11238 16464 11244 16476
rect 11296 16464 11302 16516
rect 11790 16504 11796 16516
rect 11751 16476 11796 16504
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 14844 16504 14872 16535
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16224 16572 16252 16612
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16816 16612 17233 16640
rect 16816 16600 16822 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 17954 16640 17960 16652
rect 17221 16603 17279 16609
rect 17328 16612 17960 16640
rect 16574 16572 16580 16584
rect 15979 16544 16252 16572
rect 16535 16544 16580 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16574 16532 16580 16544
rect 16632 16572 16638 16584
rect 16942 16572 16948 16584
rect 16632 16544 16948 16572
rect 16632 16532 16638 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17328 16572 17356 16612
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18230 16640 18236 16652
rect 18191 16612 18236 16640
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 18598 16640 18604 16652
rect 18559 16612 18604 16640
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 19536 16581 19564 16680
rect 20622 16668 20628 16680
rect 20680 16668 20686 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 20809 16711 20867 16717
rect 20809 16708 20821 16711
rect 20772 16680 20821 16708
rect 20772 16668 20778 16680
rect 20809 16677 20821 16680
rect 20855 16708 20867 16711
rect 22002 16708 22008 16720
rect 20855 16680 22008 16708
rect 20855 16677 20867 16680
rect 20809 16671 20867 16677
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 22649 16643 22707 16649
rect 20303 16612 22048 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 17083 16544 17356 16572
rect 19521 16575 19579 16581
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 19521 16541 19533 16575
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 22020 16581 22048 16612
rect 22649 16609 22661 16643
rect 22695 16640 22707 16643
rect 23106 16640 23112 16652
rect 22695 16612 23112 16640
rect 22695 16609 22707 16612
rect 22649 16603 22707 16609
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 24912 16612 27108 16640
rect 24912 16600 24918 16612
rect 21361 16575 21419 16581
rect 21361 16572 21373 16575
rect 21048 16544 21373 16572
rect 21048 16532 21054 16544
rect 21361 16541 21373 16544
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 23474 16572 23480 16584
rect 23435 16544 23480 16572
rect 22005 16535 22063 16541
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 27080 16581 27108 16612
rect 27065 16575 27123 16581
rect 27065 16541 27077 16575
rect 27111 16541 27123 16575
rect 27065 16535 27123 16541
rect 33781 16575 33839 16581
rect 33781 16541 33793 16575
rect 33827 16541 33839 16575
rect 33781 16535 33839 16541
rect 15378 16504 15384 16516
rect 12492 16476 12537 16504
rect 14844 16476 15384 16504
rect 12492 16464 12498 16476
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 18322 16464 18328 16516
rect 18380 16504 18386 16516
rect 18380 16476 18425 16504
rect 18380 16464 18386 16476
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19613 16507 19671 16513
rect 19613 16504 19625 16507
rect 19392 16476 19625 16504
rect 19392 16464 19398 16476
rect 19613 16473 19625 16476
rect 19659 16473 19671 16507
rect 20346 16504 20352 16516
rect 20307 16476 20352 16504
rect 19613 16467 19671 16473
rect 20346 16464 20352 16476
rect 20404 16464 20410 16516
rect 27157 16507 27215 16513
rect 27157 16473 27169 16507
rect 27203 16504 27215 16507
rect 33796 16504 33824 16535
rect 27203 16476 33824 16504
rect 27203 16473 27215 16476
rect 27157 16467 27215 16473
rect 13354 16436 13360 16448
rect 10612 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 13814 16436 13820 16448
rect 13587 16408 13820 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 21542 16436 21548 16448
rect 15160 16408 21548 16436
rect 15160 16396 15166 16408
rect 21542 16396 21548 16408
rect 21600 16396 21606 16448
rect 33597 16439 33655 16445
rect 33597 16405 33609 16439
rect 33643 16436 33655 16439
rect 34514 16436 34520 16448
rect 33643 16408 34520 16436
rect 33643 16405 33655 16408
rect 33597 16399 33655 16405
rect 34514 16396 34520 16408
rect 34572 16396 34578 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 7926 16232 7932 16244
rect 7147 16204 7932 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 9677 16235 9735 16241
rect 9677 16232 9689 16235
rect 8628 16204 9689 16232
rect 8628 16192 8634 16204
rect 9677 16201 9689 16204
rect 9723 16201 9735 16235
rect 11422 16232 11428 16244
rect 9677 16195 9735 16201
rect 10336 16204 11428 16232
rect 10336 16164 10364 16204
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 12434 16232 12440 16244
rect 11572 16204 12440 16232
rect 11572 16192 11578 16204
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 15194 16232 15200 16244
rect 15155 16204 15200 16232
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 16301 16235 16359 16241
rect 16301 16201 16313 16235
rect 16347 16232 16359 16235
rect 16666 16232 16672 16244
rect 16347 16204 16672 16232
rect 16347 16201 16359 16204
rect 16301 16195 16359 16201
rect 16666 16192 16672 16204
rect 16724 16232 16730 16244
rect 17034 16232 17040 16244
rect 16724 16204 17040 16232
rect 16724 16192 16730 16204
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17678 16232 17684 16244
rect 17543 16204 17684 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 22649 16235 22707 16241
rect 22649 16232 22661 16235
rect 20404 16204 22661 16232
rect 20404 16192 20410 16204
rect 22649 16201 22661 16204
rect 22695 16201 22707 16235
rect 22649 16195 22707 16201
rect 8588 16136 10364 16164
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 4798 16096 4804 16108
rect 1627 16068 4804 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 7098 16096 7104 16108
rect 4948 16068 7104 16096
rect 4948 16056 4954 16068
rect 7098 16056 7104 16068
rect 7156 16096 7162 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 7156 16068 7297 16096
rect 7156 16056 7162 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7650 16056 7656 16108
rect 7708 16096 7714 16108
rect 8588 16105 8616 16136
rect 10410 16124 10416 16176
rect 10468 16164 10474 16176
rect 10468 16136 11468 16164
rect 10468 16124 10474 16136
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7708 16068 7757 16096
rect 7708 16056 7714 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 9858 16096 9864 16108
rect 9819 16068 9864 16096
rect 8573 16059 8631 16065
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10284 16068 10333 16096
rect 10284 16056 10290 16068
rect 10321 16065 10333 16068
rect 10367 16096 10379 16099
rect 10778 16096 10784 16108
rect 10367 16068 10784 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11330 16096 11336 16108
rect 11195 16068 11336 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 11440 16096 11468 16136
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12802 16164 12808 16176
rect 11848 16136 12808 16164
rect 11848 16124 11854 16136
rect 12802 16124 12808 16136
rect 12860 16124 12866 16176
rect 16942 16124 16948 16176
rect 17000 16164 17006 16176
rect 19153 16167 19211 16173
rect 19153 16164 19165 16167
rect 17000 16136 19165 16164
rect 17000 16124 17006 16136
rect 19153 16133 19165 16136
rect 19199 16133 19211 16167
rect 19153 16127 19211 16133
rect 19245 16167 19303 16173
rect 19245 16133 19257 16167
rect 19291 16164 19303 16167
rect 19426 16164 19432 16176
rect 19291 16136 19432 16164
rect 19291 16133 19303 16136
rect 19245 16127 19303 16133
rect 19426 16124 19432 16136
rect 19484 16124 19490 16176
rect 20898 16164 20904 16176
rect 20859 16136 20904 16164
rect 20898 16124 20904 16136
rect 20956 16124 20962 16176
rect 21453 16167 21511 16173
rect 21453 16133 21465 16167
rect 21499 16164 21511 16167
rect 24854 16164 24860 16176
rect 21499 16136 24860 16164
rect 21499 16133 21511 16136
rect 21453 16127 21511 16133
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 11440 16068 15853 16096
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 16632 16068 18153 16096
rect 16632 16056 16638 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9766 16028 9772 16040
rect 9079 16000 9772 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 11606 16028 11612 16040
rect 10652 16000 11612 16028
rect 10652 15988 10658 16000
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 11790 15988 11796 16040
rect 11848 16028 11854 16040
rect 11885 16031 11943 16037
rect 11885 16028 11897 16031
rect 11848 16000 11897 16028
rect 11848 15988 11854 16000
rect 11885 15997 11897 16000
rect 11931 15997 11943 16031
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11885 15991 11943 15997
rect 11992 16000 12081 16028
rect 8018 15920 8024 15972
rect 8076 15960 8082 15972
rect 9858 15960 9864 15972
rect 8076 15932 9864 15960
rect 8076 15920 8082 15932
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 10410 15960 10416 15972
rect 10371 15932 10416 15960
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 11054 15920 11060 15972
rect 11112 15960 11118 15972
rect 11992 15960 12020 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12986 16028 12992 16040
rect 12947 16000 12992 16028
rect 12069 15991 12127 15997
rect 12986 15988 12992 16000
rect 13044 15988 13050 16040
rect 13170 16028 13176 16040
rect 13131 16000 13176 16028
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 14182 15988 14188 16040
rect 14240 16028 14246 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 14240 16000 14565 16028
rect 14240 15988 14246 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 14737 16031 14795 16037
rect 14737 16028 14749 16031
rect 14700 16000 14749 16028
rect 14700 15988 14706 16000
rect 14737 15997 14749 16000
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15436 16000 15669 16028
rect 15436 15988 15442 16000
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 15997 16911 16031
rect 17034 16028 17040 16040
rect 16995 16000 17040 16028
rect 16853 15991 16911 15997
rect 11112 15932 12020 15960
rect 11112 15920 11118 15932
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13357 15963 13415 15969
rect 13357 15960 13369 15963
rect 12676 15932 13369 15960
rect 12676 15920 12682 15932
rect 13357 15929 13369 15932
rect 13403 15929 13415 15963
rect 16868 15960 16896 15991
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 18782 16028 18788 16040
rect 18003 16000 18788 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 18782 15988 18788 16000
rect 18840 16028 18846 16040
rect 19978 16028 19984 16040
rect 18840 16000 19984 16028
rect 18840 15988 18846 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 16028 20867 16031
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 20855 16000 22017 16028
rect 20855 15997 20867 16000
rect 20809 15991 20867 15997
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 17494 15960 17500 15972
rect 16868 15932 17500 15960
rect 13357 15923 13415 15929
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 18046 15920 18052 15972
rect 18104 15960 18110 15972
rect 18325 15963 18383 15969
rect 18325 15960 18337 15963
rect 18104 15932 18337 15960
rect 18104 15920 18110 15932
rect 18325 15929 18337 15932
rect 18371 15929 18383 15963
rect 18325 15923 18383 15929
rect 19705 15963 19763 15969
rect 19705 15929 19717 15963
rect 19751 15929 19763 15963
rect 22112 15960 22140 16136
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 22830 16096 22836 16108
rect 22791 16068 22836 16096
rect 22830 16056 22836 16068
rect 22888 16056 22894 16108
rect 24118 16096 24124 16108
rect 24079 16068 24124 16096
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 38286 16096 38292 16108
rect 38247 16068 38292 16096
rect 38286 16056 38292 16068
rect 38344 16056 38350 16108
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 23164 16000 23305 16028
rect 23164 15988 23170 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 24026 15988 24032 16040
rect 24084 16028 24090 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24084 16000 24593 16028
rect 24084 15988 24090 16000
rect 24581 15997 24593 16000
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 19705 15923 19763 15929
rect 21468 15932 22140 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 7834 15892 7840 15904
rect 7795 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 10502 15892 10508 15904
rect 10192 15864 10508 15892
rect 10192 15852 10198 15864
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10928 15864 10977 15892
rect 10928 15852 10934 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 11974 15892 11980 15904
rect 11848 15864 11980 15892
rect 11848 15852 11854 15864
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12526 15892 12532 15904
rect 12487 15864 12532 15892
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 19720 15892 19748 15923
rect 21468 15892 21496 15932
rect 19720 15864 21496 15892
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 22186 15892 22192 15904
rect 21600 15864 22192 15892
rect 21600 15852 21606 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 23937 15895 23995 15901
rect 23937 15892 23949 15895
rect 23348 15864 23949 15892
rect 23348 15852 23354 15864
rect 23937 15861 23949 15864
rect 23983 15861 23995 15895
rect 23937 15855 23995 15861
rect 36998 15852 37004 15904
rect 37056 15892 37062 15904
rect 38105 15895 38163 15901
rect 38105 15892 38117 15895
rect 37056 15864 38117 15892
rect 37056 15852 37062 15864
rect 38105 15861 38117 15864
rect 38151 15861 38163 15895
rect 38105 15855 38163 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 8352 15660 8401 15688
rect 8352 15648 8358 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 8389 15651 8447 15657
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 13170 15688 13176 15700
rect 9640 15660 13176 15688
rect 9640 15648 9646 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 16666 15688 16672 15700
rect 14240 15660 16068 15688
rect 16627 15660 16672 15688
rect 14240 15648 14246 15660
rect 7834 15580 7840 15632
rect 7892 15620 7898 15632
rect 7892 15592 11928 15620
rect 7892 15580 7898 15592
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15552 7435 15555
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 7423 15524 10609 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 11514 15552 11520 15564
rect 10744 15524 11520 15552
rect 10744 15512 10750 15524
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 11900 15561 11928 15592
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 12069 15623 12127 15629
rect 12069 15620 12081 15623
rect 12032 15592 12081 15620
rect 12032 15580 12038 15592
rect 12069 15589 12081 15592
rect 12115 15620 12127 15623
rect 12710 15620 12716 15632
rect 12115 15592 12716 15620
rect 12115 15589 12127 15592
rect 12069 15583 12127 15589
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 14274 15620 14280 15632
rect 12912 15592 14280 15620
rect 12912 15561 12940 15592
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 14366 15580 14372 15632
rect 14424 15620 14430 15632
rect 15930 15620 15936 15632
rect 14424 15592 15936 15620
rect 14424 15580 14430 15592
rect 15930 15580 15936 15592
rect 15988 15580 15994 15632
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15521 11943 15555
rect 11885 15515 11943 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15521 12955 15555
rect 12897 15515 12955 15521
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 13136 15524 13185 15552
rect 13136 15512 13142 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 16040 15561 16068 15660
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 18966 15688 18972 15700
rect 18739 15660 18972 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 24118 15648 24124 15700
rect 24176 15688 24182 15700
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 24176 15660 24593 15688
rect 24176 15648 24182 15660
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 33318 15620 33324 15632
rect 17552 15592 20024 15620
rect 17552 15580 17558 15592
rect 14645 15555 14703 15561
rect 14645 15552 14657 15555
rect 13964 15524 14657 15552
rect 13964 15512 13970 15524
rect 14645 15521 14657 15524
rect 14691 15521 14703 15555
rect 14645 15515 14703 15521
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15552 17371 15555
rect 19334 15552 19340 15564
rect 17359 15524 19340 15552
rect 17359 15521 17371 15524
rect 17313 15515 17371 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19996 15561 20024 15592
rect 22066 15592 33324 15620
rect 19981 15555 20039 15561
rect 19981 15521 19993 15555
rect 20027 15521 20039 15555
rect 19981 15515 20039 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15552 21695 15555
rect 22066 15552 22094 15592
rect 33318 15580 33324 15592
rect 33376 15580 33382 15632
rect 23106 15552 23112 15564
rect 21683 15524 22094 15552
rect 23067 15524 23112 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23290 15552 23296 15564
rect 23251 15524 23296 15552
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 5592 15456 7297 15484
rect 5592 15444 5598 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8260 15456 8585 15484
rect 8260 15444 8266 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 8573 15447 8631 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15453 9367 15487
rect 9674 15484 9680 15496
rect 9309 15447 9367 15453
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 9325 15416 9353 15447
rect 7248 15388 9353 15416
rect 9646 15444 9680 15484
rect 9732 15444 9738 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 9916 15456 10793 15484
rect 9916 15444 9922 15456
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11701 15487 11759 15493
rect 11701 15484 11713 15487
rect 11204 15456 11713 15484
rect 11204 15444 11210 15456
rect 11701 15453 11713 15456
rect 11747 15484 11759 15487
rect 12066 15484 12072 15496
rect 11747 15456 12072 15484
rect 11747 15453 11759 15456
rect 11701 15447 11759 15453
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 16206 15484 16212 15496
rect 16167 15456 16212 15484
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 18874 15484 18880 15496
rect 18835 15456 18880 15484
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 21821 15487 21879 15493
rect 21821 15453 21833 15487
rect 21867 15484 21879 15487
rect 22094 15484 22100 15496
rect 21867 15456 22100 15484
rect 21867 15453 21879 15456
rect 21821 15447 21879 15453
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 25130 15484 25136 15496
rect 24811 15456 25136 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 25130 15444 25136 15456
rect 25188 15444 25194 15496
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 7248 15376 7254 15388
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 9646 15348 9674 15444
rect 9784 15416 9812 15444
rect 11241 15419 11299 15425
rect 9784 15388 9904 15416
rect 9766 15348 9772 15360
rect 9180 15320 9674 15348
rect 9727 15320 9772 15348
rect 9180 15308 9186 15320
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 9876 15348 9904 15388
rect 11241 15385 11253 15419
rect 11287 15416 11299 15419
rect 12526 15416 12532 15428
rect 11287 15388 12532 15416
rect 11287 15385 11299 15388
rect 11241 15379 11299 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 12982 15419 13040 15425
rect 12982 15385 12994 15419
rect 13028 15385 13040 15419
rect 14366 15416 14372 15428
rect 14327 15388 14372 15416
rect 12982 15379 13040 15385
rect 11514 15348 11520 15360
rect 9876 15320 11520 15348
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 13004 15348 13032 15379
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 14461 15419 14519 15425
rect 14461 15385 14473 15419
rect 14507 15385 14519 15419
rect 14461 15379 14519 15385
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15385 17463 15419
rect 17405 15379 17463 15385
rect 12216 15320 13032 15348
rect 12216 15308 12222 15320
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 14476 15348 14504 15379
rect 13780 15320 14504 15348
rect 13780 15308 13786 15320
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 17420 15348 17448 15379
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 17957 15419 18015 15425
rect 17957 15416 17969 15419
rect 17644 15388 17969 15416
rect 17644 15376 17650 15388
rect 17957 15385 17969 15388
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 17000 15320 17448 15348
rect 20625 15351 20683 15357
rect 17000 15308 17006 15320
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 20671 15320 22293 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 22281 15317 22293 15320
rect 22327 15348 22339 15351
rect 22554 15348 22560 15360
rect 22327 15320 22560 15348
rect 22327 15317 22339 15320
rect 22281 15311 22339 15317
rect 22554 15308 22560 15320
rect 22612 15308 22618 15360
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 23753 15351 23811 15357
rect 23753 15348 23765 15351
rect 23624 15320 23765 15348
rect 23624 15308 23630 15320
rect 23753 15317 23765 15320
rect 23799 15317 23811 15351
rect 23753 15311 23811 15317
rect 24854 15308 24860 15360
rect 24912 15348 24918 15360
rect 25225 15351 25283 15357
rect 25225 15348 25237 15351
rect 24912 15320 25237 15348
rect 24912 15308 24918 15320
rect 25225 15317 25237 15320
rect 25271 15317 25283 15351
rect 25225 15311 25283 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 9766 15144 9772 15156
rect 7024 15116 9772 15144
rect 7024 15017 7052 15116
rect 9766 15104 9772 15116
rect 9824 15144 9830 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 9824 15116 10885 15144
rect 9824 15104 9830 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 10873 15107 10931 15113
rect 11793 15147 11851 15153
rect 11793 15113 11805 15147
rect 11839 15144 11851 15147
rect 12342 15144 12348 15156
rect 11839 15116 12348 15144
rect 11839 15113 11851 15116
rect 11793 15107 11851 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 15565 15147 15623 15153
rect 12860 15116 15516 15144
rect 12860 15104 12866 15116
rect 9033 15079 9091 15085
rect 7852 15048 8984 15076
rect 7852 15017 7880 15048
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7009 14971 7067 14977
rect 7116 14980 7849 15008
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 7116 14940 7144 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 8956 15017 8984 15048
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 11054 15076 11060 15088
rect 9079 15048 11060 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 11514 15036 11520 15088
rect 11572 15076 11578 15088
rect 15378 15076 15384 15088
rect 11572 15048 12388 15076
rect 11572 15036 11578 15048
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 8168 14980 8493 15008
rect 8168 14968 8174 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9732 14980 9781 15008
rect 9732 14968 9738 14980
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 9769 14971 9827 14977
rect 9876 14980 10425 15008
rect 3200 14912 7144 14940
rect 3200 14900 3206 14912
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 9876 14940 9904 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11664 14980 11713 15008
rect 11664 14968 11670 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 12360 15017 12388 15048
rect 13924 15048 15384 15076
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 7800 14912 9904 14940
rect 10229 14943 10287 14949
rect 7800 14900 7806 14912
rect 10229 14909 10241 14943
rect 10275 14940 10287 14943
rect 11992 14940 12020 14968
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 10275 14912 12020 14940
rect 12452 14928 12541 14940
rect 12406 14912 12541 14928
rect 10275 14909 10287 14912
rect 10229 14903 10287 14909
rect 12406 14900 12480 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13924 14949 13952 15048
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 15488 15076 15516 15116
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 16574 15144 16580 15156
rect 15611 15116 16580 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 18874 15144 18880 15156
rect 18835 15116 18880 15144
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 19392 15116 20177 15144
rect 19392 15104 19398 15116
rect 20165 15113 20177 15116
rect 20211 15144 20223 15147
rect 20346 15144 20352 15156
rect 20211 15116 20352 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 20898 15144 20904 15156
rect 20671 15116 20904 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22152 15116 22197 15144
rect 22152 15104 22158 15116
rect 25406 15104 25412 15156
rect 25464 15144 25470 15156
rect 25777 15147 25835 15153
rect 25777 15144 25789 15147
rect 25464 15116 25789 15144
rect 25464 15104 25470 15116
rect 25777 15113 25789 15116
rect 25823 15113 25835 15147
rect 25777 15107 25835 15113
rect 17497 15079 17555 15085
rect 17497 15076 17509 15079
rect 15488 15048 17509 15076
rect 17497 15045 17509 15048
rect 17543 15045 17555 15079
rect 17497 15039 17555 15045
rect 17589 15079 17647 15085
rect 17589 15045 17601 15079
rect 17635 15076 17647 15079
rect 18782 15076 18788 15088
rect 17635 15048 18788 15076
rect 17635 15045 17647 15048
rect 17589 15039 17647 15045
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 20714 15076 20720 15088
rect 18984 15048 20720 15076
rect 14550 15008 14556 15020
rect 14016 14980 14556 15008
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13688 14912 13921 14940
rect 13688 14900 13694 14912
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 7653 14875 7711 14881
rect 7653 14841 7665 14875
rect 7699 14872 7711 14875
rect 9214 14872 9220 14884
rect 7699 14844 9220 14872
rect 7699 14841 7711 14844
rect 7653 14835 7711 14841
rect 9214 14832 9220 14844
rect 9272 14832 9278 14884
rect 9582 14872 9588 14884
rect 9543 14844 9588 14872
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 12406 14872 12434 14900
rect 12710 14872 12716 14884
rect 12268 14844 12434 14872
rect 12671 14844 12716 14872
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 7101 14807 7159 14813
rect 7101 14804 7113 14807
rect 5040 14776 7113 14804
rect 5040 14764 5046 14776
rect 7101 14773 7113 14776
rect 7147 14773 7159 14807
rect 8294 14804 8300 14816
rect 8255 14776 8300 14804
rect 7101 14767 7159 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 12268 14804 12296 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 14016 14872 14044 14980
rect 14550 14968 14556 14980
rect 14608 15008 14614 15020
rect 15470 15008 15476 15020
rect 14608 14980 15332 15008
rect 15431 14980 15476 15008
rect 14608 14968 14614 14980
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 13504 14844 14044 14872
rect 13504 14832 13510 14844
rect 8444 14776 12296 14804
rect 8444 14764 8450 14776
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 14108 14804 14136 14903
rect 14274 14872 14280 14884
rect 14235 14844 14280 14872
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 15304 14872 15332 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 15008 18199 15011
rect 18984 15008 19012 15048
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 18187 14980 19012 15008
rect 19061 15011 19119 15017
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 20806 15008 20812 15020
rect 19107 14980 20668 15008
rect 20767 14980 20812 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 16022 14940 16028 14952
rect 15436 14912 16028 14940
rect 15436 14900 15442 14912
rect 16022 14900 16028 14912
rect 16080 14940 16086 14952
rect 16316 14940 16344 14971
rect 18414 14940 18420 14952
rect 16080 14912 18420 14940
rect 16080 14900 16086 14912
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 19076 14940 19104 14971
rect 18984 14912 19104 14940
rect 19521 14943 19579 14949
rect 18984 14872 19012 14912
rect 19521 14909 19533 14943
rect 19567 14940 19579 14943
rect 19610 14940 19616 14952
rect 19567 14912 19616 14940
rect 19567 14909 19579 14912
rect 19521 14903 19579 14909
rect 19610 14900 19616 14912
rect 19668 14900 19674 14952
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14909 19763 14943
rect 20640 14940 20668 14980
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 21453 15011 21511 15017
rect 21453 15008 21465 15011
rect 20956 14980 21465 15008
rect 20956 14968 20962 14980
rect 21453 14977 21465 14980
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 24026 15008 24032 15020
rect 23987 14980 24032 15008
rect 22005 14971 22063 14977
rect 20990 14940 20996 14952
rect 20640 14912 20996 14940
rect 19705 14903 19763 14909
rect 15304 14844 19012 14872
rect 19720 14872 19748 14903
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21174 14900 21180 14952
rect 21232 14940 21238 14952
rect 22020 14940 22048 14971
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24854 15008 24860 15020
rect 24259 14980 24860 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24854 14968 24860 14980
rect 24912 14968 24918 15020
rect 25130 15008 25136 15020
rect 25091 14980 25136 15008
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 15008 26019 15011
rect 26050 15008 26056 15020
rect 26007 14980 26056 15008
rect 26007 14977 26019 14980
rect 25961 14971 26019 14977
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 33045 15011 33103 15017
rect 33045 14977 33057 15011
rect 33091 15008 33103 15011
rect 36998 15008 37004 15020
rect 33091 14980 37004 15008
rect 33091 14977 33103 14980
rect 33045 14971 33103 14977
rect 36998 14968 37004 14980
rect 37056 14968 37062 15020
rect 21232 14912 22048 14940
rect 22925 14943 22983 14949
rect 21232 14900 21238 14912
rect 22925 14909 22937 14943
rect 22971 14909 22983 14943
rect 22925 14903 22983 14909
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14940 23167 14943
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 23155 14912 25237 14940
rect 23155 14909 23167 14912
rect 23109 14903 23167 14909
rect 25225 14909 25237 14912
rect 25271 14909 25283 14943
rect 25225 14903 25283 14909
rect 21269 14875 21327 14881
rect 21269 14872 21281 14875
rect 19720 14844 21281 14872
rect 21269 14841 21281 14844
rect 21315 14841 21327 14875
rect 22940 14872 22968 14903
rect 22940 14844 24624 14872
rect 21269 14835 21327 14841
rect 24596 14816 24624 14844
rect 12400 14776 14136 14804
rect 16117 14807 16175 14813
rect 12400 14764 12406 14776
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 17402 14804 17408 14816
rect 16163 14776 17408 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 23566 14804 23572 14816
rect 23527 14776 23572 14804
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 24394 14804 24400 14816
rect 24355 14776 24400 14804
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 29362 14804 29368 14816
rect 24636 14776 29368 14804
rect 24636 14764 24642 14776
rect 29362 14764 29368 14776
rect 29420 14764 29426 14816
rect 33134 14804 33140 14816
rect 33095 14776 33140 14804
rect 33134 14764 33140 14776
rect 33192 14764 33198 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 4798 14600 4804 14612
rect 4759 14572 4804 14600
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 8110 14600 8116 14612
rect 6420 14572 8116 14600
rect 6420 14560 6426 14572
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 11238 14600 11244 14612
rect 8527 14572 11244 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 12250 14600 12256 14612
rect 11532 14572 12256 14600
rect 1581 14535 1639 14541
rect 1581 14501 1593 14535
rect 1627 14532 1639 14535
rect 6546 14532 6552 14544
rect 1627 14504 6552 14532
rect 1627 14501 1639 14504
rect 1581 14495 1639 14501
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 10229 14535 10287 14541
rect 10229 14501 10241 14535
rect 10275 14532 10287 14535
rect 10594 14532 10600 14544
rect 10275 14504 10600 14532
rect 10275 14501 10287 14504
rect 10229 14495 10287 14501
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 10778 14492 10784 14544
rect 10836 14532 10842 14544
rect 11532 14532 11560 14572
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12345 14603 12403 14609
rect 12345 14569 12357 14603
rect 12391 14600 12403 14603
rect 12894 14600 12900 14612
rect 12391 14572 12900 14600
rect 12391 14569 12403 14572
rect 12345 14563 12403 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 13412 14572 13553 14600
rect 13412 14560 13418 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 13541 14563 13599 14569
rect 14737 14603 14795 14609
rect 14737 14569 14749 14603
rect 14783 14600 14795 14603
rect 15286 14600 15292 14612
rect 14783 14572 15292 14600
rect 14783 14569 14795 14572
rect 14737 14563 14795 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 16574 14600 16580 14612
rect 15396 14572 16580 14600
rect 10836 14504 11560 14532
rect 11609 14535 11667 14541
rect 10836 14492 10842 14504
rect 11609 14501 11621 14535
rect 11655 14532 11667 14535
rect 13814 14532 13820 14544
rect 11655 14504 13820 14532
rect 11655 14501 11667 14504
rect 11609 14495 11667 14501
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 15396 14532 15424 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14600 16727 14603
rect 17034 14600 17040 14612
rect 16715 14572 17040 14600
rect 16715 14569 16727 14572
rect 16669 14563 16727 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17221 14603 17279 14609
rect 17221 14569 17233 14603
rect 17267 14600 17279 14603
rect 17770 14600 17776 14612
rect 17267 14572 17776 14600
rect 17267 14569 17279 14572
rect 17221 14563 17279 14569
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18322 14600 18328 14612
rect 18187 14572 18328 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 20070 14600 20076 14612
rect 18739 14572 20076 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 20349 14603 20407 14609
rect 20349 14600 20361 14603
rect 20220 14572 20361 14600
rect 20220 14560 20226 14572
rect 20349 14569 20361 14572
rect 20395 14569 20407 14603
rect 20349 14563 20407 14569
rect 24394 14560 24400 14612
rect 24452 14600 24458 14612
rect 24949 14603 25007 14609
rect 24949 14600 24961 14603
rect 24452 14572 24961 14600
rect 24452 14560 24458 14572
rect 24949 14569 24961 14572
rect 24995 14569 25007 14603
rect 24949 14563 25007 14569
rect 25866 14560 25872 14612
rect 25924 14600 25930 14612
rect 25924 14572 31754 14600
rect 25924 14560 25930 14572
rect 13924 14504 15424 14532
rect 16025 14535 16083 14541
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 9769 14467 9827 14473
rect 9769 14464 9781 14467
rect 7883 14436 9781 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 9769 14433 9781 14436
rect 9815 14433 9827 14467
rect 9769 14427 9827 14433
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 12894 14464 12900 14476
rect 11011 14436 12900 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13924 14464 13952 14504
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 17126 14532 17132 14544
rect 16071 14504 17132 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 17126 14492 17132 14504
rect 17184 14492 17190 14544
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14501 21051 14535
rect 20993 14495 21051 14501
rect 13004 14436 13952 14464
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 2774 14396 2780 14408
rect 2363 14368 2780 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 4982 14396 4988 14408
rect 4943 14368 4988 14396
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 7745 14359 7803 14365
rect 7760 14328 7788 14359
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9585 14399 9643 14405
rect 9585 14396 9597 14399
rect 8536 14368 9597 14396
rect 8536 14356 8542 14368
rect 9585 14365 9597 14368
rect 9631 14365 9643 14399
rect 11790 14396 11796 14408
rect 11751 14368 11796 14396
rect 9585 14359 9643 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12124 14368 12265 14396
rect 12124 14356 12130 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 13004 14396 13032 14436
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 15562 14464 15568 14476
rect 14516 14436 15568 14464
rect 14516 14424 14522 14436
rect 15562 14424 15568 14436
rect 15620 14464 15626 14476
rect 19610 14464 19616 14476
rect 15620 14436 16620 14464
rect 19571 14436 19616 14464
rect 15620 14424 15626 14436
rect 12492 14368 13032 14396
rect 13081 14399 13139 14405
rect 12492 14356 12498 14368
rect 13081 14365 13093 14399
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 9950 14328 9956 14340
rect 7760 14300 9956 14328
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 13096 14328 13124 14359
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13228 14368 13737 14396
rect 13228 14356 13234 14368
rect 13725 14365 13737 14368
rect 13771 14396 13783 14399
rect 14274 14396 14280 14408
rect 13771 14368 14280 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14642 14396 14648 14408
rect 14603 14368 14648 14396
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16592 14405 16620 14436
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 17402 14396 17408 14408
rect 17363 14368 17408 14396
rect 16577 14359 16635 14365
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 18046 14396 18052 14408
rect 18007 14368 18052 14396
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18472 14368 18889 14396
rect 18472 14356 18478 14368
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14396 20591 14399
rect 21008 14396 21036 14495
rect 22462 14492 22468 14544
rect 22520 14532 22526 14544
rect 23201 14535 23259 14541
rect 23201 14532 23213 14535
rect 22520 14504 23213 14532
rect 22520 14492 22526 14504
rect 23201 14501 23213 14504
rect 23247 14501 23259 14535
rect 23201 14495 23259 14501
rect 24210 14492 24216 14544
rect 24268 14532 24274 14544
rect 26329 14535 26387 14541
rect 26329 14532 26341 14535
rect 24268 14504 26341 14532
rect 24268 14492 24274 14504
rect 26329 14501 26341 14504
rect 26375 14501 26387 14535
rect 26329 14495 26387 14501
rect 22833 14467 22891 14473
rect 22833 14433 22845 14467
rect 22879 14464 22891 14467
rect 24578 14464 24584 14476
rect 22879 14436 24584 14464
rect 22879 14433 22891 14436
rect 22833 14427 22891 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 24765 14467 24823 14473
rect 24765 14433 24777 14467
rect 24811 14464 24823 14467
rect 27065 14467 27123 14473
rect 27065 14464 27077 14467
rect 24811 14436 27077 14464
rect 24811 14433 24823 14436
rect 24765 14427 24823 14433
rect 27065 14433 27077 14436
rect 27111 14433 27123 14467
rect 27065 14427 27123 14433
rect 21174 14396 21180 14408
rect 20579 14368 21036 14396
rect 21135 14368 21180 14396
rect 20579 14365 20591 14368
rect 20533 14359 20591 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 21266 14356 21272 14408
rect 21324 14396 21330 14408
rect 22005 14399 22063 14405
rect 22005 14396 22017 14399
rect 21324 14368 22017 14396
rect 21324 14356 21330 14368
rect 22005 14365 22017 14368
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14396 23075 14399
rect 24486 14396 24492 14408
rect 23063 14368 24492 14396
rect 23063 14365 23075 14368
rect 23017 14359 23075 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 25866 14396 25872 14408
rect 25827 14368 25872 14396
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 26513 14399 26571 14405
rect 26513 14365 26525 14399
rect 26559 14365 26571 14399
rect 26513 14359 26571 14365
rect 26973 14399 27031 14405
rect 26973 14365 26985 14399
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 26528 14328 26556 14359
rect 12728 14300 13124 14328
rect 25700 14300 26556 14328
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 2590 14260 2596 14272
rect 2455 14232 2596 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2590 14220 2596 14232
rect 2648 14220 2654 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 12066 14260 12072 14272
rect 9088 14232 12072 14260
rect 9088 14220 9094 14232
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12250 14220 12256 14272
rect 12308 14260 12314 14272
rect 12728 14260 12756 14300
rect 12308 14232 12756 14260
rect 12897 14263 12955 14269
rect 12308 14220 12314 14232
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 13998 14260 14004 14272
rect 12943 14232 14004 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 14792 14232 15301 14260
rect 14792 14220 14798 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 15289 14223 15347 14229
rect 21821 14263 21879 14269
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 22186 14260 22192 14272
rect 21867 14232 22192 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 25700 14269 25728 14300
rect 25685 14263 25743 14269
rect 25685 14229 25697 14263
rect 25731 14229 25743 14263
rect 25685 14223 25743 14229
rect 26050 14220 26056 14272
rect 26108 14260 26114 14272
rect 26988 14260 27016 14359
rect 31726 14328 31754 14572
rect 36446 14356 36452 14408
rect 36504 14396 36510 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 36504 14368 38025 14396
rect 36504 14356 36510 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 37826 14328 37832 14340
rect 31726 14300 37832 14328
rect 37826 14288 37832 14300
rect 37884 14288 37890 14340
rect 38194 14260 38200 14272
rect 26108 14232 27016 14260
rect 38155 14232 38200 14260
rect 26108 14220 26114 14232
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9490 14056 9496 14068
rect 9079 14028 9496 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 10686 14056 10692 14068
rect 10367 14028 10692 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 11103 14028 13308 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 5534 13988 5540 14000
rect 2976 13960 5540 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2774 13920 2780 13932
rect 2271 13892 2780 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 2976 13929 3004 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 8481 13991 8539 13997
rect 8481 13957 8493 13991
rect 8527 13988 8539 13991
rect 8527 13960 12020 13988
rect 8527 13957 8539 13960
rect 8481 13951 8539 13957
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 3602 13920 3608 13932
rect 3563 13892 3608 13920
rect 2961 13883 3019 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7374 13920 7380 13932
rect 7147 13892 7380 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7926 13920 7932 13932
rect 7887 13892 7932 13920
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8202 13920 8208 13932
rect 8115 13892 8208 13920
rect 8202 13880 8208 13892
rect 8260 13920 8266 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8260 13892 8401 13920
rect 8260 13880 8266 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 8389 13883 8447 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 9950 13920 9956 13932
rect 9907 13892 9956 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10226 13920 10232 13932
rect 10008 13892 10232 13920
rect 10008 13880 10014 13892
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10410 13920 10416 13932
rect 10284 13892 10416 13920
rect 10284 13880 10290 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 2314 13852 2320 13864
rect 2275 13824 2320 13852
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 5626 13852 5632 13864
rect 3743 13824 5632 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8220 13852 8248 13880
rect 7892 13824 8248 13852
rect 7892 13812 7898 13824
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 10520 13852 10548 13883
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 11992 13929 12020 13960
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 13280 13988 13308 14028
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14001 14059 14059 14065
rect 13412 14028 13457 14056
rect 13412 14016 13418 14028
rect 14001 14025 14013 14059
rect 14047 14056 14059 14059
rect 14737 14059 14795 14065
rect 14047 14028 14504 14056
rect 14047 14025 14059 14028
rect 14001 14019 14059 14025
rect 13722 13988 13728 14000
rect 12492 13960 12537 13988
rect 13280 13960 13728 13988
rect 12492 13948 12498 13960
rect 13722 13948 13728 13960
rect 13780 13948 13786 14000
rect 14476 13988 14504 14028
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 16206 14056 16212 14068
rect 14783 14028 16212 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 18414 14056 18420 14068
rect 18375 14028 18420 14056
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20898 14056 20904 14068
rect 20119 14028 20904 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 25869 14059 25927 14065
rect 22066 14028 25452 14056
rect 22066 14000 22094 14028
rect 15010 13988 15016 14000
rect 14476 13960 15016 13988
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 21082 13988 21088 14000
rect 15212 13960 21088 13988
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10652 13892 10977 13920
rect 10652 13880 10658 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12952 13892 13553 13920
rect 12952 13880 12958 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14056 13892 14197 13920
rect 14056 13880 14062 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 14332 13892 14657 13920
rect 14332 13880 14338 13892
rect 14645 13889 14657 13892
rect 14691 13920 14703 13923
rect 15212 13920 15240 13960
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 22002 13948 22008 14000
rect 22060 13960 22094 14000
rect 24210 13988 24216 14000
rect 24171 13960 24216 13988
rect 22060 13948 22066 13960
rect 24210 13948 24216 13960
rect 24268 13948 24274 14000
rect 17586 13920 17592 13932
rect 14691 13892 15240 13920
rect 15304 13892 17592 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 15304 13861 15332 13892
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18104 13892 18613 13920
rect 18104 13880 18110 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 19426 13920 19432 13932
rect 19387 13892 19432 13920
rect 18601 13883 18659 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 20254 13920 20260 13932
rect 20167 13892 20260 13920
rect 20254 13880 20260 13892
rect 20312 13920 20318 13932
rect 20622 13920 20628 13932
rect 20312 13892 20628 13920
rect 20312 13880 20318 13892
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21450 13920 21456 13932
rect 21411 13892 21456 13920
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 22186 13920 22192 13932
rect 22147 13892 22192 13920
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 25424 13929 25452 14028
rect 25869 14025 25881 14059
rect 25915 14056 25927 14059
rect 26602 14056 26608 14068
rect 25915 14028 26608 14056
rect 25915 14025 25927 14028
rect 25869 14019 25927 14025
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 25556 13892 26065 13920
rect 25556 13880 25562 13892
rect 26053 13889 26065 13892
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 8352 13824 10548 13852
rect 10612 13824 11805 13852
rect 8352 13812 8358 13824
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 10612 13784 10640 13824
rect 11793 13821 11805 13824
rect 11839 13852 11851 13855
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 11839 13824 15301 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 15289 13821 15301 13824
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15436 13824 15485 13852
rect 15436 13812 15442 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15896 13824 15945 13852
rect 15896 13812 15902 13824
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 17034 13852 17040 13864
rect 16995 13824 17040 13852
rect 15933 13815 15991 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17218 13852 17224 13864
rect 17179 13824 17224 13852
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 18012 13824 22017 13852
rect 18012 13812 18018 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 23106 13852 23112 13864
rect 23067 13824 23112 13852
rect 22005 13815 22063 13821
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24394 13852 24400 13864
rect 24167 13824 24400 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24762 13852 24768 13864
rect 24723 13824 24768 13852
rect 24762 13812 24768 13824
rect 24820 13812 24826 13864
rect 9364 13756 10640 13784
rect 9364 13744 9370 13756
rect 10870 13744 10876 13796
rect 10928 13784 10934 13796
rect 17126 13784 17132 13796
rect 10928 13756 17132 13784
rect 10928 13744 10934 13756
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 23198 13744 23204 13796
rect 23256 13784 23262 13796
rect 33134 13784 33140 13796
rect 23256 13756 33140 13784
rect 23256 13744 23262 13756
rect 33134 13744 33140 13756
rect 33192 13744 33198 13796
rect 1673 13719 1731 13725
rect 1673 13685 1685 13719
rect 1719 13716 1731 13719
rect 2222 13716 2228 13728
rect 1719 13688 2228 13716
rect 1719 13685 1731 13688
rect 1673 13679 1731 13685
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 10962 13716 10968 13728
rect 6420 13688 10968 13716
rect 6420 13676 6426 13688
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12802 13716 12808 13728
rect 11664 13688 12808 13716
rect 11664 13676 11670 13688
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 22646 13716 22652 13728
rect 22607 13688 22652 13716
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 23014 13676 23020 13728
rect 23072 13716 23078 13728
rect 25225 13719 25283 13725
rect 25225 13716 25237 13719
rect 23072 13688 25237 13716
rect 23072 13676 23078 13688
rect 25225 13685 25237 13688
rect 25271 13685 25283 13719
rect 25225 13679 25283 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7926 13512 7932 13524
rect 7147 13484 7932 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 11330 13512 11336 13524
rect 8435 13484 11336 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 12253 13515 12311 13521
rect 11480 13484 11525 13512
rect 11480 13472 11486 13484
rect 12253 13481 12265 13515
rect 12299 13512 12311 13515
rect 12342 13512 12348 13524
rect 12299 13484 12348 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12989 13515 13047 13521
rect 12989 13481 13001 13515
rect 13035 13512 13047 13515
rect 13035 13484 13492 13512
rect 13035 13481 13047 13484
rect 12989 13475 13047 13481
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 5810 13444 5816 13456
rect 1627 13416 5816 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 9493 13447 9551 13453
rect 6880 13416 9076 13444
rect 6880 13404 6886 13416
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 4982 13376 4988 13388
rect 2731 13348 4988 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 9048 13376 9076 13416
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 13464 13444 13492 13484
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 19521 13515 19579 13521
rect 13780 13484 18644 13512
rect 13780 13472 13786 13484
rect 9539 13416 12940 13444
rect 13464 13416 14872 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9950 13376 9956 13388
rect 9048 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13376 10287 13379
rect 12912 13376 12940 13416
rect 14844 13376 14872 13416
rect 15838 13404 15844 13456
rect 15896 13444 15902 13456
rect 15896 13416 15941 13444
rect 16316 13416 16712 13444
rect 15896 13404 15902 13416
rect 16316 13376 16344 13416
rect 16482 13376 16488 13388
rect 10275 13348 12848 13376
rect 12912 13348 13768 13376
rect 14844 13348 16344 13376
rect 16443 13348 16488 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1452 13280 1777 13308
rect 1452 13268 1458 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13308 2651 13311
rect 2774 13308 2780 13320
rect 2639 13280 2780 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 2774 13268 2780 13280
rect 2832 13308 2838 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2832 13280 3249 13308
rect 2832 13268 2838 13280
rect 3237 13277 3249 13280
rect 3283 13308 3295 13311
rect 3602 13308 3608 13320
rect 3283 13280 3608 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3602 13268 3608 13280
rect 3660 13308 3666 13320
rect 3970 13308 3976 13320
rect 3660 13280 3976 13308
rect 3660 13268 3666 13280
rect 3970 13268 3976 13280
rect 4028 13308 4034 13320
rect 4157 13311 4215 13317
rect 4157 13308 4169 13311
rect 4028 13280 4169 13308
rect 4028 13268 4034 13280
rect 4157 13277 4169 13280
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7374 13308 7380 13320
rect 7331 13280 7380 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7800 13280 7941 13308
rect 7800 13268 7806 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9858 13308 9864 13320
rect 9723 13280 9864 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 3329 13243 3387 13249
rect 3329 13209 3341 13243
rect 3375 13240 3387 13243
rect 5074 13240 5080 13252
rect 3375 13212 5080 13240
rect 3375 13209 3387 13212
rect 3329 13203 3387 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 8588 13240 8616 13271
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 7760 13212 8616 13240
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 6638 13172 6644 13184
rect 4295 13144 6644 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7760 13181 7788 13212
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 8720 13212 9674 13240
rect 8720 13200 8726 13212
rect 7745 13175 7803 13181
rect 7745 13141 7757 13175
rect 7791 13141 7803 13175
rect 7745 13135 7803 13141
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 9490 13172 9496 13184
rect 8076 13144 9496 13172
rect 8076 13132 8082 13144
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9646 13172 9674 13212
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10152 13240 10180 13271
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10781 13311 10839 13317
rect 10781 13308 10793 13311
rect 10468 13280 10793 13308
rect 10468 13268 10474 13280
rect 10781 13277 10793 13280
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 10928 13280 11621 13308
rect 10928 13268 10934 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 12434 13308 12440 13320
rect 12395 13280 12440 13308
rect 11609 13271 11667 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 10008 13212 10180 13240
rect 12820 13240 12848 13348
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13740 13317 13768 13348
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 16684 13385 16712 13416
rect 17402 13404 17408 13456
rect 17460 13444 17466 13456
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 17460 13416 17969 13444
rect 17460 13404 17466 13416
rect 17957 13413 17969 13416
rect 18003 13413 18015 13447
rect 17957 13407 18015 13413
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13345 16727 13379
rect 17586 13376 17592 13388
rect 17547 13348 17592 13376
rect 16669 13339 16727 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 13725 13311 13783 13317
rect 12952 13280 12997 13308
rect 12952 13268 12958 13280
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13277 14887 13311
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 14829 13271 14887 13277
rect 13170 13240 13176 13252
rect 12820 13212 13176 13240
rect 10008 13200 10014 13212
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 14844 13240 14872 13271
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 17034 13308 17040 13320
rect 15856 13280 17040 13308
rect 13412 13212 14872 13240
rect 13412 13200 13418 13212
rect 15010 13200 15016 13252
rect 15068 13240 15074 13252
rect 15856 13240 15884 13280
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 15068 13212 15884 13240
rect 15068 13200 15074 13212
rect 15930 13200 15936 13252
rect 15988 13240 15994 13252
rect 17788 13240 17816 13271
rect 15988 13212 17816 13240
rect 18616 13240 18644 13484
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 20806 13512 20812 13524
rect 19567 13484 20812 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 22462 13512 22468 13524
rect 22423 13484 22468 13512
rect 22462 13472 22468 13484
rect 22520 13472 22526 13524
rect 22646 13472 22652 13524
rect 22704 13512 22710 13524
rect 23290 13512 23296 13524
rect 22704 13484 23296 13512
rect 22704 13472 22710 13484
rect 23290 13472 23296 13484
rect 23348 13512 23354 13524
rect 23569 13515 23627 13521
rect 23569 13512 23581 13515
rect 23348 13484 23581 13512
rect 23348 13472 23354 13484
rect 23569 13481 23581 13484
rect 23615 13481 23627 13515
rect 23569 13475 23627 13481
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 25130 13512 25136 13524
rect 24452 13484 25136 13512
rect 24452 13472 24458 13484
rect 25130 13472 25136 13484
rect 25188 13512 25194 13524
rect 25774 13512 25780 13524
rect 25188 13484 25780 13512
rect 25188 13472 25194 13484
rect 25774 13472 25780 13484
rect 25832 13472 25838 13524
rect 18693 13447 18751 13453
rect 18693 13413 18705 13447
rect 18739 13444 18751 13447
rect 22830 13444 22836 13456
rect 18739 13416 22836 13444
rect 18739 13413 18751 13416
rect 18693 13407 18751 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 25869 13447 25927 13453
rect 25869 13444 25881 13447
rect 23400 13416 25881 13444
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 23014 13376 23020 13388
rect 22051 13348 23020 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19426 13308 19432 13320
rect 19116 13280 19432 13308
rect 19116 13268 19122 13280
rect 19426 13268 19432 13280
rect 19484 13308 19490 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19484 13280 19717 13308
rect 19484 13268 19490 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 20162 13268 20168 13320
rect 20220 13308 20226 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 20220 13280 20637 13308
rect 20220 13268 20226 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 21821 13311 21879 13317
rect 21821 13277 21833 13311
rect 21867 13308 21879 13311
rect 23106 13308 23112 13320
rect 21867 13280 23112 13308
rect 21867 13277 21879 13280
rect 21821 13271 21879 13277
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 23198 13268 23204 13320
rect 23256 13308 23262 13320
rect 23400 13317 23428 13416
rect 25869 13413 25881 13416
rect 25915 13413 25927 13447
rect 25869 13407 25927 13413
rect 24946 13336 24952 13388
rect 25004 13376 25010 13388
rect 25004 13348 25049 13376
rect 25004 13336 25010 13348
rect 23385 13311 23443 13317
rect 23256 13280 23301 13308
rect 23256 13268 23262 13280
rect 23385 13277 23397 13311
rect 23431 13277 23443 13311
rect 25774 13308 25780 13320
rect 25735 13280 25780 13308
rect 23385 13271 23443 13277
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 26602 13308 26608 13320
rect 26563 13280 26608 13308
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 21450 13240 21456 13252
rect 18616 13212 21456 13240
rect 15988 13200 15994 13212
rect 21450 13200 21456 13212
rect 21508 13240 21514 13252
rect 24394 13240 24400 13252
rect 21508 13212 24400 13240
rect 21508 13200 21514 13212
rect 24394 13200 24400 13212
rect 24452 13200 24458 13252
rect 24670 13240 24676 13252
rect 24631 13212 24676 13240
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 24765 13243 24823 13249
rect 24765 13209 24777 13243
rect 24811 13209 24823 13243
rect 24765 13203 24823 13209
rect 25424 13212 26464 13240
rect 10686 13172 10692 13184
rect 9646 13144 10692 13172
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13320 13144 13553 13172
rect 13320 13132 13326 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 14645 13175 14703 13181
rect 14645 13141 14657 13175
rect 14691 13172 14703 13175
rect 16758 13172 16764 13184
rect 14691 13144 16764 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 17129 13175 17187 13181
rect 17129 13141 17141 13175
rect 17175 13172 17187 13175
rect 18046 13172 18052 13184
rect 17175 13144 18052 13172
rect 17175 13141 17187 13144
rect 17129 13135 17187 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 20438 13172 20444 13184
rect 20399 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 20864 13144 21097 13172
rect 20864 13132 20870 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 24780 13172 24808 13203
rect 25424 13172 25452 13212
rect 26436 13181 26464 13212
rect 24780 13144 25452 13172
rect 26421 13175 26479 13181
rect 21085 13135 21143 13141
rect 26421 13141 26433 13175
rect 26467 13141 26479 13175
rect 26421 13135 26479 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 8938 12968 8944 12980
rect 5859 12940 8944 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 11057 12971 11115 12977
rect 9180 12940 11008 12968
rect 9180 12928 9186 12940
rect 6454 12900 6460 12912
rect 2746 12872 6460 12900
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2222 12792 2228 12844
rect 2280 12832 2286 12844
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 2280 12804 2421 12832
rect 2280 12792 2286 12804
rect 2409 12801 2421 12804
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 2746 12764 2774 12872
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 6546 12860 6552 12912
rect 6604 12900 6610 12912
rect 7653 12903 7711 12909
rect 6604 12872 7604 12900
rect 6604 12860 6610 12872
rect 3234 12832 3240 12844
rect 3195 12804 3240 12832
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 5994 12832 6000 12844
rect 5955 12804 6000 12832
rect 4801 12795 4859 12801
rect 1596 12736 2774 12764
rect 1596 12705 1624 12736
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4816 12764 4844 12795
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 7098 12832 7104 12844
rect 6963 12804 7104 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7098 12792 7104 12804
rect 7156 12792 7162 12844
rect 7576 12841 7604 12872
rect 7653 12869 7665 12903
rect 7699 12900 7711 12903
rect 9306 12900 9312 12912
rect 7699 12872 9312 12900
rect 7699 12869 7711 12872
rect 7653 12863 7711 12869
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 9766 12900 9772 12912
rect 9456 12872 9772 12900
rect 9456 12860 9462 12872
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 10980 12900 11008 12940
rect 11057 12937 11069 12971
rect 11103 12968 11115 12971
rect 11882 12968 11888 12980
rect 11103 12940 11888 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12345 12971 12403 12977
rect 12345 12968 12357 12971
rect 12216 12940 12357 12968
rect 12216 12928 12222 12940
rect 12345 12937 12357 12940
rect 12391 12937 12403 12971
rect 12345 12931 12403 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 15470 12968 15476 12980
rect 13127 12940 15476 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17092 12940 18736 12968
rect 17092 12928 17098 12940
rect 18708 12900 18736 12940
rect 18782 12928 18788 12980
rect 18840 12968 18846 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18840 12940 18889 12968
rect 18840 12928 18846 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 20162 12968 20168 12980
rect 20123 12940 20168 12968
rect 18877 12931 18935 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21174 12968 21180 12980
rect 20364 12940 21180 12968
rect 10980 12872 14872 12900
rect 18708 12872 19564 12900
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12801 7619 12835
rect 7561 12795 7619 12801
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 8110 12832 8116 12844
rect 7984 12804 8116 12832
rect 7984 12792 7990 12804
rect 8110 12792 8116 12804
rect 8168 12832 8174 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 8168 12804 8217 12832
rect 8168 12792 8174 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 8343 12804 10609 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11020 12804 12265 12832
rect 11020 12792 11026 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12676 12804 13001 12832
rect 12676 12792 12682 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 12989 12795 13047 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14240 12804 14473 12832
rect 14240 12792 14246 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 4028 12736 4844 12764
rect 4893 12767 4951 12773
rect 4028 12724 4034 12736
rect 4893 12733 4905 12767
rect 4939 12764 4951 12767
rect 7650 12764 7656 12776
rect 4939 12736 7656 12764
rect 4939 12733 4951 12736
rect 4893 12727 4951 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 8812 12736 8861 12764
rect 8812 12724 8818 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8849 12727 8907 12733
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12733 10471 12767
rect 10413 12727 10471 12733
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 14734 12764 14740 12776
rect 14323 12736 14740 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12665 1639 12699
rect 1581 12659 1639 12665
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 4798 12696 4804 12708
rect 3375 12668 4804 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 7009 12699 7067 12705
rect 7009 12665 7021 12699
rect 7055 12696 7067 12699
rect 9048 12696 9076 12727
rect 10428 12696 10456 12727
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14844 12764 14872 12872
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15838 12832 15844 12844
rect 15427 12804 15844 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18564 12804 18797 12832
rect 18564 12792 18570 12804
rect 18785 12801 18797 12804
rect 18831 12832 18843 12835
rect 18874 12832 18880 12844
rect 18831 12804 18880 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19536 12841 19564 12872
rect 20364 12841 20392 12940
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 26145 12971 26203 12977
rect 26145 12968 26157 12971
rect 23400 12940 26157 12968
rect 20438 12860 20444 12912
rect 20496 12900 20502 12912
rect 22186 12900 22192 12912
rect 20496 12872 21036 12900
rect 22147 12872 22192 12900
rect 20496 12860 20502 12872
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12832 19579 12835
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 19567 12804 20361 12832
rect 19567 12801 19579 12804
rect 19521 12795 19579 12801
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20806 12832 20812 12844
rect 20767 12804 20812 12832
rect 20349 12795 20407 12801
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 21008 12841 21036 12872
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 23400 12909 23428 12940
rect 26145 12937 26157 12940
rect 26191 12937 26203 12971
rect 26145 12931 26203 12937
rect 32585 12971 32643 12977
rect 32585 12937 32597 12971
rect 32631 12968 32643 12971
rect 36446 12968 36452 12980
rect 32631 12940 36452 12968
rect 32631 12937 32643 12940
rect 32585 12931 32643 12937
rect 36446 12928 36452 12940
rect 36504 12928 36510 12980
rect 23385 12903 23443 12909
rect 23385 12869 23397 12903
rect 23431 12869 23443 12903
rect 23385 12863 23443 12869
rect 24486 12860 24492 12912
rect 24544 12900 24550 12912
rect 25593 12903 25651 12909
rect 25593 12900 25605 12903
rect 24544 12872 25605 12900
rect 24544 12860 24550 12872
rect 25593 12869 25605 12872
rect 25639 12869 25651 12903
rect 25593 12863 25651 12869
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24670 12832 24676 12844
rect 24443 12804 24676 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 25498 12832 25504 12844
rect 25459 12804 25504 12832
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 14844 12736 15577 12764
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 17681 12767 17739 12773
rect 17681 12733 17693 12767
rect 17727 12764 17739 12767
rect 17770 12764 17776 12776
rect 17727 12736 17776 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 7055 12668 9076 12696
rect 9140 12668 10456 12696
rect 7055 12665 7067 12668
rect 7009 12659 7067 12665
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 8018 12628 8024 12640
rect 3927 12600 8024 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 9140 12628 9168 12668
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 12894 12696 12900 12708
rect 12492 12668 12900 12696
rect 12492 12656 12498 12668
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12696 13691 12699
rect 15378 12696 15384 12708
rect 13679 12668 15384 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 17696 12696 17724 12727
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18230 12764 18236 12776
rect 17911 12736 18236 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21416 12736 22109 12764
rect 21416 12724 21422 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23382 12764 23388 12776
rect 23339 12736 23388 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 23569 12767 23627 12773
rect 23569 12764 23581 12767
rect 23532 12736 23581 12764
rect 23532 12724 23538 12736
rect 23569 12733 23581 12736
rect 23615 12733 23627 12767
rect 23569 12727 23627 12733
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 25222 12764 25228 12776
rect 24627 12736 25228 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 18046 12696 18052 12708
rect 15488 12668 17724 12696
rect 18007 12668 18052 12696
rect 8168 12600 9168 12628
rect 9493 12631 9551 12637
rect 8168 12588 8174 12600
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 10594 12628 10600 12640
rect 9539 12600 10600 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13722 12628 13728 12640
rect 13412 12600 13728 12628
rect 13412 12588 13418 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 14424 12600 14657 12628
rect 14424 12588 14430 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 14645 12591 14703 12597
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 15488 12628 15516 12668
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 22649 12699 22707 12705
rect 22649 12665 22661 12699
rect 22695 12696 22707 12699
rect 24026 12696 24032 12708
rect 22695 12668 24032 12696
rect 22695 12665 22707 12668
rect 22649 12659 22707 12665
rect 24026 12656 24032 12668
rect 24084 12656 24090 12708
rect 26344 12696 26372 12795
rect 29086 12792 29092 12844
rect 29144 12832 29150 12844
rect 32769 12835 32827 12841
rect 32769 12832 32781 12835
rect 29144 12804 32781 12832
rect 29144 12792 29150 12804
rect 32769 12801 32781 12804
rect 32815 12801 32827 12835
rect 38010 12832 38016 12844
rect 37971 12804 38016 12832
rect 32769 12795 32827 12801
rect 38010 12792 38016 12804
rect 38068 12792 38074 12844
rect 24136 12668 26372 12696
rect 14792 12600 15516 12628
rect 16025 12631 16083 12637
rect 14792 12588 14798 12600
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 17034 12628 17040 12640
rect 16071 12600 17040 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 19613 12631 19671 12637
rect 19613 12597 19625 12631
rect 19659 12628 19671 12631
rect 20622 12628 20628 12640
rect 19659 12600 20628 12628
rect 19659 12597 19671 12600
rect 19613 12591 19671 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 21174 12628 21180 12640
rect 21135 12600 21180 12628
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 23198 12588 23204 12640
rect 23256 12628 23262 12640
rect 24136 12628 24164 12668
rect 24854 12628 24860 12640
rect 23256 12600 24164 12628
rect 24815 12600 24860 12628
rect 23256 12588 23262 12600
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5902 12424 5908 12436
rect 5592 12396 5908 12424
rect 5592 12384 5598 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 8478 12424 8484 12436
rect 6595 12396 8484 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 10042 12424 10048 12436
rect 8628 12396 10048 12424
rect 8628 12384 8634 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 12618 12424 12624 12436
rect 11480 12396 12624 12424
rect 11480 12384 11486 12396
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13630 12424 13636 12436
rect 12860 12396 13636 12424
rect 12860 12384 12866 12396
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 15930 12424 15936 12436
rect 15891 12396 15936 12424
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 17276 12396 17601 12424
rect 17276 12384 17282 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 18230 12424 18236 12436
rect 18191 12396 18236 12424
rect 17589 12387 17647 12393
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20404 12396 21005 12424
rect 20404 12384 20410 12396
rect 20993 12393 21005 12396
rect 21039 12393 21051 12427
rect 20993 12387 21051 12393
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 37829 12427 37887 12433
rect 23532 12396 31754 12424
rect 23532 12384 23538 12396
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9769 12359 9827 12365
rect 8996 12328 9444 12356
rect 8996 12316 9002 12328
rect 4614 12288 4620 12300
rect 2240 12260 4620 12288
rect 2240 12229 2268 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 6914 12288 6920 12300
rect 5307 12260 6920 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8294 12288 8300 12300
rect 7883 12260 8300 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 9306 12288 9312 12300
rect 9267 12260 9312 12288
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9416 12288 9444 12328
rect 9769 12325 9781 12359
rect 9815 12356 9827 12359
rect 11517 12359 11575 12365
rect 11517 12356 11529 12359
rect 9815 12328 11529 12356
rect 9815 12325 9827 12328
rect 9769 12319 9827 12325
rect 11517 12325 11529 12328
rect 11563 12356 11575 12359
rect 11563 12328 14412 12356
rect 11563 12325 11575 12328
rect 11517 12319 11575 12325
rect 10962 12288 10968 12300
rect 9416 12260 10968 12288
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11330 12288 11336 12300
rect 11291 12260 11336 12288
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11974 12288 11980 12300
rect 11664 12260 11980 12288
rect 11664 12248 11670 12260
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 13906 12288 13912 12300
rect 13004 12260 13912 12288
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 1780 12152 1808 12183
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2832 12192 2881 12220
rect 2832 12180 2838 12192
rect 2869 12189 2881 12192
rect 2915 12220 2927 12223
rect 3234 12220 3240 12232
rect 2915 12192 3240 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 3970 12220 3976 12232
rect 3844 12192 3976 12220
rect 3844 12180 3850 12192
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5215 12192 5825 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5813 12189 5825 12192
rect 5859 12220 5871 12223
rect 5902 12220 5908 12232
rect 5859 12192 5908 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 6454 12220 6460 12232
rect 6415 12192 6460 12220
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 7248 12192 7297 12220
rect 7248 12180 7254 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 8570 12220 8576 12232
rect 7800 12192 7845 12220
rect 8531 12192 8576 12220
rect 7800 12180 7806 12192
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8720 12192 9137 12220
rect 8720 12180 8726 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10689 12223 10747 12229
rect 10520 12220 10617 12222
rect 10689 12220 10701 12223
rect 10008 12194 10701 12220
rect 10008 12192 10548 12194
rect 10589 12192 10701 12194
rect 10008 12180 10014 12192
rect 10689 12189 10701 12192
rect 10735 12220 10747 12223
rect 10870 12220 10876 12232
rect 10735 12192 10876 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11112 12192 11161 12220
rect 11112 12180 11118 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 3050 12152 3056 12164
rect 1780 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3252 12152 3280 12180
rect 13004 12164 13032 12260
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14384 12297 14412 12328
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 23845 12359 23903 12365
rect 15436 12328 16896 12356
rect 15436 12316 15442 12328
rect 14369 12291 14427 12297
rect 14369 12257 14381 12291
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 15010 12288 15016 12300
rect 14608 12260 15016 12288
rect 14608 12248 14614 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16172 12260 16497 12288
rect 16172 12248 16178 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 16868 12288 16896 12328
rect 23845 12325 23857 12359
rect 23891 12356 23903 12359
rect 24486 12356 24492 12368
rect 23891 12328 24492 12356
rect 23891 12325 23903 12328
rect 23845 12319 23903 12325
rect 24486 12316 24492 12328
rect 24544 12356 24550 12368
rect 24949 12359 25007 12365
rect 24949 12356 24961 12359
rect 24544 12328 24961 12356
rect 24544 12316 24550 12328
rect 24949 12325 24961 12328
rect 24995 12325 25007 12359
rect 24949 12319 25007 12325
rect 20073 12291 20131 12297
rect 16724 12260 16769 12288
rect 16868 12260 20024 12288
rect 16724 12248 16730 12260
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13633 12223 13691 12229
rect 13633 12220 13645 12223
rect 13412 12192 13645 12220
rect 13412 12180 13418 12192
rect 13633 12189 13645 12192
rect 13679 12189 13691 12223
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 13633 12183 13691 12189
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17184 12192 17785 12220
rect 17184 12180 17190 12192
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 19996 12229 20024 12260
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20119 12260 20821 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 20809 12257 20821 12260
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12288 23259 12291
rect 23290 12288 23296 12300
rect 23247 12260 23296 12288
rect 23247 12257 23259 12260
rect 23201 12251 23259 12257
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 23624 12260 24593 12288
rect 23624 12248 23630 12260
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18196 12192 18429 12220
rect 18196 12180 18202 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12220 20039 12223
rect 20254 12220 20260 12232
rect 20027 12192 20260 12220
rect 20027 12189 20039 12192
rect 19981 12183 20039 12189
rect 20254 12180 20260 12192
rect 20312 12180 20318 12232
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 4065 12155 4123 12161
rect 3252 12124 4016 12152
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 2317 12087 2375 12093
rect 2317 12053 2329 12087
rect 2363 12084 2375 12087
rect 2406 12084 2412 12096
rect 2363 12056 2412 12084
rect 2363 12053 2375 12056
rect 2317 12047 2375 12053
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 2961 12087 3019 12093
rect 2961 12053 2973 12087
rect 3007 12084 3019 12087
rect 3602 12084 3608 12096
rect 3007 12056 3608 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3988 12084 4016 12124
rect 4065 12121 4077 12155
rect 4111 12152 4123 12155
rect 5534 12152 5540 12164
rect 4111 12124 5540 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 10520 12124 11928 12152
rect 4614 12084 4620 12096
rect 3988 12056 4620 12084
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 7006 12084 7012 12096
rect 5951 12056 7012 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8386 12084 8392 12096
rect 7156 12056 7201 12084
rect 8347 12056 8392 12084
rect 7156 12044 7162 12056
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 10042 12084 10048 12096
rect 8536 12056 10048 12084
rect 8536 12044 8542 12056
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10520 12093 10548 12124
rect 10505 12087 10563 12093
rect 10505 12053 10517 12087
rect 10551 12053 10563 12087
rect 11900 12084 11928 12124
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12345 12155 12403 12161
rect 12345 12152 12357 12155
rect 12032 12124 12357 12152
rect 12032 12112 12038 12124
rect 12345 12121 12357 12124
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12434 12112 12440 12164
rect 12492 12152 12498 12164
rect 12986 12152 12992 12164
rect 12492 12124 12537 12152
rect 12947 12124 12992 12152
rect 12492 12112 12498 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 14461 12155 14519 12161
rect 14461 12152 14473 12155
rect 13228 12124 14473 12152
rect 13228 12112 13234 12124
rect 14461 12121 14473 12124
rect 14507 12121 14519 12155
rect 14461 12115 14519 12121
rect 15013 12155 15071 12161
rect 15013 12121 15025 12155
rect 15059 12152 15071 12155
rect 17218 12152 17224 12164
rect 15059 12124 17224 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 17310 12112 17316 12164
rect 17368 12152 17374 12164
rect 20640 12152 20668 12183
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 22097 12223 22155 12229
rect 22097 12220 22109 12223
rect 21232 12192 22109 12220
rect 21232 12180 21238 12192
rect 22097 12189 22109 12192
rect 22143 12189 22155 12223
rect 22097 12183 22155 12189
rect 22281 12223 22339 12229
rect 22281 12189 22293 12223
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 24210 12220 24216 12232
rect 23431 12192 24216 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 22296 12152 22324 12183
rect 24210 12180 24216 12192
rect 24268 12180 24274 12232
rect 24762 12220 24768 12232
rect 24723 12192 24768 12220
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 31726 12220 31754 12396
rect 37829 12393 37841 12427
rect 37875 12424 37887 12427
rect 38010 12424 38016 12436
rect 37875 12396 38016 12424
rect 37875 12393 37887 12396
rect 37829 12387 37887 12393
rect 38010 12384 38016 12396
rect 38068 12384 38074 12436
rect 36909 12223 36967 12229
rect 36909 12220 36921 12223
rect 31726 12192 36921 12220
rect 36909 12189 36921 12192
rect 36955 12189 36967 12223
rect 36909 12183 36967 12189
rect 37001 12223 37059 12229
rect 37001 12189 37013 12223
rect 37047 12220 37059 12223
rect 38013 12223 38071 12229
rect 38013 12220 38025 12223
rect 37047 12192 38025 12220
rect 37047 12189 37059 12192
rect 37001 12183 37059 12189
rect 38013 12189 38025 12192
rect 38059 12189 38071 12223
rect 38013 12183 38071 12189
rect 17368 12124 17816 12152
rect 20640 12124 22094 12152
rect 22296 12124 22876 12152
rect 17368 12112 17374 12124
rect 12250 12084 12256 12096
rect 11900 12056 12256 12084
rect 10505 12047 10563 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 12952 12056 13461 12084
rect 12952 12044 12958 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 15562 12084 15568 12096
rect 14332 12056 15568 12084
rect 14332 12044 14338 12056
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 17092 12056 17141 12084
rect 17092 12044 17098 12056
rect 17129 12053 17141 12056
rect 17175 12084 17187 12087
rect 17678 12084 17684 12096
rect 17175 12056 17684 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17788 12084 17816 12124
rect 21910 12084 21916 12096
rect 17788 12056 21916 12084
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22066 12084 22094 12124
rect 22462 12084 22468 12096
rect 22066 12056 22468 12084
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 22738 12084 22744 12096
rect 22699 12056 22744 12084
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 22848 12084 22876 12124
rect 22922 12112 22928 12164
rect 22980 12152 22986 12164
rect 25685 12155 25743 12161
rect 25685 12152 25697 12155
rect 22980 12124 25697 12152
rect 22980 12112 22986 12124
rect 25685 12121 25697 12124
rect 25731 12121 25743 12155
rect 25685 12115 25743 12121
rect 23750 12084 23756 12096
rect 22848 12056 23756 12084
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 7101 11883 7159 11889
rect 1636 11852 5856 11880
rect 1636 11840 1642 11852
rect 5350 11812 5356 11824
rect 4370 11784 5356 11812
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1544 11716 1777 11744
rect 1544 11704 1550 11716
rect 1765 11713 1777 11716
rect 1811 11713 1823 11747
rect 2406 11744 2412 11756
rect 2367 11716 2412 11744
rect 1765 11707 1823 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 5828 11753 5856 11852
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 8294 11880 8300 11892
rect 7147 11852 8300 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 8536 11852 8892 11880
rect 8536 11840 8542 11852
rect 8864 11812 8892 11852
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9398 11880 9404 11892
rect 8996 11852 9404 11880
rect 8996 11840 9002 11852
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9677 11883 9735 11889
rect 9677 11849 9689 11883
rect 9723 11880 9735 11883
rect 11974 11880 11980 11892
rect 9723 11852 11980 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12434 11880 12440 11892
rect 12124 11852 12440 11880
rect 12124 11840 12130 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 18138 11880 18144 11892
rect 18099 11852 18144 11880
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18230 11840 18236 11892
rect 18288 11880 18294 11892
rect 20254 11880 20260 11892
rect 18288 11852 20260 11880
rect 18288 11840 18294 11852
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 21174 11880 21180 11892
rect 21131 11852 21180 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 22002 11880 22008 11892
rect 21963 11852 22008 11880
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 24946 11880 24952 11892
rect 22520 11852 24952 11880
rect 22520 11840 22526 11852
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25222 11880 25228 11892
rect 25183 11852 25228 11880
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 25869 11883 25927 11889
rect 25869 11849 25881 11883
rect 25915 11849 25927 11883
rect 25869 11843 25927 11849
rect 12621 11815 12679 11821
rect 12621 11812 12633 11815
rect 8864 11784 12633 11812
rect 12621 11781 12633 11784
rect 12667 11781 12679 11815
rect 14182 11812 14188 11824
rect 12621 11775 12679 11781
rect 14016 11784 14188 11812
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4672 11716 5181 11744
rect 4672 11704 4678 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7331 11716 7420 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 5718 11676 5724 11688
rect 3191 11648 5724 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 5718 11636 5724 11648
rect 5776 11676 5782 11688
rect 7190 11676 7196 11688
rect 5776 11648 7196 11676
rect 5776 11636 5782 11648
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7392 11676 7420 11716
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 7745 11747 7803 11753
rect 7745 11744 7757 11747
rect 7616 11716 7757 11744
rect 7616 11704 7622 11716
rect 7745 11713 7757 11716
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 8573 11747 8631 11753
rect 9217 11748 9275 11753
rect 8573 11713 8585 11747
rect 8619 11713 8631 11747
rect 9140 11747 9275 11748
rect 9140 11744 9229 11747
rect 9048 11742 9229 11744
rect 8573 11707 8631 11713
rect 8864 11720 9229 11742
rect 8864 11716 9168 11720
rect 8864 11714 9076 11716
rect 7466 11676 7472 11688
rect 7392 11648 7472 11676
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 8294 11676 8300 11688
rect 7760 11648 8300 11676
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 1627 11580 2774 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 1912 11512 2237 11540
rect 1912 11500 1918 11512
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2746 11540 2774 11580
rect 4154 11568 4160 11620
rect 4212 11608 4218 11620
rect 5261 11611 5319 11617
rect 5261 11608 5273 11611
rect 4212 11580 5273 11608
rect 4212 11568 4218 11580
rect 5261 11577 5273 11580
rect 5307 11577 5319 11611
rect 5261 11571 5319 11577
rect 5905 11611 5963 11617
rect 5905 11577 5917 11611
rect 5951 11608 5963 11611
rect 7760 11608 7788 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8588 11676 8616 11707
rect 8662 11676 8668 11688
rect 8588 11648 8668 11676
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 5951 11580 7788 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8202 11608 8208 11620
rect 7984 11580 8208 11608
rect 7984 11568 7990 11580
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8389 11611 8447 11617
rect 8389 11577 8401 11611
rect 8435 11608 8447 11611
rect 8864 11608 8892 11714
rect 9217 11713 9229 11720
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 9364 11716 10517 11744
rect 9364 11704 9370 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10962 11744 10968 11756
rect 10923 11716 10968 11744
rect 10505 11707 10563 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11514 11744 11520 11756
rect 11103 11716 11520 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 14016 11753 14044 11784
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 14274 11772 14280 11824
rect 14332 11812 14338 11824
rect 19886 11812 19892 11824
rect 14332 11784 14377 11812
rect 15502 11784 17816 11812
rect 14332 11772 14338 11784
rect 14001 11747 14059 11753
rect 11624 11716 11928 11744
rect 9398 11676 9404 11688
rect 9048 11648 9404 11676
rect 9048 11617 9076 11648
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 9766 11676 9772 11688
rect 9640 11648 9772 11676
rect 9640 11636 9646 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 11624 11676 11652 11716
rect 11790 11676 11796 11688
rect 10152 11648 11652 11676
rect 11751 11648 11796 11676
rect 8435 11580 8892 11608
rect 9033 11611 9091 11617
rect 8435 11577 8447 11580
rect 8389 11571 8447 11577
rect 9033 11577 9045 11611
rect 9079 11577 9091 11611
rect 10152 11608 10180 11648
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11900 11676 11928 11716
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 15838 11704 15844 11756
rect 15896 11744 15902 11756
rect 17310 11744 17316 11756
rect 15896 11716 17316 11744
rect 15896 11704 15902 11716
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 17788 11744 17816 11784
rect 18340 11784 19892 11812
rect 18340 11756 18368 11784
rect 19886 11772 19892 11784
rect 19944 11772 19950 11824
rect 20162 11812 20168 11824
rect 19996 11784 20168 11812
rect 18230 11744 18236 11756
rect 17788 11716 18236 11744
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 18380 11716 18425 11744
rect 18380 11704 18386 11716
rect 18598 11704 18604 11756
rect 18656 11744 18662 11756
rect 19996 11753 20024 11784
rect 20162 11772 20168 11784
rect 20220 11812 20226 11824
rect 21818 11812 21824 11824
rect 20220 11784 21824 11812
rect 20220 11772 20226 11784
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 23014 11812 23020 11824
rect 22975 11784 23020 11812
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 24213 11815 24271 11821
rect 24213 11781 24225 11815
rect 24259 11812 24271 11815
rect 25314 11812 25320 11824
rect 24259 11784 25320 11812
rect 24259 11781 24271 11784
rect 24213 11775 24271 11781
rect 25314 11772 25320 11784
rect 25372 11772 25378 11824
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 18656 11716 18797 11744
rect 18656 11704 18662 11716
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11713 20039 11747
rect 20622 11744 20628 11756
rect 20583 11716 20628 11744
rect 19981 11707 20039 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 25409 11747 25467 11753
rect 25409 11713 25421 11747
rect 25455 11744 25467 11747
rect 25884 11744 25912 11843
rect 26050 11744 26056 11756
rect 25455 11716 25912 11744
rect 26011 11716 26056 11744
rect 25455 11713 25467 11716
rect 25409 11707 25467 11713
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 11900 11648 12541 11676
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 9033 11571 9091 11577
rect 9232 11580 10180 11608
rect 10321 11611 10379 11617
rect 3878 11540 3884 11552
rect 2746 11512 3884 11540
rect 2225 11503 2283 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4614 11540 4620 11552
rect 4575 11512 4620 11540
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 7558 11540 7564 11552
rect 6236 11512 7564 11540
rect 6236 11500 6242 11512
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 9232 11540 9260 11580
rect 10321 11577 10333 11611
rect 10367 11608 10379 11611
rect 10410 11608 10416 11620
rect 10367 11580 10416 11608
rect 10367 11577 10379 11580
rect 10321 11571 10379 11577
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 12544 11608 12572 11639
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12768 11648 12817 11676
rect 12768 11636 12774 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 20438 11676 20444 11688
rect 12805 11639 12863 11645
rect 12912 11648 20444 11676
rect 12912 11608 12940 11648
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 12544 11580 12940 11608
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 22204 11608 22232 11707
rect 26050 11704 26056 11716
rect 26108 11704 26114 11756
rect 22922 11676 22928 11688
rect 22883 11648 22928 11676
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23569 11679 23627 11685
rect 23569 11645 23581 11679
rect 23615 11676 23627 11679
rect 23658 11676 23664 11688
rect 23615 11648 23664 11676
rect 23615 11645 23627 11648
rect 23569 11639 23627 11645
rect 23658 11636 23664 11648
rect 23716 11676 23722 11688
rect 23934 11676 23940 11688
rect 23716 11648 23940 11676
rect 23716 11636 23722 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11676 24179 11679
rect 24854 11676 24860 11688
rect 24167 11648 24860 11676
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 24854 11636 24860 11648
rect 24912 11676 24918 11688
rect 25038 11676 25044 11688
rect 24912 11648 25044 11676
rect 24912 11636 24918 11648
rect 25038 11636 25044 11648
rect 25096 11636 25102 11688
rect 23842 11608 23848 11620
rect 16172 11580 23848 11608
rect 16172 11568 16178 11580
rect 23842 11568 23848 11580
rect 23900 11568 23906 11620
rect 24302 11568 24308 11620
rect 24360 11608 24366 11620
rect 24670 11608 24676 11620
rect 24360 11580 24676 11608
rect 24360 11568 24366 11580
rect 24670 11568 24676 11580
rect 24728 11568 24734 11620
rect 7883 11512 9260 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10502 11540 10508 11552
rect 9824 11512 10508 11540
rect 9824 11500 9830 11512
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 15470 11540 15476 11552
rect 11848 11512 15476 11540
rect 11848 11500 11854 11512
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15749 11543 15807 11549
rect 15749 11509 15761 11543
rect 15795 11540 15807 11543
rect 15930 11540 15936 11552
rect 15795 11512 15936 11540
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 15930 11500 15936 11512
rect 15988 11540 15994 11552
rect 16390 11540 16396 11552
rect 15988 11512 16396 11540
rect 15988 11500 15994 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18840 11512 18889 11540
rect 18840 11500 18846 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 20346 11540 20352 11552
rect 19843 11512 20352 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 25866 11540 25872 11552
rect 20588 11512 25872 11540
rect 20588 11500 20594 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 4062 11336 4068 11348
rect 1627 11308 4068 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4236 11339 4294 11345
rect 4236 11305 4248 11339
rect 4282 11336 4294 11339
rect 8202 11336 8208 11348
rect 4282 11308 8208 11336
rect 4282 11305 4294 11308
rect 4236 11299 4294 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 12066 11336 12072 11348
rect 9456 11308 12072 11336
rect 9456 11296 9462 11308
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15856 11308 16037 11336
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11237 2651 11271
rect 2593 11231 2651 11237
rect 2608 11200 2636 11231
rect 3510 11228 3516 11280
rect 3568 11268 3574 11280
rect 3970 11268 3976 11280
rect 3568 11240 3976 11268
rect 3568 11228 3574 11240
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 5718 11268 5724 11280
rect 5679 11240 5724 11268
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 10594 11268 10600 11280
rect 8352 11240 10456 11268
rect 10555 11240 10600 11268
rect 8352 11228 8358 11240
rect 2608 11172 3280 11200
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 3252 11141 3280 11172
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 6273 11203 6331 11209
rect 3936 11172 6224 11200
rect 3936 11160 3942 11172
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11101 3295 11135
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3237 11095 3295 11101
rect 2792 11064 2820 11095
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 6086 11132 6092 11144
rect 5382 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6196 11141 6224 11172
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 9766 11200 9772 11212
rect 6319 11172 9772 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10318 11200 10324 11212
rect 9999 11172 10324 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10428 11200 10456 11240
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 11054 11228 11060 11280
rect 11112 11228 11118 11280
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 13541 11271 13599 11277
rect 12492 11240 12940 11268
rect 12492 11228 12498 11240
rect 11072 11200 11100 11228
rect 10428 11172 11100 11200
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11422 11200 11428 11212
rect 11379 11172 11428 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 11940 11172 12817 11200
rect 11940 11160 11946 11172
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 6788 11104 6837 11132
rect 6788 11092 6794 11104
rect 6825 11101 6837 11104
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 9490 11132 9496 11144
rect 8444 11104 9496 11132
rect 8444 11092 8450 11104
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9732 11104 10149 11132
rect 9732 11092 9738 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 10137 11095 10195 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 12912 11132 12940 11240
rect 13541 11237 13553 11271
rect 13587 11237 13599 11271
rect 13541 11231 13599 11237
rect 13556 11200 13584 11231
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 15856 11268 15884 11308
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 16850 11336 16856 11348
rect 16025 11299 16083 11305
rect 16132 11308 16856 11336
rect 15804 11240 15884 11268
rect 15804 11228 15810 11240
rect 16132 11200 16160 11308
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 20530 11336 20536 11348
rect 19484 11308 20536 11336
rect 19484 11296 19490 11308
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 21821 11339 21879 11345
rect 21821 11305 21833 11339
rect 21867 11336 21879 11339
rect 22186 11336 22192 11348
rect 21867 11308 22192 11336
rect 21867 11305 21879 11308
rect 21821 11299 21879 11305
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 24581 11339 24639 11345
rect 22480 11308 23704 11336
rect 16390 11228 16396 11280
rect 16448 11268 16454 11280
rect 18966 11268 18972 11280
rect 16448 11240 18972 11268
rect 16448 11228 16454 11240
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 19705 11271 19763 11277
rect 19705 11237 19717 11271
rect 19751 11268 19763 11271
rect 20990 11268 20996 11280
rect 19751 11240 20996 11268
rect 19751 11237 19763 11240
rect 19705 11231 19763 11237
rect 20990 11228 20996 11240
rect 21048 11228 21054 11280
rect 22480 11268 22508 11308
rect 21744 11240 22508 11268
rect 13556 11172 16160 11200
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 16264 11172 16589 11200
rect 16264 11160 16270 11172
rect 16577 11169 16589 11172
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 16758 11160 16764 11212
rect 16816 11200 16822 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16816 11172 16865 11200
rect 16816 11160 16822 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 20349 11203 20407 11209
rect 20349 11169 20361 11203
rect 20395 11200 20407 11203
rect 20438 11200 20444 11212
rect 20395 11172 20444 11200
rect 20395 11169 20407 11172
rect 20349 11163 20407 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 12912 11104 13737 11132
rect 13725 11101 13737 11104
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14240 11104 14289 11132
rect 14240 11092 14246 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 16390 11132 16396 11144
rect 15686 11104 16396 11132
rect 14277 11095 14335 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 19889 11135 19947 11141
rect 18288 11104 19840 11132
rect 18288 11092 18294 11104
rect 3329 11067 3387 11073
rect 2792 11036 3280 11064
rect 3252 10996 3280 11036
rect 3329 11033 3341 11067
rect 3375 11064 3387 11067
rect 3375 11036 4660 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 4522 10996 4528 11008
rect 3252 10968 4528 10996
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 4632 10996 4660 11036
rect 5552 11036 7052 11064
rect 5552 10996 5580 11036
rect 4632 10968 5580 10996
rect 7024 10996 7052 11036
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 7156 11036 7201 11064
rect 7156 11024 7162 11036
rect 7558 11024 7564 11076
rect 7616 11024 7622 11076
rect 8404 11036 11744 11064
rect 8404 10996 8432 11036
rect 7024 10968 8432 10996
rect 8573 10999 8631 11005
rect 8573 10965 8585 10999
rect 8619 10996 8631 10999
rect 8662 10996 8668 11008
rect 8619 10968 8668 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 8662 10956 8668 10968
rect 8720 10996 8726 11008
rect 10410 10996 10416 11008
rect 8720 10968 10416 10996
rect 8720 10956 8726 10968
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 11716 10996 11744 11036
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 14553 11067 14611 11073
rect 14553 11033 14565 11067
rect 14599 11064 14611 11067
rect 14599 11036 14964 11064
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 13814 10996 13820 11008
rect 11716 10968 13820 10996
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 14826 10996 14832 11008
rect 13964 10968 14832 10996
rect 13964 10956 13970 10968
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 14936 10996 14964 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16669 11067 16727 11073
rect 16669 11064 16681 11067
rect 15896 11036 16681 11064
rect 15896 11024 15902 11036
rect 16669 11033 16681 11036
rect 16715 11033 16727 11067
rect 16669 11027 16727 11033
rect 17494 11024 17500 11076
rect 17552 11064 17558 11076
rect 17773 11067 17831 11073
rect 17773 11064 17785 11067
rect 17552 11036 17785 11064
rect 17552 11024 17558 11036
rect 17773 11033 17785 11036
rect 17819 11033 17831 11067
rect 17773 11027 17831 11033
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 18325 11067 18383 11073
rect 18325 11064 18337 11067
rect 17920 11036 18337 11064
rect 17920 11024 17926 11036
rect 18325 11033 18337 11036
rect 18371 11033 18383 11067
rect 19812 11064 19840 11104
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 19978 11132 19984 11144
rect 19935 11104 19984 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20530 11132 20536 11144
rect 20491 11104 20536 11132
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 21744 11141 21772 11240
rect 22554 11228 22560 11280
rect 22612 11228 22618 11280
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 22572 11200 22600 11228
rect 22419 11172 22600 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 20640 11104 21741 11132
rect 20640 11064 20668 11104
rect 21729 11101 21741 11104
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 23676 11141 23704 11308
rect 24581 11305 24593 11339
rect 24627 11336 24639 11339
rect 24762 11336 24768 11348
rect 24627 11308 24768 11336
rect 24627 11305 24639 11308
rect 24581 11299 24639 11305
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 25314 11336 25320 11348
rect 25275 11308 25320 11336
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 25961 11339 26019 11345
rect 25961 11305 25973 11339
rect 26007 11336 26019 11339
rect 29086 11336 29092 11348
rect 26007 11308 29092 11336
rect 26007 11305 26019 11308
rect 25961 11299 26019 11305
rect 29086 11296 29092 11308
rect 29144 11296 29150 11348
rect 23842 11228 23848 11280
rect 23900 11268 23906 11280
rect 25498 11268 25504 11280
rect 23900 11240 25504 11268
rect 23900 11228 23906 11240
rect 25498 11228 25504 11240
rect 25556 11228 25562 11280
rect 38194 11268 38200 11280
rect 38155 11240 38200 11268
rect 38194 11228 38200 11240
rect 38252 11228 38258 11280
rect 25774 11200 25780 11212
rect 25240 11172 25780 11200
rect 25240 11144 25268 11172
rect 25774 11160 25780 11172
rect 25832 11160 25838 11212
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22520 11104 22569 11132
rect 22520 11092 22526 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 23661 11135 23719 11141
rect 23661 11101 23673 11135
rect 23707 11101 23719 11135
rect 24762 11132 24768 11144
rect 24723 11104 24768 11132
rect 23661 11095 23719 11101
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 25222 11132 25228 11144
rect 25183 11104 25228 11132
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 25866 11132 25872 11144
rect 25827 11104 25872 11132
rect 25866 11092 25872 11104
rect 25924 11092 25930 11144
rect 26973 11135 27031 11141
rect 26973 11101 26985 11135
rect 27019 11101 27031 11135
rect 26973 11095 27031 11101
rect 19812 11036 20668 11064
rect 20993 11067 21051 11073
rect 18325 11027 18383 11033
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 22094 11064 22100 11076
rect 21039 11036 22100 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 22738 11024 22744 11076
rect 22796 11064 22802 11076
rect 23017 11067 23075 11073
rect 23017 11064 23029 11067
rect 22796 11036 23029 11064
rect 22796 11024 22802 11036
rect 23017 11033 23029 11036
rect 23063 11064 23075 11067
rect 26988 11064 27016 11095
rect 36078 11092 36084 11144
rect 36136 11132 36142 11144
rect 38013 11135 38071 11141
rect 38013 11132 38025 11135
rect 36136 11104 38025 11132
rect 36136 11092 36142 11104
rect 38013 11101 38025 11104
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 23063 11036 27016 11064
rect 27065 11067 27123 11073
rect 23063 11033 23075 11036
rect 23017 11027 23075 11033
rect 27065 11033 27077 11067
rect 27111 11064 27123 11067
rect 28902 11064 28908 11076
rect 27111 11036 28908 11064
rect 27111 11033 27123 11036
rect 27065 11027 27123 11033
rect 28902 11024 28908 11036
rect 28960 11024 28966 11076
rect 16114 10996 16120 11008
rect 14936 10968 16120 10996
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 17954 10996 17960 11008
rect 16264 10968 17960 10996
rect 16264 10956 16270 10968
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 18414 10956 18420 11008
rect 18472 10996 18478 11008
rect 23290 10996 23296 11008
rect 18472 10968 23296 10996
rect 18472 10956 18478 10968
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 23474 10996 23480 11008
rect 23435 10968 23480 10996
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 3694 10792 3700 10804
rect 1627 10764 3700 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 7009 10795 7067 10801
rect 4212 10764 5948 10792
rect 4212 10752 4218 10764
rect 5718 10724 5724 10736
rect 4554 10696 5724 10724
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2498 10616 2504 10668
rect 2556 10656 2562 10668
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 2556 10628 2605 10656
rect 2556 10616 2562 10628
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 2593 10619 2651 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 5920 10656 5948 10764
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 11057 10795 11115 10801
rect 7055 10764 9812 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 8386 10724 8392 10736
rect 7576 10696 8392 10724
rect 7576 10665 7604 10696
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 9784 10724 9812 10764
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 15838 10792 15844 10804
rect 11103 10764 15844 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16114 10792 16120 10804
rect 15979 10764 16120 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 20165 10795 20223 10801
rect 16408 10764 20116 10792
rect 12342 10724 12348 10736
rect 8536 10696 8970 10724
rect 9784 10696 12348 10724
rect 8536 10684 8542 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12802 10684 12808 10736
rect 12860 10684 12866 10736
rect 16408 10724 16436 10764
rect 15686 10696 16436 10724
rect 16850 10684 16856 10736
rect 16908 10724 16914 10736
rect 16945 10727 17003 10733
rect 16945 10724 16957 10727
rect 16908 10696 16957 10724
rect 16908 10684 16914 10696
rect 16945 10693 16957 10696
rect 16991 10693 17003 10727
rect 16945 10687 17003 10693
rect 17310 10684 17316 10736
rect 17368 10724 17374 10736
rect 19886 10724 19892 10736
rect 17368 10696 19892 10724
rect 17368 10684 17374 10696
rect 19886 10684 19892 10696
rect 19944 10684 19950 10736
rect 20088 10724 20116 10764
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20530 10792 20536 10804
rect 20211 10764 20536 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 23750 10792 23756 10804
rect 23711 10764 23756 10792
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 25038 10792 25044 10804
rect 24999 10764 25044 10792
rect 25038 10752 25044 10764
rect 25096 10752 25102 10804
rect 20622 10724 20628 10736
rect 20088 10696 20628 10724
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 22649 10727 22707 10733
rect 22649 10724 22661 10727
rect 22152 10696 22661 10724
rect 22152 10684 22158 10696
rect 22649 10693 22661 10696
rect 22695 10693 22707 10727
rect 22649 10687 22707 10693
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10724 22799 10727
rect 25593 10727 25651 10733
rect 25593 10724 25605 10727
rect 22787 10696 25605 10724
rect 22787 10693 22799 10696
rect 22741 10687 22799 10693
rect 25593 10693 25605 10696
rect 25639 10693 25651 10727
rect 25593 10687 25651 10693
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 5920 10628 6929 10656
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 10192 10628 10241 10656
rect 10192 10616 10198 10628
rect 10229 10625 10241 10628
rect 10275 10656 10287 10659
rect 10686 10656 10692 10668
rect 10275 10628 10692 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10836 10628 10977 10656
rect 10836 10616 10842 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 10965 10619 11023 10625
rect 11900 10628 11989 10656
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 3016 10560 3065 10588
rect 3016 10548 3022 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3418 10588 3424 10600
rect 3375 10560 3424 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3418 10548 3424 10560
rect 3476 10588 3482 10600
rect 7742 10588 7748 10600
rect 3476 10560 7748 10588
rect 3476 10548 3482 10560
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 8202 10588 8208 10600
rect 8163 10560 8208 10588
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 10594 10588 10600 10600
rect 8527 10560 10600 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11900 10588 11928 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 20346 10656 20352 10668
rect 11977 10619 12035 10625
rect 17512 10628 19656 10656
rect 20307 10628 20352 10656
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11112 10560 11928 10588
rect 11992 10560 12265 10588
rect 11112 10548 11118 10560
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 8110 10520 8116 10532
rect 5951 10492 8116 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 11882 10520 11888 10532
rect 9548 10492 11888 10520
rect 9548 10480 9554 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 1728 10424 2421 10452
rect 1728 10412 1734 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2409 10415 2467 10421
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 7466 10452 7472 10464
rect 4847 10424 7472 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7653 10455 7711 10461
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 9122 10452 9128 10464
rect 7699 10424 9128 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10686 10452 10692 10464
rect 10100 10424 10692 10452
rect 10100 10412 10106 10424
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11992 10452 12020 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 12253 10551 12311 10557
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 15528 10560 16865 10588
rect 15528 10548 15534 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 17126 10588 17132 10600
rect 17087 10560 17132 10588
rect 16853 10551 16911 10557
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17512 10588 17540 10628
rect 18598 10588 18604 10600
rect 17276 10560 17540 10588
rect 18559 10560 18604 10588
rect 17276 10548 17282 10560
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 18785 10591 18843 10597
rect 18785 10557 18797 10591
rect 18831 10557 18843 10591
rect 19518 10588 19524 10600
rect 19479 10560 19524 10588
rect 18785 10551 18843 10557
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 13872 10492 14320 10520
rect 13872 10480 13878 10492
rect 10928 10424 12020 10452
rect 13725 10455 13783 10461
rect 10928 10412 10934 10424
rect 13725 10421 13737 10455
rect 13771 10452 13783 10455
rect 13906 10452 13912 10464
rect 13771 10424 13912 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 14292 10452 14320 10492
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16206 10520 16212 10532
rect 15620 10492 16212 10520
rect 15620 10480 15626 10492
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 18800 10520 18828 10551
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 19628 10588 19656 10628
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10656 23351 10659
rect 23382 10656 23388 10668
rect 23339 10628 23388 10656
rect 23339 10625 23351 10628
rect 23293 10619 23351 10625
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 23934 10656 23940 10668
rect 23895 10628 23940 10656
rect 23934 10616 23940 10628
rect 23992 10616 23998 10668
rect 24026 10616 24032 10668
rect 24084 10656 24090 10668
rect 25501 10659 25559 10665
rect 25501 10656 25513 10659
rect 24084 10628 25513 10656
rect 24084 10616 24090 10628
rect 25501 10625 25513 10628
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 24118 10588 24124 10600
rect 19628 10560 24124 10588
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24397 10591 24455 10597
rect 24397 10557 24409 10591
rect 24443 10557 24455 10591
rect 24397 10551 24455 10557
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 25314 10588 25320 10600
rect 24627 10560 25320 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 17788 10492 18828 10520
rect 17788 10461 17816 10492
rect 18874 10480 18880 10532
rect 18932 10520 18938 10532
rect 23382 10520 23388 10532
rect 18932 10492 23388 10520
rect 18932 10480 18938 10492
rect 23382 10480 23388 10492
rect 23440 10480 23446 10532
rect 24412 10520 24440 10551
rect 25314 10548 25320 10560
rect 25372 10548 25378 10600
rect 33686 10520 33692 10532
rect 24412 10492 33692 10520
rect 33686 10480 33692 10492
rect 33744 10480 33750 10532
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 14292 10424 17785 10452
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 17773 10415 17831 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 20162 10452 20168 10464
rect 18564 10424 20168 10452
rect 18564 10412 18570 10424
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20809 10455 20867 10461
rect 20809 10421 20821 10455
rect 20855 10452 20867 10455
rect 20990 10452 20996 10464
rect 20855 10424 20996 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1936 10251 1994 10257
rect 1936 10217 1948 10251
rect 1982 10248 1994 10251
rect 3418 10248 3424 10260
rect 1982 10220 3280 10248
rect 3379 10220 3424 10248
rect 1982 10217 1994 10220
rect 1936 10211 1994 10217
rect 3252 10180 3280 10220
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 5258 10248 5264 10260
rect 4764 10220 5264 10248
rect 4764 10208 4770 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 8110 10248 8116 10260
rect 6972 10220 8116 10248
rect 6972 10208 6978 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9388 10251 9446 10257
rect 9388 10217 9400 10251
rect 9434 10248 9446 10251
rect 10870 10248 10876 10260
rect 9434 10220 10876 10248
rect 9434 10217 9446 10220
rect 9388 10211 9446 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 22186 10248 22192 10260
rect 10980 10220 22192 10248
rect 4062 10180 4068 10192
rect 3252 10152 4068 10180
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 8662 10180 8668 10192
rect 8128 10152 8668 10180
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2958 10112 2964 10124
rect 1719 10084 2964 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2958 10072 2964 10084
rect 3016 10112 3022 10124
rect 4525 10115 4583 10121
rect 3016 10084 4016 10112
rect 3016 10072 3022 10084
rect 3988 10056 4016 10084
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 5994 10112 6000 10124
rect 4571 10084 6000 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 8128 10112 8156 10152
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 10410 10140 10416 10192
rect 10468 10180 10474 10192
rect 10980 10180 11008 10220
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 22741 10251 22799 10257
rect 22741 10217 22753 10251
rect 22787 10248 22799 10251
rect 23014 10248 23020 10260
rect 22787 10220 23020 10248
rect 22787 10217 22799 10220
rect 22741 10211 22799 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23198 10208 23204 10260
rect 23256 10248 23262 10260
rect 23385 10251 23443 10257
rect 23385 10248 23397 10251
rect 23256 10220 23397 10248
rect 23256 10208 23262 10220
rect 23385 10217 23397 10220
rect 23431 10217 23443 10251
rect 23385 10211 23443 10217
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24673 10251 24731 10257
rect 24673 10248 24685 10251
rect 24268 10220 24685 10248
rect 24268 10208 24274 10220
rect 24673 10217 24685 10220
rect 24719 10217 24731 10251
rect 25314 10248 25320 10260
rect 25275 10220 25320 10248
rect 24673 10211 24731 10217
rect 25314 10208 25320 10220
rect 25372 10208 25378 10260
rect 34885 10251 34943 10257
rect 34885 10217 34897 10251
rect 34931 10248 34943 10251
rect 36078 10248 36084 10260
rect 34931 10220 36084 10248
rect 34931 10217 34943 10220
rect 34885 10211 34943 10217
rect 36078 10208 36084 10220
rect 36136 10208 36142 10260
rect 10468 10152 11008 10180
rect 10468 10140 10474 10152
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13357 10183 13415 10189
rect 13357 10180 13369 10183
rect 13228 10152 13369 10180
rect 13228 10140 13234 10152
rect 13357 10149 13369 10152
rect 13403 10180 13415 10183
rect 13722 10180 13728 10192
rect 13403 10152 13728 10180
rect 13403 10149 13415 10152
rect 13357 10143 13415 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 23106 10180 23112 10192
rect 16908 10152 23112 10180
rect 16908 10140 16914 10152
rect 23106 10140 23112 10152
rect 23164 10140 23170 10192
rect 23290 10140 23296 10192
rect 23348 10180 23354 10192
rect 23348 10152 24900 10180
rect 23348 10140 23354 10152
rect 6871 10084 8156 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8260 10084 9137 10112
rect 8260 10072 8266 10084
rect 9125 10081 9137 10084
rect 9171 10112 9183 10115
rect 11054 10112 11060 10124
rect 9171 10084 11060 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 11054 10072 11060 10084
rect 11112 10112 11118 10124
rect 11609 10115 11667 10121
rect 11609 10112 11621 10115
rect 11112 10084 11621 10112
rect 11112 10072 11118 10084
rect 11609 10081 11621 10084
rect 11655 10081 11667 10115
rect 11882 10112 11888 10124
rect 11843 10084 11888 10112
rect 11609 10075 11667 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 17218 10112 17224 10124
rect 13280 10084 17224 10112
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 4028 10016 4261 10044
rect 4028 10004 4034 10016
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6564 9976 6592 10007
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8570 10044 8576 10056
rect 8352 10016 8576 10044
rect 8352 10004 8358 10016
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 10744 10016 11284 10044
rect 10744 10004 10750 10016
rect 6730 9976 6736 9988
rect 3174 9948 4476 9976
rect 4448 9908 4476 9948
rect 5920 9948 6500 9976
rect 6564 9948 6736 9976
rect 5920 9908 5948 9948
rect 4448 9880 5948 9908
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6086 9908 6092 9920
rect 6043 9880 6092 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 6086 9868 6092 9880
rect 6144 9908 6150 9920
rect 6270 9908 6276 9920
rect 6144 9880 6276 9908
rect 6144 9868 6150 9880
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 6472 9908 6500 9948
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 7282 9936 7288 9988
rect 7340 9936 7346 9988
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8168 9948 9890 9976
rect 8168 9936 8174 9948
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 11149 9979 11207 9985
rect 11149 9976 11161 9979
rect 11020 9948 11161 9976
rect 11020 9936 11026 9948
rect 11149 9945 11161 9948
rect 11195 9945 11207 9979
rect 11256 9976 11284 10016
rect 11256 9948 12374 9976
rect 11149 9939 11207 9945
rect 13280 9908 13308 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10112 17739 10115
rect 17862 10112 17868 10124
rect 17727 10084 17868 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18874 10112 18880 10124
rect 18012 10084 18880 10112
rect 18012 10072 18018 10084
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19518 10112 19524 10124
rect 19479 10084 19524 10112
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19668 10084 19809 10112
rect 19668 10072 19674 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 20990 10112 20996 10124
rect 20951 10084 20996 10112
rect 19797 10075 19855 10081
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 22848 10084 24624 10112
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 16482 10044 16488 10056
rect 15686 10016 16488 10044
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 16724 10016 16957 10044
rect 16724 10004 16730 10016
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 20806 10044 20812 10056
rect 17092 10016 17540 10044
rect 20767 10016 20812 10044
rect 17092 10004 17098 10016
rect 14553 9979 14611 9985
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14826 9976 14832 9988
rect 14599 9948 14832 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 17310 9976 17316 9988
rect 15856 9948 17316 9976
rect 6472 9880 13308 9908
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 15856 9908 15884 9948
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 17512 9976 17540 10016
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 22186 10004 22192 10056
rect 22244 10044 22250 10056
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 22244 10016 22293 10044
rect 22244 10004 22250 10016
rect 22281 10013 22293 10016
rect 22327 10044 22339 10047
rect 22370 10044 22376 10056
rect 22327 10016 22376 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22848 9988 22876 10084
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10044 22983 10047
rect 23474 10044 23480 10056
rect 22971 10016 23480 10044
rect 22971 10013 22983 10016
rect 22925 10007 22983 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10044 23627 10047
rect 24026 10044 24032 10056
rect 23615 10016 24032 10044
rect 23615 10013 23627 10016
rect 23569 10007 23627 10013
rect 17773 9979 17831 9985
rect 17773 9976 17785 9979
rect 17512 9948 17785 9976
rect 17773 9945 17785 9948
rect 17819 9945 17831 9979
rect 17773 9939 17831 9945
rect 19606 9979 19664 9985
rect 19606 9945 19618 9979
rect 19652 9945 19664 9979
rect 19606 9939 19664 9945
rect 14516 9880 15884 9908
rect 16025 9911 16083 9917
rect 14516 9868 14522 9880
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16206 9908 16212 9920
rect 16071 9880 16212 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9908 17095 9911
rect 17586 9908 17592 9920
rect 17083 9880 17592 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 17586 9868 17592 9880
rect 17644 9908 17650 9920
rect 17862 9908 17868 9920
rect 17644 9880 17868 9908
rect 17644 9868 17650 9880
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19628 9908 19656 9939
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 22830 9976 22836 9988
rect 19944 9948 22836 9976
rect 19944 9936 19950 9948
rect 22830 9936 22836 9948
rect 22888 9936 22894 9988
rect 23106 9936 23112 9988
rect 23164 9976 23170 9988
rect 23584 9976 23612 10007
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24596 10053 24624 10084
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10013 24639 10047
rect 24872 10044 24900 10152
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 24872 10016 25237 10044
rect 24581 10007 24639 10013
rect 25225 10013 25237 10016
rect 25271 10044 25283 10047
rect 26050 10044 26056 10056
rect 25271 10016 26056 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 28902 10004 28908 10056
rect 28960 10044 28966 10056
rect 34333 10047 34391 10053
rect 34333 10044 34345 10047
rect 28960 10016 34345 10044
rect 28960 10004 28966 10016
rect 34333 10013 34345 10016
rect 34379 10013 34391 10047
rect 35066 10044 35072 10056
rect 35027 10016 35072 10044
rect 34333 10007 34391 10013
rect 35066 10004 35072 10016
rect 35124 10004 35130 10056
rect 23164 9948 23612 9976
rect 23164 9936 23170 9948
rect 21450 9908 21456 9920
rect 19484 9880 19656 9908
rect 21411 9880 21456 9908
rect 19484 9868 19490 9880
rect 21450 9868 21456 9880
rect 21508 9868 21514 9920
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 23934 9908 23940 9920
rect 22143 9880 23940 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 23934 9868 23940 9880
rect 23992 9868 23998 9920
rect 34149 9911 34207 9917
rect 34149 9877 34161 9911
rect 34195 9908 34207 9911
rect 34790 9908 34796 9920
rect 34195 9880 34796 9908
rect 34195 9877 34207 9880
rect 34149 9871 34207 9877
rect 34790 9868 34796 9880
rect 34848 9868 34854 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 4890 9704 4896 9716
rect 4672 9676 4896 9704
rect 4672 9664 4678 9676
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 8478 9704 8484 9716
rect 7576 9676 8484 9704
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2455 9608 3924 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2774 9568 2780 9580
rect 2363 9540 2780 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2774 9528 2780 9540
rect 2832 9568 2838 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2832 9540 2973 9568
rect 2832 9528 2838 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3620 9500 3648 9531
rect 2924 9472 3648 9500
rect 2924 9460 2930 9472
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 3418 9432 3424 9444
rect 1811 9404 3424 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 3418 9392 3424 9404
rect 3476 9392 3482 9444
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3234 9364 3240 9376
rect 3099 9336 3240 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3660 9336 3709 9364
rect 3660 9324 3666 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3896 9364 3924 9608
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 7576 9636 7604 9676
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 8665 9707 8723 9713
rect 8665 9673 8677 9707
rect 8711 9704 8723 9707
rect 16850 9704 16856 9716
rect 8711 9676 16856 9704
rect 8711 9673 8723 9676
rect 8665 9667 8723 9673
rect 4120 9608 5014 9636
rect 5828 9608 7604 9636
rect 4120 9596 4126 9608
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4028 9472 4261 9500
rect 4028 9460 4034 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5718 9500 5724 9512
rect 4571 9472 5724 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 5828 9364 5856 9608
rect 7650 9596 7656 9648
rect 7708 9596 7714 9648
rect 9416 9645 9444 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 18414 9704 18420 9716
rect 17828 9676 18420 9704
rect 17828 9664 17834 9676
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19076 9676 19380 9704
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9605 9459 9639
rect 9401 9599 9459 9605
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 12342 9636 12348 9648
rect 11195 9608 12348 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 13814 9636 13820 9648
rect 13478 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 13998 9636 14004 9648
rect 13959 9608 14004 9636
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14737 9639 14795 9645
rect 14737 9605 14749 9639
rect 14783 9636 14795 9639
rect 14826 9636 14832 9648
rect 14783 9608 14832 9636
rect 14783 9605 14795 9608
rect 14737 9599 14795 9605
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 16114 9596 16120 9648
rect 16172 9636 16178 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 16172 9608 17049 9636
rect 16172 9596 16178 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 19076 9636 19104 9676
rect 19242 9636 19248 9648
rect 17037 9599 17095 9605
rect 18340 9608 19104 9636
rect 19203 9608 19248 9636
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 11238 9568 11244 9580
rect 10534 9540 11244 9568
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 5994 9500 6000 9512
rect 5955 9472 6000 9500
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6788 9472 6929 9500
rect 6788 9460 6794 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 8220 9500 8248 9528
rect 7239 9472 8248 9500
rect 9125 9503 9183 9509
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 6822 9432 6828 9444
rect 5960 9404 6828 9432
rect 5960 9392 5966 9404
rect 6822 9392 6828 9404
rect 6880 9392 6886 9444
rect 3896 9336 5856 9364
rect 6932 9364 6960 9463
rect 9140 9364 9168 9463
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11992 9500 12020 9531
rect 11112 9472 12020 9500
rect 12253 9503 12311 9509
rect 11112 9460 11118 9472
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 13998 9500 14004 9512
rect 12299 9472 14004 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14332 9472 14473 9500
rect 14332 9460 14338 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 15746 9500 15752 9512
rect 14461 9463 14519 9469
rect 14568 9472 15752 9500
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 11698 9432 11704 9444
rect 11204 9404 11704 9432
rect 11204 9392 11210 9404
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 14568 9432 14596 9472
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 13872 9404 14596 9432
rect 15856 9432 15884 9554
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 16080 9472 16221 9500
rect 16080 9460 16086 9472
rect 16209 9469 16221 9472
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16632 9472 16957 9500
rect 16632 9460 16638 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 18340 9500 18368 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19352 9636 19380 9676
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20438 9704 20444 9716
rect 20128 9676 20444 9704
rect 20128 9664 20134 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20864 9676 20913 9704
rect 20864 9664 20870 9676
rect 20901 9673 20913 9676
rect 20947 9673 20959 9707
rect 20901 9667 20959 9673
rect 22186 9636 22192 9648
rect 19352 9608 22192 9636
rect 22186 9596 22192 9608
rect 22244 9596 22250 9648
rect 22462 9636 22468 9648
rect 22423 9608 22468 9636
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 23937 9639 23995 9645
rect 23937 9636 23949 9639
rect 23256 9608 23949 9636
rect 23256 9596 23262 9608
rect 23937 9605 23949 9608
rect 23983 9636 23995 9639
rect 27525 9639 27583 9645
rect 23983 9608 27476 9636
rect 23983 9605 23995 9608
rect 23937 9599 23995 9605
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20441 9571 20499 9577
rect 20441 9568 20453 9571
rect 20128 9540 20453 9568
rect 20128 9528 20134 9540
rect 20441 9537 20453 9540
rect 20487 9537 20499 9571
rect 22370 9568 22376 9580
rect 22331 9540 22376 9568
rect 20441 9531 20499 9537
rect 22370 9528 22376 9540
rect 22428 9528 22434 9580
rect 25498 9528 25504 9580
rect 25556 9568 25562 9580
rect 27448 9577 27476 9608
rect 27525 9605 27537 9639
rect 27571 9636 27583 9639
rect 35066 9636 35072 9648
rect 27571 9608 35072 9636
rect 27571 9605 27583 9608
rect 27525 9599 27583 9605
rect 35066 9596 35072 9608
rect 35124 9596 35130 9648
rect 25685 9571 25743 9577
rect 25685 9568 25697 9571
rect 25556 9540 25697 9568
rect 25556 9528 25562 9540
rect 25685 9537 25697 9540
rect 25731 9537 25743 9571
rect 25685 9531 25743 9537
rect 26145 9571 26203 9577
rect 26145 9537 26157 9571
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 16945 9463 17003 9469
rect 17420 9472 18368 9500
rect 18417 9503 18475 9509
rect 17420 9432 17448 9472
rect 18417 9469 18429 9503
rect 18463 9500 18475 9503
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18463 9472 19165 9500
rect 18463 9469 18475 9472
rect 18417 9463 18475 9469
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9469 19487 9503
rect 23290 9500 23296 9512
rect 23251 9472 23296 9500
rect 19429 9463 19487 9469
rect 15856 9404 17448 9432
rect 17497 9435 17555 9441
rect 13872 9392 13878 9404
rect 17497 9401 17509 9435
rect 17543 9432 17555 9435
rect 19444 9432 19472 9463
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 23474 9500 23480 9512
rect 23435 9472 23480 9500
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 24394 9500 24400 9512
rect 24355 9472 24400 9500
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 24578 9500 24584 9512
rect 24539 9472 24584 9500
rect 24578 9460 24584 9472
rect 24636 9460 24642 9512
rect 26160 9432 26188 9531
rect 17543 9404 26188 9432
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 6932 9336 9168 9364
rect 3697 9327 3755 9333
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 12894 9364 12900 9376
rect 10928 9336 12900 9364
rect 10928 9324 10934 9336
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 17954 9364 17960 9376
rect 13412 9336 17960 9364
rect 13412 9324 13418 9336
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 20257 9367 20315 9373
rect 20257 9364 20269 9367
rect 18288 9336 20269 9364
rect 18288 9324 18294 9336
rect 20257 9333 20269 9336
rect 20303 9333 20315 9367
rect 20257 9327 20315 9333
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 24857 9367 24915 9373
rect 24857 9364 24869 9367
rect 23992 9336 24869 9364
rect 23992 9324 23998 9336
rect 24857 9333 24869 9336
rect 24903 9333 24915 9367
rect 25498 9364 25504 9376
rect 25459 9336 25504 9364
rect 24857 9327 24915 9333
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 26237 9367 26295 9373
rect 26237 9333 26249 9367
rect 26283 9364 26295 9367
rect 30190 9364 30196 9376
rect 26283 9336 30196 9364
rect 26283 9333 26295 9336
rect 26237 9327 26295 9333
rect 30190 9324 30196 9336
rect 30248 9324 30254 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 5721 9163 5779 9169
rect 3476 9132 5304 9160
rect 3476 9120 3482 9132
rect 3602 9052 3608 9104
rect 3660 9052 3666 9104
rect 5276 9092 5304 9132
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 9401 9163 9459 9169
rect 5767 9132 9352 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 6546 9092 6552 9104
rect 5276 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 9324 9092 9352 9132
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 9674 9160 9680 9172
rect 9447 9132 9680 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11412 9163 11470 9169
rect 9784 9132 11291 9160
rect 9784 9092 9812 9132
rect 9324 9064 9812 9092
rect 2866 9024 2872 9036
rect 1964 8996 2872 9024
rect 1964 8965 1992 8996
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 3418 9024 3424 9036
rect 2924 8996 3424 9024
rect 2924 8984 2930 8996
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 3620 9024 3648 9052
rect 7101 9027 7159 9033
rect 3620 8996 5580 9024
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2774 8956 2780 8968
rect 2639 8928 2780 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 3050 8888 3056 8900
rect 1360 8860 3056 8888
rect 1360 8848 1366 8860
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3252 8888 3280 8919
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 3970 8956 3976 8968
rect 3660 8928 3976 8956
rect 3660 8916 3666 8928
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4249 8891 4307 8897
rect 3252 8860 4200 8888
rect 4172 8832 4200 8860
rect 4249 8857 4261 8891
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2464 8792 2697 8820
rect 2464 8780 2470 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 2924 8792 3341 8820
rect 2924 8780 2930 8792
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3329 8783 3387 8789
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 4264 8820 4292 8851
rect 5258 8820 5264 8832
rect 4264 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5368 8820 5396 8942
rect 5552 8888 5580 8996
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 10962 9024 10968 9036
rect 7147 8996 10968 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11112 8996 11161 9024
rect 11112 8984 11118 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11263 9024 11291 9132
rect 11412 9129 11424 9163
rect 11458 9160 11470 9163
rect 11882 9160 11888 9172
rect 11458 9132 11888 9160
rect 11458 9129 11470 9132
rect 11412 9123 11470 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 16114 9160 16120 9172
rect 12768 9132 16120 9160
rect 12768 9120 12774 9132
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16448 9132 18184 9160
rect 16448 9120 16454 9132
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 13262 9092 13268 9104
rect 12492 9064 13268 9092
rect 12492 9052 12498 9064
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 14090 9052 14096 9104
rect 14148 9092 14154 9104
rect 14366 9092 14372 9104
rect 14148 9064 14372 9092
rect 14148 9052 14154 9064
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 18049 9095 18107 9101
rect 18049 9061 18061 9095
rect 18095 9061 18107 9095
rect 18156 9092 18184 9132
rect 18598 9120 18604 9172
rect 18656 9160 18662 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18656 9132 18705 9160
rect 18656 9120 18662 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 19426 9160 19432 9172
rect 19387 9132 19432 9160
rect 18693 9123 18751 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 22005 9163 22063 9169
rect 20404 9132 21772 9160
rect 20404 9120 20410 9132
rect 21634 9092 21640 9104
rect 18156 9064 21640 9092
rect 18049 9055 18107 9061
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 11263 8996 14657 9024
rect 11149 8987 11207 8993
rect 14645 8993 14657 8996
rect 14691 9024 14703 9027
rect 18064 9024 18092 9055
rect 21634 9052 21640 9064
rect 21692 9052 21698 9104
rect 21744 9092 21772 9132
rect 22005 9129 22017 9163
rect 22051 9160 22063 9163
rect 22094 9160 22100 9172
rect 22051 9132 22100 9160
rect 22051 9129 22063 9132
rect 22005 9123 22063 9129
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22649 9163 22707 9169
rect 22649 9129 22661 9163
rect 22695 9160 22707 9163
rect 22695 9132 23428 9160
rect 22695 9129 22707 9132
rect 22649 9123 22707 9129
rect 23400 9092 23428 9132
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 25225 9163 25283 9169
rect 25225 9160 25237 9163
rect 23532 9132 25237 9160
rect 23532 9120 23538 9132
rect 25225 9129 25237 9132
rect 25271 9129 25283 9163
rect 25225 9123 25283 9129
rect 24762 9092 24768 9104
rect 21744 9064 23336 9092
rect 23400 9064 24768 9092
rect 14691 8996 16896 9024
rect 18064 8996 18920 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5776 8928 6193 8956
rect 5776 8916 5782 8928
rect 6181 8925 6193 8928
rect 6227 8956 6239 8959
rect 6546 8956 6552 8968
rect 6227 8928 6552 8956
rect 6227 8925 6239 8928
rect 6181 8919 6239 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6788 8928 6837 8956
rect 6788 8916 6794 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 9582 8956 9588 8968
rect 9543 8928 9588 8956
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9824 8928 10057 8956
rect 9824 8916 9830 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10226 8956 10232 8968
rect 10187 8928 10232 8956
rect 10045 8919 10103 8925
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13538 8956 13544 8968
rect 13228 8928 13544 8956
rect 13228 8916 13234 8928
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 8754 8888 8760 8900
rect 5552 8860 7512 8888
rect 5810 8820 5816 8832
rect 5368 8792 5816 8820
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 7374 8820 7380 8832
rect 6319 8792 7380 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7484 8820 7512 8860
rect 8588 8860 8760 8888
rect 8386 8820 8392 8832
rect 7484 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8588 8829 8616 8860
rect 8754 8848 8760 8860
rect 8812 8888 8818 8900
rect 9416 8888 9444 8916
rect 8812 8860 9444 8888
rect 10689 8891 10747 8897
rect 8812 8848 8818 8860
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 11146 8888 11152 8900
rect 10735 8860 11152 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 11532 8860 11914 8888
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 11532 8820 11560 8860
rect 12894 8820 12900 8832
rect 9364 8792 11560 8820
rect 12855 8792 12900 8820
rect 9364 8780 9370 8792
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13228 8792 13553 8820
rect 13228 8780 13234 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13740 8820 13768 8919
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 14332 8928 14381 8956
rect 14332 8916 14338 8928
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 16390 8956 16396 8968
rect 15778 8928 16396 8956
rect 14369 8919 14427 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 16574 8956 16580 8968
rect 16535 8928 16580 8956
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16758 8956 16764 8968
rect 16719 8928 16764 8956
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16868 8956 16896 8996
rect 18892 8965 18920 8996
rect 19058 8984 19064 9036
rect 19116 9024 19122 9036
rect 21545 9027 21603 9033
rect 19116 8996 20300 9024
rect 19116 8984 19122 8996
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 16868 8928 18245 8956
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 20070 8956 20076 8968
rect 19659 8928 20076 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 17494 8888 17500 8900
rect 17052 8860 17500 8888
rect 17052 8820 17080 8860
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 18248 8888 18276 8919
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 20272 8965 20300 8996
rect 21545 8993 21557 9027
rect 21591 9024 21603 9027
rect 21591 8996 22784 9024
rect 21591 8993 21603 8996
rect 21545 8987 21603 8993
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20714 8956 20720 8968
rect 20675 8928 20720 8956
rect 20257 8919 20315 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8956 21419 8959
rect 22462 8956 22468 8968
rect 21407 8928 22468 8956
rect 21407 8925 21419 8928
rect 21361 8919 21419 8925
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 22370 8888 22376 8900
rect 18248 8860 22376 8888
rect 22370 8848 22376 8860
rect 22428 8848 22434 8900
rect 22756 8888 22784 8996
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 23308 8965 23336 9064
rect 24762 9052 24768 9064
rect 24820 9052 24826 9104
rect 23293 8959 23351 8965
rect 22888 8928 22933 8956
rect 22888 8916 22894 8928
rect 23293 8925 23305 8959
rect 23339 8925 23351 8959
rect 23293 8919 23351 8925
rect 24486 8916 24492 8968
rect 24544 8956 24550 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24544 8928 24593 8956
rect 24544 8916 24550 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24670 8916 24676 8968
rect 24728 8956 24734 8968
rect 25409 8959 25467 8965
rect 25409 8956 25421 8959
rect 24728 8928 25421 8956
rect 24728 8916 24734 8928
rect 25409 8925 25421 8928
rect 25455 8925 25467 8959
rect 25409 8919 25467 8925
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 34848 8928 38025 8956
rect 34848 8916 34854 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 23385 8891 23443 8897
rect 23385 8888 23397 8891
rect 22756 8860 23397 8888
rect 23385 8857 23397 8860
rect 23431 8857 23443 8891
rect 23385 8851 23443 8857
rect 17218 8820 17224 8832
rect 13740 8792 17080 8820
rect 17179 8792 17224 8820
rect 13541 8783 13599 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 20809 8823 20867 8829
rect 20809 8820 20821 8823
rect 17368 8792 20821 8820
rect 17368 8780 17374 8792
rect 20809 8789 20821 8792
rect 20855 8789 20867 8823
rect 20809 8783 20867 8789
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 23532 8792 24685 8820
rect 23532 8780 23538 8792
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 24673 8783 24731 8789
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 4062 8616 4068 8628
rect 1811 8588 4068 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 6454 8616 6460 8628
rect 4212 8588 6460 8616
rect 4212 8576 4218 8588
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7156 8588 9168 8616
rect 7156 8576 7162 8588
rect 4982 8548 4988 8560
rect 4462 8520 4988 8548
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 7650 8548 7656 8560
rect 5316 8520 7656 8548
rect 5316 8508 5322 8520
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 9140 8548 9168 8588
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 12434 8616 12440 8628
rect 9456 8588 12440 8616
rect 9456 8576 9462 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 16117 8619 16175 8625
rect 16117 8585 16129 8619
rect 16163 8616 16175 8619
rect 17034 8616 17040 8628
rect 16163 8588 17040 8616
rect 16163 8585 16175 8588
rect 16117 8579 16175 8585
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 19242 8616 19248 8628
rect 17420 8588 18920 8616
rect 19203 8588 19248 8616
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 9140 8520 9321 8548
rect 9309 8517 9321 8520
rect 9355 8517 9367 8551
rect 9309 8511 9367 8517
rect 11900 8520 12434 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 2866 8480 2872 8492
rect 2547 8452 2872 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 1688 8412 1716 8443
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 2958 8412 2964 8424
rect 1688 8384 2820 8412
rect 2919 8384 2964 8412
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 2317 8347 2375 8353
rect 2317 8344 2329 8347
rect 1636 8316 2329 8344
rect 1636 8304 1642 8316
rect 2317 8313 2329 8316
rect 2363 8313 2375 8347
rect 2317 8307 2375 8313
rect 2792 8276 2820 8384
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 3068 8384 3249 8412
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3068 8344 3096 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 5184 8412 5212 8443
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5776 8452 5825 8480
rect 5776 8440 5782 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 7006 8480 7012 8492
rect 5813 8443 5871 8449
rect 5920 8452 7012 8480
rect 3752 8384 5212 8412
rect 5261 8415 5319 8421
rect 3752 8372 3758 8384
rect 5261 8381 5273 8415
rect 5307 8412 5319 8415
rect 5442 8412 5448 8424
rect 5307 8384 5448 8412
rect 5307 8381 5319 8384
rect 5261 8375 5319 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5920 8412 5948 8452
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 11900 8480 11928 8520
rect 5552 8384 5948 8412
rect 2924 8316 3096 8344
rect 2924 8304 2930 8316
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 4709 8347 4767 8353
rect 4709 8344 4721 8347
rect 4580 8316 4721 8344
rect 4580 8304 4586 8316
rect 4709 8313 4721 8316
rect 4755 8313 4767 8347
rect 5552 8344 5580 8384
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6788 8384 7113 8412
rect 6788 8372 6794 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8412 7435 8415
rect 8110 8412 8116 8424
rect 7423 8384 8116 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 4709 8307 4767 8313
rect 4816 8316 5580 8344
rect 3878 8276 3884 8288
rect 2792 8248 3884 8276
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4816 8276 4844 8316
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5684 8316 5917 8344
rect 5684 8304 5690 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 8496 8344 8524 8466
rect 8864 8452 11928 8480
rect 11977 8483 12035 8489
rect 8864 8421 8892 8452
rect 11977 8449 11989 8483
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12158 8480 12164 8492
rect 12115 8452 12164 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 10962 8412 10968 8424
rect 8849 8375 8907 8381
rect 9324 8384 10968 8412
rect 9324 8344 9352 8384
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 8496 8316 9352 8344
rect 5905 8307 5963 8313
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 9456 8316 10609 8344
rect 9456 8304 9462 8316
rect 10597 8313 10609 8316
rect 10643 8344 10655 8347
rect 11146 8344 11152 8356
rect 10643 8316 11152 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11992 8344 12020 8443
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12406 8412 12434 8520
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 12713 8551 12771 8557
rect 12713 8548 12725 8551
rect 12584 8520 12725 8548
rect 12584 8508 12590 8520
rect 12713 8517 12725 8520
rect 12759 8517 12771 8551
rect 12713 8511 12771 8517
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 12986 8548 12992 8560
rect 12851 8520 12992 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13354 8548 13360 8560
rect 13315 8520 13360 8548
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 14366 8548 14372 8560
rect 13464 8520 14372 8548
rect 13464 8412 13492 8520
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 12406 8384 13492 8412
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14458 8412 14464 8424
rect 14139 8384 14464 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 13740 8344 13768 8372
rect 11992 8316 13768 8344
rect 4028 8248 4844 8276
rect 4028 8236 4034 8248
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 13722 8276 13728 8288
rect 5500 8248 13728 8276
rect 5500 8236 5506 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13832 8276 13860 8375
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 15212 8344 15240 8466
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15620 8452 16313 8480
rect 15620 8440 15626 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17310 8480 17316 8492
rect 16991 8452 17316 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 16390 8412 16396 8424
rect 15528 8384 16396 8412
rect 15528 8372 15534 8384
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17420 8412 17448 8588
rect 18230 8548 18236 8560
rect 18191 8520 18236 8548
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18414 8508 18420 8560
rect 18472 8548 18478 8560
rect 18785 8551 18843 8557
rect 18785 8548 18797 8551
rect 18472 8520 18797 8548
rect 18472 8508 18478 8520
rect 18785 8517 18797 8520
rect 18831 8517 18843 8551
rect 18892 8548 18920 8588
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 23198 8616 23204 8628
rect 23159 8588 23204 8616
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 23661 8619 23719 8625
rect 23661 8616 23673 8619
rect 23348 8588 23673 8616
rect 23348 8576 23354 8588
rect 23661 8585 23673 8588
rect 23707 8585 23719 8619
rect 23661 8579 23719 8585
rect 24305 8619 24363 8625
rect 24305 8585 24317 8619
rect 24351 8616 24363 8619
rect 24578 8616 24584 8628
rect 24351 8588 24584 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 24578 8576 24584 8588
rect 24636 8576 24642 8628
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 25004 8588 25053 8616
rect 25004 8576 25010 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 33686 8616 33692 8628
rect 33647 8588 33692 8616
rect 25041 8579 25099 8585
rect 33686 8576 33692 8588
rect 33744 8576 33750 8628
rect 21818 8548 21824 8560
rect 18892 8520 21824 8548
rect 18785 8511 18843 8517
rect 21818 8508 21824 8520
rect 21876 8508 21882 8560
rect 25498 8548 25504 8560
rect 24504 8520 25504 8548
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19208 8452 19441 8480
rect 19208 8440 19214 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 19429 8443 19487 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 24302 8480 24308 8492
rect 21223 8452 24308 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24504 8489 24532 8520
rect 25498 8508 25504 8520
rect 25556 8508 25562 8560
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 24949 8483 25007 8489
rect 24949 8449 24961 8483
rect 24995 8480 25007 8483
rect 29730 8480 29736 8492
rect 24995 8452 29736 8480
rect 24995 8449 25007 8452
rect 24949 8443 25007 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8480 33655 8483
rect 34698 8480 34704 8492
rect 33643 8452 34704 8480
rect 33643 8449 33655 8452
rect 33597 8443 33655 8449
rect 34698 8440 34704 8452
rect 34756 8440 34762 8492
rect 17175 8384 17448 8412
rect 18141 8415 18199 8421
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 18141 8381 18153 8415
rect 18187 8412 18199 8415
rect 19334 8412 19340 8424
rect 18187 8384 19340 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 19444 8384 21281 8412
rect 17310 8344 17316 8356
rect 15212 8316 17172 8344
rect 17271 8316 17316 8344
rect 14274 8276 14280 8288
rect 13832 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 15565 8279 15623 8285
rect 15565 8276 15577 8279
rect 15528 8248 15577 8276
rect 15528 8236 15534 8248
rect 15565 8245 15577 8248
rect 15611 8245 15623 8279
rect 15565 8239 15623 8245
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 17034 8276 17040 8288
rect 16264 8248 17040 8276
rect 16264 8236 16270 8248
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17144 8276 17172 8316
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 17494 8304 17500 8356
rect 17552 8344 17558 8356
rect 19444 8344 19472 8384
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 22554 8412 22560 8424
rect 22515 8384 22560 8412
rect 21269 8375 21327 8381
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 22741 8415 22799 8421
rect 22741 8381 22753 8415
rect 22787 8412 22799 8415
rect 23842 8412 23848 8424
rect 22787 8384 23848 8412
rect 22787 8381 22799 8384
rect 22741 8375 22799 8381
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 17552 8316 19472 8344
rect 17552 8304 17558 8316
rect 17954 8276 17960 8288
rect 17144 8248 17960 8276
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 19150 8276 19156 8288
rect 18840 8248 19156 8276
rect 18840 8236 18846 8248
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 20073 8279 20131 8285
rect 20073 8245 20085 8279
rect 20119 8276 20131 8279
rect 20806 8276 20812 8288
rect 20119 8248 20812 8276
rect 20119 8245 20131 8248
rect 20073 8239 20131 8245
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 5258 8072 5264 8084
rect 2740 8044 5264 8072
rect 2740 8032 2746 8044
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10226 8072 10232 8084
rect 9815 8044 10232 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 16025 8075 16083 8081
rect 10367 8044 15608 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 8113 8007 8171 8013
rect 8113 8004 8125 8007
rect 6748 7976 8125 8004
rect 6748 7948 6776 7976
rect 8113 7973 8125 7976
rect 8159 7973 8171 8007
rect 8113 7967 8171 7973
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 15580 8004 15608 8044
rect 16025 8041 16037 8075
rect 16071 8072 16083 8075
rect 16298 8072 16304 8084
rect 16071 8044 16304 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 20530 8072 20536 8084
rect 16868 8044 20536 8072
rect 16758 8004 16764 8016
rect 12952 7976 14412 8004
rect 15580 7976 16764 8004
rect 12952 7964 12958 7976
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 6730 7936 6736 7948
rect 4295 7908 6736 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 6822 7896 6828 7948
rect 6880 7896 6886 7948
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 14384 7936 14412 7976
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 15010 7936 15016 7948
rect 11011 7908 14320 7936
rect 14384 7908 15016 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 6840 7868 6868 7896
rect 14292 7880 14320 7908
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 16868 7936 16896 8044
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21450 8072 21456 8084
rect 21315 8044 21456 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 21818 8072 21824 8084
rect 21779 8044 21824 8072
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 23842 8072 23848 8084
rect 23803 8044 23848 8072
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 34698 8032 34704 8084
rect 34756 8072 34762 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 34756 8044 38117 8072
rect 34756 8032 34762 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17092 7976 18184 8004
rect 17092 7964 17098 7976
rect 15672 7908 16896 7936
rect 16945 7939 17003 7945
rect 6319 7840 6868 7868
rect 9677 7871 9735 7877
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9858 7868 9864 7880
rect 9723 7840 9864 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9858 7828 9864 7840
rect 9916 7868 9922 7880
rect 10226 7868 10232 7880
rect 9916 7840 10232 7868
rect 9916 7828 9922 7840
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12584 7840 13001 7868
rect 12584 7828 12590 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 13541 7831 13599 7837
rect 1670 7800 1676 7812
rect 1631 7772 1676 7800
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3421 7803 3479 7809
rect 3421 7800 3433 7803
rect 3016 7772 3433 7800
rect 3016 7760 3022 7772
rect 3421 7769 3433 7772
rect 3467 7800 3479 7803
rect 3602 7800 3608 7812
rect 3467 7772 3608 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 4525 7803 4583 7809
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 4614 7800 4620 7812
rect 4571 7772 4620 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 5534 7760 5540 7812
rect 5592 7760 5598 7812
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7769 6883 7803
rect 6825 7763 6883 7769
rect 11248 7803 11306 7809
rect 11248 7769 11260 7803
rect 11294 7769 11306 7803
rect 11248 7763 11306 7769
rect 1688 7732 1716 7760
rect 6840 7732 6868 7763
rect 9398 7732 9404 7744
rect 1688 7704 9404 7732
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 11256 7732 11284 7763
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 13556 7800 13584 7831
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 15672 7854 15700 7908
rect 16945 7905 16957 7939
rect 16991 7936 17003 7939
rect 17402 7936 17408 7948
rect 16991 7908 17408 7936
rect 16991 7905 17003 7908
rect 16945 7899 17003 7905
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 18046 7936 18052 7948
rect 18007 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18156 7936 18184 7976
rect 18598 7964 18604 8016
rect 18656 8004 18662 8016
rect 19242 8004 19248 8016
rect 18656 7976 19248 8004
rect 18656 7964 18662 7976
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 19702 7964 19708 8016
rect 19760 8004 19766 8016
rect 23109 8007 23167 8013
rect 19760 7976 22508 8004
rect 19760 7964 19766 7976
rect 19426 7948 19432 7960
rect 19352 7936 19432 7948
rect 18156 7920 19432 7936
rect 18156 7908 19380 7920
rect 19426 7908 19432 7920
rect 19484 7908 19490 7960
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 20864 7908 20909 7936
rect 20864 7896 20870 7908
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 19334 7868 19340 7880
rect 19306 7828 19340 7868
rect 19392 7828 19398 7880
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 21910 7868 21916 7880
rect 21775 7840 21916 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 12676 7772 14565 7800
rect 12676 7760 12682 7772
rect 14553 7769 14565 7772
rect 14599 7800 14611 7803
rect 14642 7800 14648 7812
rect 14599 7772 14648 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 17034 7760 17040 7812
rect 17092 7800 17098 7812
rect 17586 7800 17592 7812
rect 17092 7772 17137 7800
rect 17499 7772 17592 7800
rect 17092 7760 17098 7772
rect 17586 7760 17592 7772
rect 17644 7800 17650 7812
rect 17644 7772 19012 7800
rect 17644 7760 17650 7772
rect 12158 7732 12164 7744
rect 11256 7704 12164 7732
rect 12158 7692 12164 7704
rect 12216 7732 12222 7744
rect 13262 7732 13268 7744
rect 12216 7704 13268 7732
rect 12216 7692 12222 7704
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 13633 7735 13691 7741
rect 13633 7701 13645 7735
rect 13679 7732 13691 7735
rect 16022 7732 16028 7744
rect 13679 7704 16028 7732
rect 13679 7701 13691 7704
rect 13633 7695 13691 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 18138 7732 18144 7744
rect 16172 7704 18144 7732
rect 16172 7692 16178 7704
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 18690 7732 18696 7744
rect 18651 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 18984 7732 19012 7772
rect 19058 7760 19064 7812
rect 19116 7800 19122 7812
rect 19306 7800 19334 7828
rect 19116 7772 19334 7800
rect 19521 7803 19579 7809
rect 19116 7760 19122 7772
rect 19521 7769 19533 7803
rect 19567 7769 19579 7803
rect 19521 7763 19579 7769
rect 19334 7732 19340 7744
rect 18984 7704 19340 7732
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 19536 7732 19564 7763
rect 19610 7760 19616 7812
rect 19668 7800 19674 7812
rect 20165 7803 20223 7809
rect 19668 7772 19713 7800
rect 19668 7760 19674 7772
rect 20165 7769 20177 7803
rect 20211 7800 20223 7803
rect 20211 7772 20576 7800
rect 20211 7769 20223 7772
rect 20165 7763 20223 7769
rect 20548 7744 20576 7772
rect 20438 7732 20444 7744
rect 19536 7704 20444 7732
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 20640 7732 20668 7831
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22370 7868 22376 7880
rect 22331 7840 22376 7868
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 22480 7868 22508 7976
rect 23109 7973 23121 8007
rect 23155 8004 23167 8007
rect 24670 8004 24676 8016
rect 23155 7976 24676 8004
rect 23155 7973 23167 7976
rect 23109 7967 23167 7973
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 23293 7871 23351 7877
rect 23293 7868 23305 7871
rect 22480 7840 23305 7868
rect 23293 7837 23305 7840
rect 23339 7868 23351 7871
rect 23753 7871 23811 7877
rect 23753 7868 23765 7871
rect 23339 7840 23765 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 23753 7837 23765 7840
rect 23799 7837 23811 7871
rect 23753 7831 23811 7837
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7868 24639 7871
rect 25406 7868 25412 7880
rect 24627 7840 25412 7868
rect 24627 7837 24639 7840
rect 24581 7831 24639 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 22465 7803 22523 7809
rect 22465 7800 22477 7803
rect 21416 7772 22477 7800
rect 21416 7760 21422 7772
rect 22465 7769 22477 7772
rect 22511 7769 22523 7803
rect 22465 7763 22523 7769
rect 24486 7732 24492 7744
rect 20640 7704 24492 7732
rect 24486 7692 24492 7704
rect 24544 7692 24550 7744
rect 24670 7732 24676 7744
rect 24631 7704 24676 7732
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2682 7528 2688 7540
rect 2363 7500 2688 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 7190 7528 7196 7540
rect 3007 7500 7196 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7834 7528 7840 7540
rect 7392 7500 7840 7528
rect 1394 7420 1400 7472
rect 1452 7460 1458 7472
rect 1854 7460 1860 7472
rect 1452 7432 1860 7460
rect 1452 7420 1458 7432
rect 1854 7420 1860 7432
rect 1912 7420 1918 7472
rect 2240 7432 3464 7460
rect 2240 7401 2268 7432
rect 3436 7404 3464 7432
rect 3694 7420 3700 7472
rect 3752 7460 3758 7472
rect 7009 7463 7067 7469
rect 3752 7432 4922 7460
rect 3752 7420 3758 7432
rect 7009 7429 7021 7463
rect 7055 7460 7067 7463
rect 7392 7460 7420 7500
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 12618 7528 12624 7540
rect 8527 7500 12624 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13173 7531 13231 7537
rect 12768 7500 13124 7528
rect 12768 7488 12774 7500
rect 9398 7460 9404 7472
rect 7055 7432 7420 7460
rect 9359 7432 9404 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 9398 7420 9404 7432
rect 9456 7420 9462 7472
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11054 7460 11060 7472
rect 11011 7432 11060 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 12526 7460 12532 7472
rect 11808 7432 12532 7460
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 1627 7364 2237 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2832 7364 2881 7392
rect 2832 7352 2838 7364
rect 2869 7361 2881 7364
rect 2915 7392 2927 7395
rect 2958 7392 2964 7404
rect 2915 7364 2964 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3476 7364 3525 7392
rect 3476 7352 3482 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3660 7364 4169 7392
rect 3660 7352 3666 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 4157 7355 4215 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 10870 7392 10876 7404
rect 8142 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 5166 7324 5172 7336
rect 4479 7296 5172 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5902 7324 5908 7336
rect 5815 7296 5908 7324
rect 5902 7284 5908 7296
rect 5960 7324 5966 7336
rect 7466 7324 7472 7336
rect 5960 7296 7472 7324
rect 5960 7284 5966 7296
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 11698 7324 11704 7336
rect 9732 7296 11704 7324
rect 9732 7284 9738 7296
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 4062 7256 4068 7268
rect 1719 7228 4068 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 11808 7265 11836 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12894 7392 12900 7404
rect 12023 7364 12900 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13096 7401 13124 7500
rect 13173 7497 13185 7531
rect 13219 7528 13231 7531
rect 13219 7500 17080 7528
rect 13219 7497 13231 7500
rect 13173 7491 13231 7497
rect 13998 7460 14004 7472
rect 13959 7432 14004 7460
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 16482 7460 16488 7472
rect 15226 7432 16488 7460
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 17052 7469 17080 7500
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 18288 7500 20177 7528
rect 18288 7488 18294 7500
rect 20165 7497 20177 7500
rect 20211 7497 20223 7531
rect 20165 7491 20223 7497
rect 20438 7488 20444 7540
rect 20496 7528 20502 7540
rect 22278 7528 22284 7540
rect 20496 7500 22284 7528
rect 20496 7488 20502 7500
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 24394 7488 24400 7540
rect 24452 7528 24458 7540
rect 28813 7531 28871 7537
rect 28813 7528 28825 7531
rect 24452 7500 28825 7528
rect 24452 7488 24458 7500
rect 28813 7497 28825 7500
rect 28859 7497 28871 7531
rect 28813 7491 28871 7497
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7429 17095 7463
rect 17037 7423 17095 7429
rect 17589 7463 17647 7469
rect 17589 7429 17601 7463
rect 17635 7460 17647 7463
rect 18598 7460 18604 7472
rect 17635 7432 18604 7460
rect 17635 7429 17647 7432
rect 17589 7423 17647 7429
rect 18598 7420 18604 7432
rect 18656 7420 18662 7472
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 19610 7460 19616 7472
rect 18748 7432 19616 7460
rect 18748 7420 18754 7432
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 21450 7460 21456 7472
rect 19996 7432 21456 7460
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13722 7392 13728 7404
rect 13683 7364 13728 7392
rect 13081 7355 13139 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 16574 7392 16580 7404
rect 15212 7364 16580 7392
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 15212 7324 15240 7364
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 18138 7352 18144 7404
rect 18196 7392 18202 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 18196 7364 18245 7392
rect 18196 7352 18202 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7392 19027 7395
rect 19996 7392 20024 7432
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 19015 7364 20024 7392
rect 20073 7395 20131 7401
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 21174 7392 21180 7404
rect 20763 7364 21180 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 15746 7324 15752 7336
rect 12483 7296 15240 7324
rect 15707 7296 15752 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 18322 7324 18328 7336
rect 16991 7296 18328 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 20088 7324 20116 7355
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22922 7392 22928 7404
rect 22883 7364 22928 7392
rect 22005 7355 22063 7361
rect 20898 7324 20904 7336
rect 20088 7296 20904 7324
rect 20898 7284 20904 7296
rect 20956 7324 20962 7336
rect 21818 7324 21824 7336
rect 20956 7296 21824 7324
rect 20956 7284 20962 7296
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 22020 7324 22048 7355
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 23661 7395 23719 7401
rect 23661 7361 23673 7395
rect 23707 7392 23719 7395
rect 28721 7395 28779 7401
rect 23707 7364 27752 7392
rect 23707 7361 23719 7364
rect 23661 7355 23719 7361
rect 23566 7324 23572 7336
rect 22020 7296 23572 7324
rect 23566 7284 23572 7296
rect 23624 7284 23630 7336
rect 23845 7327 23903 7333
rect 23845 7293 23857 7327
rect 23891 7324 23903 7327
rect 24670 7324 24676 7336
rect 23891 7296 24676 7324
rect 23891 7293 23903 7296
rect 23845 7287 23903 7293
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 27724 7324 27752 7364
rect 28721 7361 28733 7395
rect 28767 7392 28779 7395
rect 35802 7392 35808 7404
rect 28767 7364 35808 7392
rect 28767 7361 28779 7364
rect 28721 7355 28779 7361
rect 35802 7352 35808 7364
rect 35860 7352 35866 7404
rect 31938 7324 31944 7336
rect 27724 7296 31944 7324
rect 31938 7284 31944 7296
rect 31996 7284 32002 7336
rect 11793 7259 11851 7265
rect 11793 7225 11805 7259
rect 11839 7225 11851 7259
rect 11793 7219 11851 7225
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 18049 7259 18107 7265
rect 12584 7228 13584 7256
rect 12584 7216 12590 7228
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 5442 7188 5448 7200
rect 3651 7160 5448 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 7558 7188 7564 7200
rect 6052 7160 7564 7188
rect 6052 7148 6058 7160
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 13446 7188 13452 7200
rect 10560 7160 13452 7188
rect 10560 7148 10566 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13556 7188 13584 7228
rect 18049 7225 18061 7259
rect 18095 7256 18107 7259
rect 19426 7256 19432 7268
rect 18095 7228 19432 7256
rect 18095 7225 18107 7228
rect 18049 7219 18107 7225
rect 19426 7216 19432 7228
rect 19484 7216 19490 7268
rect 19610 7216 19616 7268
rect 19668 7256 19674 7268
rect 19668 7228 20944 7256
rect 19668 7216 19674 7228
rect 15746 7188 15752 7200
rect 13556 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 20438 7188 20444 7200
rect 16540 7160 20444 7188
rect 16540 7148 16546 7160
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 20916 7188 20944 7228
rect 20990 7216 20996 7268
rect 21048 7256 21054 7268
rect 22097 7259 22155 7265
rect 22097 7256 22109 7259
rect 21048 7228 22109 7256
rect 21048 7216 21054 7228
rect 22097 7225 22109 7228
rect 22143 7225 22155 7259
rect 22097 7219 22155 7225
rect 23017 7259 23075 7265
rect 23017 7225 23029 7259
rect 23063 7256 23075 7259
rect 26510 7256 26516 7268
rect 23063 7228 26516 7256
rect 23063 7225 23075 7228
rect 23017 7219 23075 7225
rect 26510 7216 26516 7228
rect 26568 7216 26574 7268
rect 23106 7188 23112 7200
rect 20916 7160 23112 7188
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23934 7148 23940 7200
rect 23992 7188 23998 7200
rect 24029 7191 24087 7197
rect 24029 7188 24041 7191
rect 23992 7160 24041 7188
rect 23992 7148 23998 7160
rect 24029 7157 24041 7160
rect 24075 7157 24087 7191
rect 24029 7151 24087 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 5902 6984 5908 6996
rect 3752 6956 5908 6984
rect 3752 6944 3758 6956
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 7088 6987 7146 6993
rect 7088 6953 7100 6987
rect 7134 6984 7146 6987
rect 10134 6984 10140 6996
rect 7134 6956 10140 6984
rect 7134 6953 7146 6956
rect 7088 6947 7146 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10578 6987 10636 6993
rect 10578 6984 10590 6987
rect 10376 6956 10590 6984
rect 10376 6944 10382 6956
rect 10578 6953 10590 6956
rect 10624 6984 10636 6987
rect 12250 6984 12256 6996
rect 10624 6956 12256 6984
rect 10624 6953 10636 6956
rect 10578 6947 10636 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 12952 6956 13553 6984
rect 12952 6944 12958 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14274 6984 14280 6996
rect 13780 6956 14280 6984
rect 13780 6944 13786 6956
rect 14274 6944 14280 6956
rect 14332 6984 14338 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 14332 6956 15577 6984
rect 14332 6944 14338 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 17218 6984 17224 6996
rect 15565 6947 15623 6953
rect 15672 6956 17224 6984
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 6086 6916 6092 6928
rect 5316 6888 6092 6916
rect 5316 6876 5322 6888
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 15102 6916 15108 6928
rect 12492 6888 15108 6916
rect 12492 6876 12498 6888
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 15672 6916 15700 6956
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 22646 6984 22652 6996
rect 17460 6956 22652 6984
rect 17460 6944 17466 6956
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 24486 6944 24492 6996
rect 24544 6984 24550 6996
rect 28445 6987 28503 6993
rect 28445 6984 28457 6987
rect 24544 6956 28457 6984
rect 24544 6944 24550 6956
rect 28445 6953 28457 6956
rect 28491 6953 28503 6987
rect 28445 6947 28503 6953
rect 15212 6888 15700 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1762 6848 1768 6860
rect 1636 6820 1768 6848
rect 1636 6808 1642 6820
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 5718 6848 5724 6860
rect 3292 6820 5580 6848
rect 5631 6820 5724 6848
rect 3292 6808 3298 6820
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3467 6752 3985 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1636 6684 1685 6712
rect 1636 6672 1642 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3436 6644 3464 6743
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 2740 6616 3464 6644
rect 4264 6644 4292 6675
rect 4890 6672 4896 6724
rect 4948 6672 4954 6724
rect 5552 6712 5580 6820
rect 5718 6808 5724 6820
rect 5776 6848 5782 6860
rect 6362 6848 6368 6860
rect 5776 6820 6368 6848
rect 5776 6808 5782 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 8573 6851 8631 6857
rect 7524 6820 8340 6848
rect 7524 6808 7530 6820
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6270 6780 6276 6792
rect 6227 6752 6276 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 8312 6780 8340 6820
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 9214 6848 9220 6860
rect 8619 6820 9220 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9950 6848 9956 6860
rect 9324 6820 9956 6848
rect 9324 6780 9352 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 11054 6848 11060 6860
rect 10367 6820 11060 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 12342 6848 12348 6860
rect 11204 6820 11928 6848
rect 12303 6820 12348 6848
rect 11204 6808 11210 6820
rect 8312 6752 9352 6780
rect 6825 6743 6883 6749
rect 6840 6712 6868 6743
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9456 6752 9689 6780
rect 9456 6740 9462 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 11900 6724 11928 6820
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 14550 6848 14556 6860
rect 12400 6820 14556 6848
rect 12400 6808 12406 6820
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15212 6848 15240 6888
rect 16482 6876 16488 6928
rect 16540 6916 16546 6928
rect 16850 6916 16856 6928
rect 16540 6888 16856 6916
rect 16540 6876 16546 6888
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 17129 6919 17187 6925
rect 17129 6885 17141 6919
rect 17175 6916 17187 6919
rect 17586 6916 17592 6928
rect 17175 6888 17592 6916
rect 17175 6885 17187 6888
rect 17129 6879 17187 6885
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 20990 6916 20996 6928
rect 17696 6888 20996 6916
rect 17696 6860 17724 6888
rect 20990 6876 20996 6888
rect 21048 6876 21054 6928
rect 33597 6919 33655 6925
rect 33597 6916 33609 6919
rect 30392 6888 33609 6916
rect 14700 6820 15240 6848
rect 16577 6851 16635 6857
rect 14700 6808 14706 6820
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 17310 6848 17316 6860
rect 16623 6820 17316 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 17678 6848 17684 6860
rect 17639 6820 17684 6848
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 18322 6848 18328 6860
rect 18283 6820 18328 6848
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 19426 6848 19432 6860
rect 19387 6820 19432 6848
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 20254 6848 20260 6860
rect 19576 6820 20260 6848
rect 19576 6808 19582 6820
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 20548 6820 20760 6848
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13722 6780 13728 6792
rect 13044 6752 13089 6780
rect 13683 6752 13728 6780
rect 13044 6740 13050 6752
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 16206 6780 16212 6792
rect 14056 6752 16212 6780
rect 14056 6740 14062 6752
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6780 17923 6783
rect 19886 6780 19892 6792
rect 17911 6752 19892 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 20548 6789 20576 6820
rect 20732 6790 20760 6820
rect 22462 6808 22468 6860
rect 22520 6848 22526 6860
rect 22520 6820 25176 6848
rect 22520 6808 22526 6820
rect 20533 6783 20591 6789
rect 20533 6749 20545 6783
rect 20579 6749 20591 6783
rect 20732 6780 20852 6790
rect 21174 6780 21180 6792
rect 20732 6762 21180 6780
rect 20824 6752 21180 6762
rect 20533 6743 20591 6749
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21818 6740 21824 6792
rect 21876 6780 21882 6792
rect 22005 6783 22063 6789
rect 22005 6780 22017 6783
rect 21876 6752 22017 6780
rect 21876 6740 21882 6752
rect 22005 6749 22017 6752
rect 22051 6749 22063 6783
rect 22646 6780 22652 6792
rect 22607 6752 22652 6780
rect 22005 6743 22063 6749
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 23106 6780 23112 6792
rect 23067 6752 23112 6780
rect 23106 6740 23112 6752
rect 23164 6740 23170 6792
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 23937 6783 23995 6789
rect 23440 6752 23888 6780
rect 23440 6740 23446 6752
rect 7006 6712 7012 6724
rect 5552 6684 6776 6712
rect 6840 6684 7012 6712
rect 5258 6644 5264 6656
rect 4264 6616 5264 6644
rect 2740 6604 2746 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6748 6644 6776 6684
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7248 6684 7590 6712
rect 7248 6672 7254 6684
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8444 6684 9996 6712
rect 8444 6672 8450 6684
rect 9490 6644 9496 6656
rect 6748 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 9858 6644 9864 6656
rect 9815 6616 9864 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 9968 6644 9996 6684
rect 10704 6684 11086 6712
rect 10704 6644 10732 6684
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 14277 6715 14335 6721
rect 14277 6712 14289 6715
rect 11940 6684 14289 6712
rect 11940 6672 11946 6684
rect 14277 6681 14289 6684
rect 14323 6681 14335 6715
rect 14277 6675 14335 6681
rect 14918 6672 14924 6724
rect 14976 6712 14982 6724
rect 15838 6712 15844 6724
rect 14976 6684 15844 6712
rect 14976 6672 14982 6684
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 16574 6672 16580 6724
rect 16632 6712 16638 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16632 6684 16681 6712
rect 16632 6672 16638 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 20162 6712 20168 6724
rect 16669 6675 16727 6681
rect 18800 6684 20168 6712
rect 9968 6616 10732 6644
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 12250 6644 12256 6656
rect 10928 6616 12256 6644
rect 10928 6604 10934 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 16114 6644 16120 6656
rect 12768 6616 16120 6644
rect 12768 6604 12774 6616
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 18800 6644 18828 6684
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 18196 6616 18828 6644
rect 18196 6604 18202 6616
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 20254 6644 20260 6656
rect 19024 6616 20260 6644
rect 19024 6604 19030 6616
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 20680 6616 20725 6644
rect 20680 6604 20686 6616
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 21269 6647 21327 6653
rect 21269 6644 21281 6647
rect 20956 6616 21281 6644
rect 20956 6604 20962 6616
rect 21269 6613 21281 6616
rect 21315 6613 21327 6647
rect 21269 6607 21327 6613
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 21821 6647 21879 6653
rect 21821 6644 21833 6647
rect 21416 6616 21833 6644
rect 21416 6604 21422 6616
rect 21821 6613 21833 6616
rect 21867 6613 21879 6647
rect 21821 6607 21879 6613
rect 21910 6604 21916 6656
rect 21968 6644 21974 6656
rect 22465 6647 22523 6653
rect 22465 6644 22477 6647
rect 21968 6616 22477 6644
rect 21968 6604 21974 6616
rect 22465 6613 22477 6616
rect 22511 6613 22523 6647
rect 23198 6644 23204 6656
rect 23159 6616 23204 6644
rect 22465 6607 22523 6613
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 23753 6647 23811 6653
rect 23753 6644 23765 6647
rect 23348 6616 23765 6644
rect 23348 6604 23354 6616
rect 23753 6613 23765 6616
rect 23799 6613 23811 6647
rect 23860 6644 23888 6752
rect 23937 6749 23949 6783
rect 23983 6780 23995 6783
rect 24026 6780 24032 6792
rect 23983 6752 24032 6780
rect 23983 6749 23995 6752
rect 23937 6743 23995 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 25148 6712 25176 6820
rect 28353 6783 28411 6789
rect 28353 6749 28365 6783
rect 28399 6780 28411 6783
rect 30282 6780 30288 6792
rect 28399 6752 30288 6780
rect 28399 6749 28411 6752
rect 28353 6743 28411 6749
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 30392 6712 30420 6888
rect 33597 6885 33609 6888
rect 33643 6885 33655 6919
rect 33597 6879 33655 6885
rect 33505 6783 33563 6789
rect 33505 6749 33517 6783
rect 33551 6780 33563 6783
rect 36354 6780 36360 6792
rect 33551 6752 36360 6780
rect 33551 6749 33563 6752
rect 33505 6743 33563 6749
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 36449 6783 36507 6789
rect 36449 6749 36461 6783
rect 36495 6749 36507 6783
rect 36449 6743 36507 6749
rect 25148 6684 30420 6712
rect 36464 6644 36492 6743
rect 23860 6616 36492 6644
rect 36541 6647 36599 6653
rect 23753 6607 23811 6613
rect 36541 6613 36553 6647
rect 36587 6644 36599 6647
rect 38010 6644 38016 6656
rect 36587 6616 38016 6644
rect 36587 6613 36599 6616
rect 36541 6607 36599 6613
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1670 6440 1676 6452
rect 1452 6412 1676 6440
rect 1452 6400 1458 6412
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 2639 6412 2774 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 2746 6372 2774 6412
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 2924 6412 4629 6440
rect 2924 6400 2930 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 4890 6440 4896 6452
rect 4764 6412 4896 6440
rect 4764 6400 4770 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 7006 6440 7012 6452
rect 6564 6412 7012 6440
rect 3602 6372 3608 6384
rect 2746 6344 3608 6372
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 5258 6372 5264 6384
rect 4370 6358 5264 6372
rect 4356 6344 5264 6358
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1762 6304 1768 6316
rect 1627 6276 1768 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 2682 6236 2688 6248
rect 1544 6208 2688 6236
rect 1544 6196 1550 6208
rect 2682 6196 2688 6208
rect 2740 6236 2746 6248
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2740 6208 2881 6236
rect 2740 6196 2746 6208
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 2869 6199 2927 6205
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 4356 6236 4384 6344
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5902 6304 5908 6316
rect 5859 6276 5908 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 3660 6208 4384 6236
rect 3660 6196 3666 6208
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 5184 6168 5212 6267
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 6564 6313 6592 6412
rect 7006 6400 7012 6412
rect 7064 6440 7070 6452
rect 7064 6412 8984 6440
rect 7064 6400 7070 6412
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 6788 6344 7314 6372
rect 6788 6332 6794 6344
rect 8956 6313 8984 6412
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 11790 6440 11796 6452
rect 9916 6412 11796 6440
rect 9916 6400 9922 6412
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 13722 6440 13728 6452
rect 12032 6412 13728 6440
rect 12032 6400 12038 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 14240 6412 14289 6440
rect 14240 6400 14246 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 18601 6443 18659 6449
rect 18601 6440 18613 6443
rect 14608 6412 18613 6440
rect 14608 6400 14614 6412
rect 18601 6409 18613 6412
rect 18647 6409 18659 6443
rect 20254 6440 20260 6452
rect 18601 6403 18659 6409
rect 19168 6412 20260 6440
rect 9214 6372 9220 6384
rect 9175 6344 9220 6372
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9766 6332 9772 6384
rect 9824 6332 9830 6384
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 12894 6372 12900 6384
rect 10560 6344 12900 6372
rect 10560 6332 10566 6344
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13814 6332 13820 6384
rect 13872 6332 13878 6384
rect 15746 6372 15752 6384
rect 15707 6344 15752 6372
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 15930 6332 15936 6384
rect 15988 6372 15994 6384
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 15988 6344 17141 6372
rect 15988 6332 15994 6344
rect 17129 6341 17141 6344
rect 17175 6341 17187 6375
rect 19168 6372 19196 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 21324 6412 21373 6440
rect 21324 6400 21330 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 21361 6403 21419 6409
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 22612 6412 22661 6440
rect 22612 6400 22618 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 18354 6344 19196 6372
rect 19245 6375 19303 6381
rect 17129 6335 17187 6341
rect 19245 6341 19257 6375
rect 19291 6372 19303 6375
rect 19426 6372 19432 6384
rect 19291 6344 19432 6372
rect 19291 6341 19303 6344
rect 19245 6335 19303 6341
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 19797 6375 19855 6381
rect 19797 6341 19809 6375
rect 19843 6372 19855 6375
rect 19978 6372 19984 6384
rect 19843 6344 19984 6372
rect 19843 6341 19855 6344
rect 19797 6335 19855 6341
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 24578 6372 24584 6384
rect 20088 6344 24584 6372
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11790 6304 11796 6316
rect 11747 6276 11796 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 14918 6304 14924 6316
rect 14879 6276 14924 6304
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16482 6304 16488 6316
rect 16347 6276 16488 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 16842 6307 16900 6313
rect 16842 6304 16854 6307
rect 16724 6276 16854 6304
rect 16724 6264 16730 6276
rect 16842 6273 16854 6276
rect 16888 6273 16900 6307
rect 16842 6267 16900 6273
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 20088 6304 20116 6344
rect 24578 6332 24584 6344
rect 24636 6332 24642 6384
rect 20622 6304 20628 6316
rect 19944 6276 20116 6304
rect 20583 6276 20628 6304
rect 19944 6264 19950 6276
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 21269 6307 21327 6313
rect 21269 6304 21281 6307
rect 21232 6276 21281 6304
rect 21232 6264 21238 6276
rect 21269 6273 21281 6276
rect 21315 6273 21327 6307
rect 21269 6267 21327 6273
rect 21450 6264 21456 6316
rect 21508 6304 21514 6316
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 21508 6276 22201 6304
rect 21508 6264 21514 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6304 23351 6307
rect 23474 6304 23480 6316
rect 23339 6276 23480 6304
rect 23339 6273 23351 6276
rect 23293 6267 23351 6273
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 37734 6304 37740 6316
rect 37695 6276 37740 6304
rect 37734 6264 37740 6276
rect 37792 6264 37798 6316
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 6362 6236 6368 6248
rect 5307 6208 6368 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 8662 6236 8668 6248
rect 6871 6208 8668 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9272 6208 10272 6236
rect 9272 6196 9278 6208
rect 6546 6168 6552 6180
rect 5184 6140 6552 6168
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 10244 6168 10272 6208
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10744 6208 10977 6236
rect 10744 6196 10750 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 12526 6236 12532 6248
rect 12487 6208 12532 6236
rect 10965 6199 11023 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 13354 6236 13360 6248
rect 12851 6208 13360 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 16114 6196 16120 6248
rect 16172 6236 16178 6248
rect 16172 6208 18460 6236
rect 16172 6196 16178 6208
rect 11793 6171 11851 6177
rect 11793 6168 11805 6171
rect 7852 6140 8432 6168
rect 10244 6140 11805 6168
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 4706 6100 4712 6112
rect 2648 6072 4712 6100
rect 2648 6060 2654 6072
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6100 5963 6103
rect 7852 6100 7880 6140
rect 8294 6100 8300 6112
rect 5951 6072 7880 6100
rect 8255 6072 8300 6100
rect 5951 6069 5963 6072
rect 5905 6063 5963 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8404 6100 8432 6140
rect 11793 6137 11805 6140
rect 11839 6137 11851 6171
rect 18432 6168 18460 6208
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 18564 6208 19165 6236
rect 18564 6196 18570 6208
rect 19153 6205 19165 6208
rect 19199 6205 19211 6239
rect 21542 6236 21548 6248
rect 19153 6199 19211 6205
rect 19720 6208 21548 6236
rect 19720 6168 19748 6208
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6236 22063 6239
rect 24762 6236 24768 6248
rect 22051 6208 24768 6236
rect 22051 6205 22063 6208
rect 22005 6199 22063 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 37458 6236 37464 6248
rect 37419 6208 37464 6236
rect 37458 6196 37464 6208
rect 37516 6196 37522 6248
rect 20898 6168 20904 6180
rect 11793 6131 11851 6137
rect 13832 6140 16896 6168
rect 18432 6140 19748 6168
rect 19812 6140 20904 6168
rect 9858 6100 9864 6112
rect 8404 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 11974 6100 11980 6112
rect 10836 6072 11980 6100
rect 10836 6060 10842 6072
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 13832 6100 13860 6140
rect 12492 6072 13860 6100
rect 15013 6103 15071 6109
rect 12492 6060 12498 6072
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 16758 6100 16764 6112
rect 15059 6072 16764 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 16868 6100 16896 6140
rect 19812 6100 19840 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 16868 6072 19840 6100
rect 20717 6103 20775 6109
rect 20717 6069 20729 6103
rect 20763 6100 20775 6103
rect 21266 6100 21272 6112
rect 20763 6072 21272 6100
rect 20763 6069 20775 6072
rect 20717 6063 20775 6069
rect 21266 6060 21272 6072
rect 21324 6060 21330 6112
rect 23109 6103 23167 6109
rect 23109 6069 23121 6103
rect 23155 6100 23167 6103
rect 24670 6100 24676 6112
rect 23155 6072 24676 6100
rect 23155 6069 23167 6072
rect 23109 6063 23167 6069
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 4614 5896 4620 5908
rect 3375 5868 4620 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5644 5868 7512 5896
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 2648 5732 3985 5760
rect 2648 5720 2654 5732
rect 3973 5729 3985 5732
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4982 5760 4988 5772
rect 4295 5732 4988 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4982 5720 4988 5732
rect 5040 5760 5046 5772
rect 5644 5760 5672 5868
rect 5721 5831 5779 5837
rect 5721 5797 5733 5831
rect 5767 5828 5779 5831
rect 5994 5828 6000 5840
rect 5767 5800 6000 5828
rect 5767 5797 5779 5800
rect 5721 5791 5779 5797
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 7484 5828 7512 5868
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7892 5868 7941 5896
rect 7892 5856 7898 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 10502 5896 10508 5908
rect 7929 5859 7987 5865
rect 8036 5868 10508 5896
rect 8036 5828 8064 5868
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11480 5868 11713 5896
rect 11480 5856 11486 5868
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 12710 5896 12716 5908
rect 11701 5859 11759 5865
rect 11808 5868 12716 5896
rect 7484 5800 8064 5828
rect 10410 5788 10416 5840
rect 10468 5828 10474 5840
rect 11808 5828 11836 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 15562 5896 15568 5908
rect 12943 5868 15568 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 18233 5899 18291 5905
rect 16540 5868 17816 5896
rect 16540 5856 16546 5868
rect 14090 5828 14096 5840
rect 10468 5800 11836 5828
rect 12406 5800 14096 5828
rect 10468 5788 10474 5800
rect 5040 5732 5672 5760
rect 6181 5763 6239 5769
rect 5040 5720 5046 5732
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 7006 5760 7012 5772
rect 6227 5732 7012 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7248 5732 7696 5760
rect 7248 5720 7254 5732
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 7668 5692 7696 5732
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 7984 5732 9413 5760
rect 7984 5720 7990 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 12406 5760 12434 5800
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 16025 5831 16083 5837
rect 16025 5828 16037 5831
rect 15896 5800 16037 5828
rect 15896 5788 15902 5800
rect 16025 5797 16037 5800
rect 16071 5828 16083 5831
rect 17788 5828 17816 5868
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18414 5896 18420 5908
rect 18279 5868 18420 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 19150 5896 19156 5908
rect 18739 5868 19156 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 19150 5856 19156 5868
rect 19208 5856 19214 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 20404 5868 21925 5896
rect 20404 5856 20410 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 22554 5896 22560 5908
rect 21913 5859 21971 5865
rect 22066 5868 22560 5896
rect 19886 5828 19892 5840
rect 16071 5800 16620 5828
rect 17788 5800 19892 5828
rect 16071 5797 16083 5800
rect 16025 5791 16083 5797
rect 9548 5732 12434 5760
rect 9548 5720 9554 5732
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 14274 5760 14280 5772
rect 12584 5732 14280 5760
rect 12584 5720 12590 5732
rect 14274 5720 14280 5732
rect 14332 5760 14338 5772
rect 16482 5760 16488 5772
rect 14332 5732 16488 5760
rect 14332 5720 14338 5732
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16592 5760 16620 5800
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 20073 5831 20131 5837
rect 20073 5797 20085 5831
rect 20119 5828 20131 5831
rect 22066 5828 22094 5868
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 23750 5856 23756 5908
rect 23808 5896 23814 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23808 5868 23857 5896
rect 23808 5856 23814 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 20119 5800 22094 5828
rect 22204 5800 22692 5828
rect 20119 5797 20131 5800
rect 20073 5791 20131 5797
rect 18046 5760 18052 5772
rect 16592 5732 18052 5760
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 21358 5760 21364 5772
rect 18892 5732 21364 5760
rect 8386 5692 8392 5704
rect 7668 5664 8392 5692
rect 1581 5655 1639 5661
rect 8386 5652 8392 5664
rect 8444 5692 8450 5704
rect 8938 5692 8944 5704
rect 8444 5664 8944 5692
rect 8444 5652 8450 5664
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10928 5664 11161 5692
rect 10928 5652 10934 5664
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 1857 5627 1915 5633
rect 1857 5593 1869 5627
rect 1903 5593 1915 5627
rect 1857 5587 1915 5593
rect 1872 5556 1900 5587
rect 2314 5584 2320 5636
rect 2372 5584 2378 5636
rect 6362 5624 6368 5636
rect 5474 5596 6368 5624
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 6457 5627 6515 5633
rect 6457 5593 6469 5627
rect 6503 5624 6515 5627
rect 8202 5624 8208 5636
rect 6503 5596 6868 5624
rect 7682 5596 8208 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 6638 5556 6644 5568
rect 1872 5528 6644 5556
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6840 5556 6868 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 9490 5624 9496 5636
rect 8312 5596 9496 5624
rect 8312 5556 8340 5596
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 9858 5584 9864 5636
rect 9916 5584 9922 5636
rect 8478 5556 8484 5568
rect 6840 5528 8340 5556
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 10888 5556 10916 5652
rect 11624 5624 11652 5655
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 11974 5692 11980 5704
rect 11848 5664 11980 5692
rect 11848 5652 11854 5664
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5692 12495 5695
rect 12483 5664 12940 5692
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 12912 5624 12940 5664
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 13044 5664 13093 5692
rect 13044 5652 13050 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 18892 5701 18920 5732
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13596 5664 13737 5692
rect 13596 5652 13602 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19392 5664 19441 5692
rect 19392 5652 19398 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19978 5692 19984 5704
rect 19659 5664 19984 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 20530 5692 20536 5704
rect 20443 5664 20536 5692
rect 20530 5652 20536 5664
rect 20588 5692 20594 5704
rect 21174 5692 21180 5704
rect 20588 5664 21180 5692
rect 20588 5652 20594 5664
rect 21174 5652 21180 5664
rect 21232 5692 21238 5704
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 21232 5664 21833 5692
rect 21232 5652 21238 5664
rect 21821 5661 21833 5664
rect 21867 5692 21879 5695
rect 22204 5692 22232 5800
rect 22557 5763 22615 5769
rect 22557 5760 22569 5763
rect 21867 5664 22232 5692
rect 22388 5732 22569 5760
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 11624 5596 12848 5624
rect 12912 5596 13860 5624
rect 8720 5528 10916 5556
rect 12253 5559 12311 5565
rect 8720 5516 8726 5528
rect 12253 5525 12265 5559
rect 12299 5556 12311 5559
rect 12710 5556 12716 5568
rect 12299 5528 12716 5556
rect 12299 5525 12311 5528
rect 12253 5519 12311 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 12820 5556 12848 5596
rect 12894 5556 12900 5568
rect 12820 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 13541 5559 13599 5565
rect 13541 5556 13553 5559
rect 13504 5528 13553 5556
rect 13504 5516 13510 5528
rect 13541 5525 13553 5528
rect 13587 5525 13599 5559
rect 13832 5556 13860 5596
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 14553 5627 14611 5633
rect 14553 5624 14565 5627
rect 13964 5596 14565 5624
rect 13964 5584 13970 5596
rect 14553 5593 14565 5596
rect 14599 5593 14611 5627
rect 15778 5596 16252 5624
rect 14553 5587 14611 5593
rect 15930 5556 15936 5568
rect 13832 5528 15936 5556
rect 13541 5519 13599 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16224 5556 16252 5596
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16761 5627 16819 5633
rect 16761 5624 16773 5627
rect 16356 5596 16773 5624
rect 16356 5584 16362 5596
rect 16761 5593 16773 5596
rect 16807 5593 16819 5627
rect 20806 5624 20812 5636
rect 17986 5596 20812 5624
rect 16761 5587 16819 5593
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 20898 5584 20904 5636
rect 20956 5624 20962 5636
rect 22388 5624 22416 5732
rect 22557 5729 22569 5732
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22664 5692 22692 5800
rect 23014 5692 23020 5704
rect 22511 5664 23020 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 23109 5695 23167 5701
rect 23109 5661 23121 5695
rect 23155 5692 23167 5695
rect 23474 5692 23480 5704
rect 23155 5664 23480 5692
rect 23155 5661 23167 5664
rect 23109 5655 23167 5661
rect 23474 5652 23480 5664
rect 23532 5692 23538 5704
rect 23753 5695 23811 5701
rect 23753 5692 23765 5695
rect 23532 5664 23765 5692
rect 23532 5652 23538 5664
rect 23753 5661 23765 5664
rect 23799 5661 23811 5695
rect 23753 5655 23811 5661
rect 30190 5652 30196 5704
rect 30248 5692 30254 5704
rect 30653 5695 30711 5701
rect 30653 5692 30665 5695
rect 30248 5664 30665 5692
rect 30248 5652 30254 5664
rect 30653 5661 30665 5664
rect 30699 5661 30711 5695
rect 30653 5655 30711 5661
rect 23201 5627 23259 5633
rect 23201 5624 23213 5627
rect 20956 5596 22416 5624
rect 22480 5596 23213 5624
rect 20956 5584 20962 5596
rect 20346 5556 20352 5568
rect 16224 5528 20352 5556
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 20625 5559 20683 5565
rect 20625 5525 20637 5559
rect 20671 5556 20683 5559
rect 20714 5556 20720 5568
rect 20671 5528 20720 5556
rect 20671 5525 20683 5528
rect 20625 5519 20683 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 21082 5516 21088 5568
rect 21140 5556 21146 5568
rect 21269 5559 21327 5565
rect 21269 5556 21281 5559
rect 21140 5528 21281 5556
rect 21140 5516 21146 5528
rect 21269 5525 21281 5528
rect 21315 5525 21327 5559
rect 21269 5519 21327 5525
rect 22002 5516 22008 5568
rect 22060 5556 22066 5568
rect 22480 5556 22508 5596
rect 23201 5593 23213 5596
rect 23247 5593 23259 5627
rect 23201 5587 23259 5593
rect 22060 5528 22508 5556
rect 30469 5559 30527 5565
rect 22060 5516 22066 5528
rect 30469 5525 30481 5559
rect 30515 5556 30527 5559
rect 33042 5556 33048 5568
rect 30515 5528 33048 5556
rect 30515 5525 30527 5528
rect 30469 5519 30527 5525
rect 33042 5516 33048 5528
rect 33100 5516 33106 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 5718 5352 5724 5364
rect 3896 5324 5724 5352
rect 3896 5293 3924 5324
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 7282 5352 7288 5364
rect 6779 5324 7288 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 8202 5352 8208 5364
rect 7800 5324 8208 5352
rect 7800 5312 7806 5324
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9030 5352 9036 5364
rect 8991 5324 9036 5352
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10686 5352 10692 5364
rect 9916 5324 10692 5352
rect 9916 5312 9922 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 11057 5355 11115 5361
rect 11057 5352 11069 5355
rect 11020 5324 11069 5352
rect 11020 5312 11026 5324
rect 11057 5321 11069 5324
rect 11103 5321 11115 5355
rect 11057 5315 11115 5321
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12158 5352 12164 5364
rect 11931 5324 12164 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 13998 5352 14004 5364
rect 13648 5324 14004 5352
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5253 3939 5287
rect 3881 5247 3939 5253
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 7548 5287 7606 5293
rect 7548 5284 7560 5287
rect 7248 5256 7560 5284
rect 7248 5244 7254 5256
rect 7548 5253 7560 5256
rect 7594 5253 7606 5287
rect 7548 5247 7606 5253
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 11146 5284 11152 5296
rect 7892 5256 8050 5284
rect 8864 5256 11152 5284
rect 7892 5244 7898 5256
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 1670 5216 1676 5228
rect 1627 5188 1676 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2280 5188 2329 5216
rect 2280 5176 2286 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 2740 5188 3617 5216
rect 2740 5176 2746 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 5092 5188 6653 5216
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 5092 5148 5120 5188
rect 6641 5185 6653 5188
rect 6687 5216 6699 5219
rect 6822 5216 6828 5228
rect 6687 5188 6828 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7064 5188 7297 5216
rect 7064 5176 7070 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 4672 5120 5120 5148
rect 5629 5151 5687 5157
rect 4672 5108 4678 5120
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5718 5148 5724 5160
rect 5675 5120 5724 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 8864 5148 8892 5256
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 12802 5244 12808 5296
rect 12860 5284 12866 5296
rect 12860 5256 12905 5284
rect 12860 5244 12866 5256
rect 12986 5244 12992 5296
rect 13044 5284 13050 5296
rect 13648 5293 13676 5324
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 15102 5352 15108 5364
rect 15063 5324 15108 5352
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 17034 5352 17040 5364
rect 16255 5324 17040 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 18874 5352 18880 5364
rect 17512 5324 18880 5352
rect 13633 5287 13691 5293
rect 13633 5284 13645 5287
rect 13044 5256 13645 5284
rect 13044 5244 13050 5256
rect 13633 5253 13645 5256
rect 13679 5253 13691 5287
rect 13633 5247 13691 5253
rect 14090 5244 14096 5296
rect 14148 5244 14154 5296
rect 17512 5284 17540 5324
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19484 5324 19809 5352
rect 19484 5312 19490 5324
rect 19797 5321 19809 5324
rect 19843 5321 19855 5355
rect 19797 5315 19855 5321
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 20533 5355 20591 5361
rect 20533 5352 20545 5355
rect 20496 5324 20545 5352
rect 20496 5312 20502 5324
rect 20533 5321 20545 5324
rect 20579 5321 20591 5355
rect 20533 5315 20591 5321
rect 20714 5312 20720 5364
rect 20772 5352 20778 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 20772 5324 24041 5352
rect 20772 5312 20778 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24029 5315 24087 5321
rect 24118 5312 24124 5364
rect 24176 5352 24182 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24176 5324 24685 5352
rect 24176 5312 24182 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 21910 5284 21916 5296
rect 16684 5256 17540 5284
rect 18354 5256 21916 5284
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 10134 5216 10140 5228
rect 9723 5188 10140 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10318 5216 10324 5228
rect 10279 5188 10324 5216
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 10410 5176 10416 5228
rect 10468 5216 10474 5228
rect 10962 5216 10968 5228
rect 10468 5188 10968 5216
rect 10468 5176 10474 5188
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 12158 5216 12164 5228
rect 11572 5188 12164 5216
rect 11572 5176 11578 5188
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12721 5217 12779 5223
rect 12721 5183 12733 5217
rect 12767 5214 12779 5217
rect 12894 5216 12900 5228
rect 12820 5214 12900 5216
rect 12767 5188 12900 5214
rect 12767 5186 12848 5188
rect 12767 5183 12779 5186
rect 12721 5177 12779 5183
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 16114 5216 16120 5228
rect 15068 5188 16120 5216
rect 15068 5176 15074 5188
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 6932 5120 8892 5148
rect 2038 5040 2044 5092
rect 2096 5080 2102 5092
rect 6932 5080 6960 5120
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 12434 5148 12440 5160
rect 9548 5120 12440 5148
rect 9548 5108 9554 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12584 5120 13369 5148
rect 12584 5108 12590 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 16684 5148 16712 5256
rect 21910 5244 21916 5256
rect 21968 5244 21974 5296
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 24486 5284 24492 5296
rect 22244 5256 24492 5284
rect 22244 5244 22250 5256
rect 24486 5244 24492 5256
rect 24544 5244 24550 5296
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19702 5216 19708 5228
rect 19663 5188 19708 5216
rect 19245 5179 19303 5185
rect 16850 5148 16856 5160
rect 13357 5111 13415 5117
rect 13464 5120 16712 5148
rect 16811 5120 16856 5148
rect 10413 5083 10471 5089
rect 10413 5080 10425 5083
rect 2096 5052 3740 5080
rect 2096 5040 2102 5052
rect 14 4972 20 5024
rect 72 5012 78 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 72 4984 1777 5012
rect 72 4972 78 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 2774 5012 2780 5024
rect 2547 4984 2780 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 3712 5012 3740 5052
rect 4908 5052 6960 5080
rect 8588 5052 10425 5080
rect 4908 5012 4936 5052
rect 3712 4984 4936 5012
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 8588 5012 8616 5052
rect 10413 5049 10425 5052
rect 10459 5049 10471 5083
rect 13464 5080 13492 5120
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 16960 5120 17141 5148
rect 10413 5043 10471 5049
rect 12544 5052 13492 5080
rect 6420 4984 8616 5012
rect 6420 4972 6426 4984
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 12544 5012 12572 5052
rect 14826 5040 14832 5092
rect 14884 5080 14890 5092
rect 16960 5080 16988 5120
rect 17129 5117 17141 5120
rect 17175 5148 17187 5151
rect 18598 5148 18604 5160
rect 17175 5120 18604 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 19260 5148 19288 5179
rect 19702 5176 19708 5188
rect 19760 5176 19766 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20530 5216 20536 5228
rect 20487 5188 20536 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 21266 5216 21272 5228
rect 21227 5188 21272 5216
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22060 5188 22661 5216
rect 22060 5186 22103 5188
rect 22060 5176 22066 5186
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 23750 5216 23756 5228
rect 23339 5188 23756 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23750 5176 23756 5188
rect 23808 5216 23814 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23808 5188 23949 5216
rect 23808 5176 23814 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24581 5219 24639 5225
rect 24581 5185 24593 5219
rect 24627 5185 24639 5219
rect 26510 5216 26516 5228
rect 26471 5188 26516 5216
rect 24581 5179 24639 5185
rect 21818 5148 21824 5160
rect 19260 5120 21824 5148
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 21968 5120 23397 5148
rect 21968 5108 21974 5120
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 24596 5148 24624 5179
rect 26510 5176 26516 5188
rect 26568 5176 26574 5228
rect 38010 5216 38016 5228
rect 37971 5188 38016 5216
rect 38010 5176 38016 5188
rect 38068 5176 38074 5228
rect 23532 5120 24624 5148
rect 23532 5108 23538 5120
rect 23934 5080 23940 5092
rect 14884 5052 16988 5080
rect 18524 5052 23940 5080
rect 14884 5040 14890 5052
rect 10376 4984 12572 5012
rect 10376 4972 10382 4984
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 16482 5012 16488 5024
rect 12676 4984 16488 5012
rect 12676 4972 12682 4984
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 18524 5012 18552 5052
rect 23934 5040 23940 5052
rect 23992 5040 23998 5092
rect 16724 4984 18552 5012
rect 18601 5015 18659 5021
rect 16724 4972 16730 4984
rect 18601 4981 18613 5015
rect 18647 5012 18659 5015
rect 19242 5012 19248 5024
rect 18647 4984 19248 5012
rect 18647 4981 18659 4984
rect 18601 4975 18659 4981
rect 19242 4972 19248 4984
rect 19300 5012 19306 5024
rect 19702 5012 19708 5024
rect 19300 4984 19708 5012
rect 19300 4972 19306 4984
rect 19702 4972 19708 4984
rect 19760 4972 19766 5024
rect 21082 5012 21088 5024
rect 21043 4984 21088 5012
rect 21082 4972 21088 4984
rect 21140 4972 21146 5024
rect 21634 4972 21640 5024
rect 21692 5012 21698 5024
rect 21910 5012 21916 5024
rect 21692 4984 21916 5012
rect 21692 4972 21698 4984
rect 21910 4972 21916 4984
rect 21968 4972 21974 5024
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 22738 5012 22744 5024
rect 22152 4984 22197 5012
rect 22699 4984 22744 5012
rect 22152 4972 22158 4984
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 26329 5015 26387 5021
rect 26329 4981 26341 5015
rect 26375 5012 26387 5015
rect 32306 5012 32312 5024
rect 26375 4984 32312 5012
rect 26375 4981 26387 4984
rect 26329 4975 26387 4981
rect 32306 4972 32312 4984
rect 32364 4972 32370 5024
rect 37829 5015 37887 5021
rect 37829 4981 37841 5015
rect 37875 5012 37887 5015
rect 38010 5012 38016 5024
rect 37875 4984 38016 5012
rect 37875 4981 37887 4984
rect 37829 4975 37887 4981
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 6086 4808 6092 4820
rect 4755 4780 6092 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 8481 4811 8539 4817
rect 6196 4780 8432 4808
rect 3050 4740 3056 4752
rect 2884 4712 3056 4740
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2884 4672 2912 4712
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 6196 4740 6224 4780
rect 3200 4712 6224 4740
rect 7837 4743 7895 4749
rect 3200 4700 3206 4712
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 7926 4740 7932 4752
rect 7883 4712 7932 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 7926 4700 7932 4712
rect 7984 4700 7990 4752
rect 8404 4740 8432 4780
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 9306 4808 9312 4820
rect 8527 4780 9312 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 13262 4808 13268 4820
rect 9416 4780 10640 4808
rect 13223 4780 13268 4808
rect 9416 4740 9444 4780
rect 8404 4712 9444 4740
rect 10612 4740 10640 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 16022 4808 16028 4820
rect 15983 4780 16028 4808
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 18046 4808 18052 4820
rect 16448 4780 18052 4808
rect 16448 4768 16454 4780
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18506 4808 18512 4820
rect 18467 4780 18512 4808
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 18598 4768 18604 4820
rect 18656 4808 18662 4820
rect 21085 4811 21143 4817
rect 18656 4780 21036 4808
rect 18656 4768 18662 4780
rect 11422 4740 11428 4752
rect 10612 4712 11428 4740
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 17221 4743 17279 4749
rect 17221 4709 17233 4743
rect 17267 4740 17279 4743
rect 20622 4740 20628 4752
rect 17267 4712 20628 4740
rect 17267 4709 17279 4712
rect 17221 4703 17279 4709
rect 20622 4700 20628 4712
rect 20680 4700 20686 4752
rect 21008 4740 21036 4780
rect 21085 4777 21097 4811
rect 21131 4808 21143 4811
rect 21450 4808 21456 4820
rect 21131 4780 21456 4808
rect 21131 4777 21143 4780
rect 21085 4771 21143 4777
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 23382 4808 23388 4820
rect 21560 4780 23388 4808
rect 21560 4740 21588 4780
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 24762 4768 24768 4820
rect 24820 4808 24826 4820
rect 28261 4811 28319 4817
rect 28261 4808 28273 4811
rect 24820 4780 28273 4808
rect 24820 4768 24826 4780
rect 28261 4777 28273 4780
rect 28307 4777 28319 4811
rect 31938 4808 31944 4820
rect 31899 4780 31944 4808
rect 28261 4771 28319 4777
rect 31938 4768 31944 4780
rect 31996 4768 32002 4820
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 38105 4811 38163 4817
rect 38105 4808 38117 4811
rect 35860 4780 38117 4808
rect 35860 4768 35866 4780
rect 38105 4777 38117 4780
rect 38151 4777 38163 4811
rect 38105 4771 38163 4777
rect 23753 4743 23811 4749
rect 23753 4740 23765 4743
rect 21008 4712 21588 4740
rect 22066 4712 23765 4740
rect 1903 4644 2912 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3418 4672 3424 4684
rect 3292 4644 3424 4672
rect 3292 4632 3298 4644
rect 3418 4632 3424 4644
rect 3476 4672 3482 4684
rect 6089 4675 6147 4681
rect 3476 4644 4660 4672
rect 3476 4632 3482 4644
rect 4632 4616 4660 4644
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6454 4672 6460 4684
rect 6135 4644 6460 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6454 4632 6460 4644
rect 6512 4672 6518 4684
rect 7006 4672 7012 4684
rect 6512 4644 7012 4672
rect 6512 4632 6518 4644
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 9122 4672 9128 4684
rect 7852 4644 9128 4672
rect 7852 4616 7880 4644
rect 9122 4632 9128 4644
rect 9180 4672 9186 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 9180 4644 9321 4672
rect 9180 4632 9186 4644
rect 9309 4641 9321 4644
rect 9355 4672 9367 4675
rect 10134 4672 10140 4684
rect 9355 4644 10140 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 10134 4632 10140 4644
rect 10192 4672 10198 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 10192 4644 11529 4672
rect 10192 4632 10198 4644
rect 11517 4641 11529 4644
rect 11563 4672 11575 4675
rect 11790 4672 11796 4684
rect 11563 4644 11796 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 12216 4644 13308 4672
rect 12216 4632 12222 4644
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1544 4576 1593 4604
rect 1544 4564 1550 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 4157 4567 4215 4573
rect 3510 4536 3516 4548
rect 3082 4508 3516 4536
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 4172 4536 4200 4567
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5442 4604 5448 4616
rect 5215 4576 5448 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 11330 4564 11336 4616
rect 11388 4564 11394 4616
rect 13280 4604 13308 4644
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14274 4672 14280 4684
rect 14056 4644 14280 4672
rect 14056 4632 14062 4644
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 14550 4672 14556 4684
rect 14511 4644 14556 4672
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 16666 4672 16672 4684
rect 16627 4644 16672 4672
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 22066 4672 22094 4712
rect 23753 4709 23765 4712
rect 23799 4709 23811 4743
rect 23753 4703 23811 4709
rect 23842 4700 23848 4752
rect 23900 4740 23906 4752
rect 27614 4740 27620 4752
rect 23900 4712 27620 4740
rect 23900 4700 23906 4712
rect 27614 4700 27620 4712
rect 27672 4700 27678 4752
rect 18095 4644 22094 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 14182 4604 14188 4616
rect 13280 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 18874 4564 18880 4616
rect 18932 4604 18938 4616
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 18932 4576 19993 4604
rect 18932 4564 18938 4576
rect 19981 4573 19993 4576
rect 20027 4604 20039 4607
rect 20162 4604 20168 4616
rect 20027 4576 20168 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 21266 4604 21272 4616
rect 21227 4576 21272 4604
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22002 4604 22008 4616
rect 21867 4576 22008 4604
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 22002 4564 22008 4576
rect 22060 4604 22066 4616
rect 22465 4607 22523 4613
rect 22465 4604 22477 4607
rect 22060 4576 22477 4604
rect 22060 4564 22066 4576
rect 22465 4573 22477 4576
rect 22511 4604 22523 4607
rect 23109 4607 23167 4613
rect 23109 4604 23121 4607
rect 22511 4576 23121 4604
rect 22511 4573 22523 4576
rect 22465 4567 22523 4573
rect 23109 4573 23121 4576
rect 23155 4573 23167 4607
rect 23934 4604 23940 4616
rect 23895 4576 23940 4604
rect 23109 4567 23167 4573
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 28169 4607 28227 4613
rect 28169 4573 28181 4607
rect 28215 4604 28227 4607
rect 31849 4607 31907 4613
rect 28215 4576 31754 4604
rect 28215 4573 28227 4576
rect 28169 4567 28227 4573
rect 4172 4508 6316 4536
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 4614 4468 4620 4480
rect 4295 4440 4620 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5626 4468 5632 4480
rect 5587 4440 5632 4468
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 6288 4468 6316 4508
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 6420 4508 6465 4536
rect 6420 4496 6426 4508
rect 6914 4496 6920 4548
rect 6972 4496 6978 4548
rect 7760 4508 9536 4536
rect 7760 4468 7788 4508
rect 6288 4440 7788 4468
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 8662 4468 8668 4480
rect 8260 4440 8668 4468
rect 8260 4428 8266 4440
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 9508 4468 9536 4508
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 10870 4536 10876 4548
rect 9640 4508 9685 4536
rect 10810 4508 10876 4536
rect 9640 4496 9646 4508
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 11348 4536 11376 4564
rect 11072 4508 11376 4536
rect 10318 4468 10324 4480
rect 9508 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 11072 4477 11100 4508
rect 11514 4496 11520 4548
rect 11572 4536 11578 4548
rect 11793 4539 11851 4545
rect 11793 4536 11805 4539
rect 11572 4508 11805 4536
rect 11572 4496 11578 4508
rect 11793 4505 11805 4508
rect 11839 4505 11851 4539
rect 11793 4499 11851 4505
rect 12250 4496 12256 4548
rect 12308 4496 12314 4548
rect 13832 4508 14964 4536
rect 15778 4508 16712 4536
rect 11057 4471 11115 4477
rect 11057 4437 11069 4471
rect 11103 4437 11115 4471
rect 11057 4431 11115 4437
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 13832 4468 13860 4508
rect 11388 4440 13860 4468
rect 11388 4428 11394 4440
rect 13906 4428 13912 4480
rect 13964 4468 13970 4480
rect 14826 4468 14832 4480
rect 13964 4440 14832 4468
rect 13964 4428 13970 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 14936 4468 14964 4508
rect 15470 4468 15476 4480
rect 14936 4440 15476 4468
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 16684 4468 16712 4508
rect 16758 4496 16764 4548
rect 16816 4536 16822 4548
rect 16816 4508 16861 4536
rect 16816 4496 16822 4508
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 23201 4539 23259 4545
rect 23201 4536 23213 4539
rect 18012 4508 23213 4536
rect 18012 4496 18018 4508
rect 23201 4505 23213 4508
rect 23247 4505 23259 4539
rect 31726 4536 31754 4576
rect 31849 4573 31861 4607
rect 31895 4604 31907 4607
rect 33870 4604 33876 4616
rect 31895 4576 33876 4604
rect 31895 4573 31907 4576
rect 31849 4567 31907 4573
rect 33870 4564 33876 4576
rect 33928 4564 33934 4616
rect 38286 4604 38292 4616
rect 38247 4576 38292 4604
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 33594 4536 33600 4548
rect 31726 4508 33600 4536
rect 23201 4499 23259 4505
rect 33594 4496 33600 4508
rect 33652 4496 33658 4548
rect 19150 4468 19156 4480
rect 16684 4440 19156 4468
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 20070 4468 20076 4480
rect 20031 4440 20076 4468
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 21910 4468 21916 4480
rect 21871 4440 21916 4468
rect 21910 4428 21916 4440
rect 21968 4428 21974 4480
rect 22554 4468 22560 4480
rect 22515 4440 22560 4468
rect 22554 4428 22560 4440
rect 22612 4428 22618 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2464 4236 2774 4264
rect 2464 4224 2470 4236
rect 1578 4196 1584 4208
rect 1539 4168 1584 4196
rect 1578 4156 1584 4168
rect 1636 4156 1642 4208
rect 2746 4196 2774 4236
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 7650 4264 7656 4276
rect 4120 4236 7656 4264
rect 4120 4224 4126 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 8404 4236 9536 4264
rect 2746 4168 4554 4196
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 6362 4196 6368 4208
rect 6052 4168 6368 4196
rect 6052 4156 6058 4168
rect 6362 4156 6368 4168
rect 6420 4196 6426 4208
rect 8404 4196 8432 4236
rect 6420 4168 8432 4196
rect 6420 4156 6426 4168
rect 8662 4156 8668 4208
rect 8720 4156 8726 4208
rect 9508 4196 9536 4236
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 12158 4264 12164 4276
rect 9640 4236 12164 4264
rect 9640 4224 9646 4236
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12250 4224 12256 4276
rect 12308 4264 12314 4276
rect 14090 4264 14096 4276
rect 12308 4236 14096 4264
rect 12308 4224 12314 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 22738 4264 22744 4276
rect 14660 4236 22744 4264
rect 11330 4196 11336 4208
rect 9508 4168 11336 4196
rect 11330 4156 11336 4168
rect 11388 4156 11394 4208
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 12342 4196 12348 4208
rect 11572 4168 12348 4196
rect 11572 4156 11578 4168
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 14660 4196 14688 4236
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 23845 4267 23903 4273
rect 23845 4233 23857 4267
rect 23891 4264 23903 4267
rect 23934 4264 23940 4276
rect 23891 4236 23940 4264
rect 23891 4233 23903 4236
rect 23845 4227 23903 4233
rect 23934 4224 23940 4236
rect 23992 4224 23998 4276
rect 24486 4224 24492 4276
rect 24544 4264 24550 4276
rect 24581 4267 24639 4273
rect 24581 4264 24593 4267
rect 24544 4236 24593 4264
rect 24544 4224 24550 4236
rect 24581 4233 24593 4236
rect 24627 4233 24639 4267
rect 24581 4227 24639 4233
rect 22554 4196 22560 4208
rect 13294 4168 14688 4196
rect 15502 4168 22560 4196
rect 22554 4156 22560 4168
rect 22612 4156 22618 4208
rect 23382 4156 23388 4208
rect 23440 4196 23446 4208
rect 23440 4168 23520 4196
rect 23440 4156 23446 4168
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 2740 4100 3801 4128
rect 2740 4088 2746 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 7190 4128 7196 4140
rect 5859 4100 7196 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7892 4100 7941 4128
rect 7892 4088 7898 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 10318 4128 10324 4140
rect 10279 4100 10324 4128
rect 7929 4091 7987 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11238 4128 11244 4140
rect 11103 4100 11244 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13280 4100 14013 4128
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 3752 4032 4077 4060
rect 3752 4020 3758 4032
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 5960 4032 6561 4060
rect 5960 4020 5966 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 6825 4023 6883 4029
rect 8036 4032 8217 4060
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 6086 3924 6092 3936
rect 1912 3896 6092 3924
rect 1912 3884 1918 3896
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6840 3924 6868 4023
rect 7926 3952 7932 4004
rect 7984 3992 7990 4004
rect 8036 3992 8064 4032
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 11698 4060 11704 4072
rect 9640 4032 11704 4060
rect 9640 4020 9646 4032
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 9950 3992 9956 4004
rect 7984 3964 8064 3992
rect 9600 3964 9956 3992
rect 7984 3952 7990 3964
rect 9600 3924 9628 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 6840 3896 9628 3924
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9766 3924 9772 3936
rect 9723 3896 9772 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11808 3924 11836 4088
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 13280 3924 13308 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 14001 4091 14059 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17276 4100 17969 4128
rect 17276 4088 17282 4100
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18104 4100 19165 4128
rect 18104 4088 18110 4100
rect 19153 4097 19165 4100
rect 19199 4128 19211 4131
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19199 4100 19625 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 19978 4128 19984 4140
rect 19751 4100 19984 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 20128 4100 20269 4128
rect 20128 4088 20134 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20404 4100 20449 4128
rect 20404 4088 20410 4100
rect 20990 4088 20996 4140
rect 21048 4128 21054 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21048 4100 21281 4128
rect 21048 4088 21054 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23014 4128 23020 4140
rect 22327 4100 23020 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 23492 4128 23520 4168
rect 23750 4156 23756 4208
rect 23808 4196 23814 4208
rect 23808 4168 24624 4196
rect 23808 4156 23814 4168
rect 24029 4131 24087 4137
rect 24029 4128 24041 4131
rect 23348 4100 23393 4128
rect 23492 4100 24041 4128
rect 23348 4088 23354 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 24029 4091 24087 4097
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4097 24547 4131
rect 24596 4128 24624 4168
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 24596 4100 25145 4128
rect 24489 4091 24547 4097
rect 25133 4097 25145 4100
rect 25179 4097 25191 4131
rect 25133 4091 25191 4097
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 13630 4060 13636 4072
rect 13587 4032 13636 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 13630 4020 13636 4032
rect 13688 4060 13694 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13688 4032 14289 4060
rect 13688 4020 13694 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 20530 4060 20536 4072
rect 14277 4023 14335 4029
rect 15304 4032 20536 4060
rect 11572 3896 13308 3924
rect 11572 3884 11578 3896
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 15304 3924 15332 4032
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 20772 4032 22569 4060
rect 20772 4020 20778 4032
rect 22557 4029 22569 4032
rect 22603 4060 22615 4063
rect 23750 4060 23756 4072
rect 22603 4032 23756 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 15378 3952 15384 4004
rect 15436 3992 15442 4004
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 15436 3964 15761 3992
rect 15436 3952 15442 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 15749 3955 15807 3961
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 15988 3964 17233 3992
rect 15988 3952 15994 3964
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17221 3955 17279 3961
rect 17773 3995 17831 4001
rect 17773 3961 17785 3995
rect 17819 3992 17831 3995
rect 18782 3992 18788 4004
rect 17819 3964 18788 3992
rect 17819 3961 17831 3964
rect 17773 3955 17831 3961
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 18969 3995 19027 4001
rect 18969 3961 18981 3995
rect 19015 3992 19027 3995
rect 21266 3992 21272 4004
rect 19015 3964 21272 3992
rect 19015 3961 19027 3964
rect 18969 3955 19027 3961
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 24504 3992 24532 4091
rect 37182 4088 37188 4140
rect 37240 4128 37246 4140
rect 38289 4131 38347 4137
rect 38289 4128 38301 4131
rect 37240 4100 38301 4128
rect 37240 4088 37246 4100
rect 38289 4097 38301 4100
rect 38335 4097 38347 4131
rect 38289 4091 38347 4097
rect 21600 3964 24532 3992
rect 21600 3952 21606 3964
rect 36354 3952 36360 4004
rect 36412 3992 36418 4004
rect 38105 3995 38163 4001
rect 38105 3992 38117 3995
rect 36412 3964 38117 3992
rect 36412 3952 36418 3964
rect 38105 3961 38117 3964
rect 38151 3961 38163 3995
rect 38105 3955 38163 3961
rect 14148 3896 15332 3924
rect 14148 3884 14154 3896
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 21082 3924 21088 3936
rect 15528 3896 21088 3924
rect 15528 3884 15534 3896
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 21361 3927 21419 3933
rect 21361 3924 21373 3927
rect 21232 3896 21373 3924
rect 21232 3884 21238 3896
rect 21361 3893 21373 3896
rect 21407 3893 21419 3927
rect 25222 3924 25228 3936
rect 25183 3896 25228 3924
rect 21361 3887 21419 3893
rect 25222 3884 25228 3896
rect 25280 3884 25286 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 5350 3720 5356 3732
rect 3375 3692 5356 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 7926 3720 7932 3732
rect 5776 3692 7932 3720
rect 5776 3680 5782 3692
rect 7926 3680 7932 3692
rect 7984 3720 7990 3732
rect 9582 3720 9588 3732
rect 7984 3692 9588 3720
rect 7984 3680 7990 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 16574 3720 16580 3732
rect 13320 3692 16580 3720
rect 13320 3680 13326 3692
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 16684 3692 19625 3720
rect 11974 3612 11980 3664
rect 12032 3652 12038 3664
rect 14090 3652 14096 3664
rect 12032 3624 14096 3652
rect 12032 3612 12038 3624
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15988 3624 16037 3652
rect 15988 3612 15994 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 16025 3615 16083 3621
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 16684 3652 16712 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 19613 3683 19671 3689
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 23474 3720 23480 3732
rect 20404 3692 23480 3720
rect 20404 3680 20410 3692
rect 22278 3652 22284 3664
rect 16540 3624 16712 3652
rect 17880 3624 22284 3652
rect 16540 3612 16546 3624
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3384 3556 3985 3584
rect 3384 3544 3390 3556
rect 3973 3553 3985 3556
rect 4019 3584 4031 3587
rect 6454 3584 6460 3596
rect 4019 3556 6460 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 8478 3584 8484 3596
rect 6779 3556 8484 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10192 3556 10425 3584
rect 10192 3544 10198 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 12250 3584 12256 3596
rect 10735 3556 12256 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 12400 3556 12449 3584
rect 12400 3544 12406 3556
rect 12437 3553 12449 3556
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 14056 3556 14289 3584
rect 14056 3544 14062 3556
rect 14277 3553 14289 3556
rect 14323 3584 14335 3587
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 14323 3556 16589 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 16577 3553 16589 3556
rect 16623 3584 16635 3587
rect 16850 3584 16856 3596
rect 16623 3556 16856 3584
rect 16623 3553 16635 3556
rect 16577 3547 16635 3553
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17880 3584 17908 3624
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 21542 3584 21548 3596
rect 17276 3556 17908 3584
rect 21503 3556 21548 3584
rect 17276 3544 17282 3556
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 22480 3593 22508 3692
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 33870 3680 33876 3732
rect 33928 3720 33934 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 33928 3692 38117 3720
rect 33928 3680 33934 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 23198 3612 23204 3664
rect 23256 3652 23262 3664
rect 23256 3624 23428 3652
rect 23256 3612 23262 3624
rect 23400 3593 23428 3624
rect 23566 3612 23572 3664
rect 23624 3652 23630 3664
rect 25225 3655 25283 3661
rect 25225 3652 25237 3655
rect 23624 3624 25237 3652
rect 23624 3612 23630 3624
rect 25225 3621 25237 3624
rect 25271 3621 25283 3655
rect 25225 3615 25283 3621
rect 22465 3587 22523 3593
rect 22465 3553 22477 3587
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 23385 3587 23443 3593
rect 23385 3553 23397 3587
rect 23431 3553 23443 3587
rect 23385 3547 23443 3553
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9674 3516 9680 3528
rect 9355 3488 9680 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9824 3488 9869 3516
rect 9824 3476 9830 3488
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 12768 3488 13461 3516
rect 12768 3476 12774 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 19518 3516 19524 3528
rect 19479 3488 19524 3516
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 20162 3476 20168 3488
rect 20220 3516 20226 3528
rect 20714 3516 20720 3528
rect 20220 3488 20720 3516
rect 20220 3476 20226 3488
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21048 3488 21281 3516
rect 21048 3476 21054 3488
rect 21269 3485 21281 3488
rect 21315 3516 21327 3519
rect 22002 3516 22008 3528
rect 21315 3488 22008 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 22281 3519 22339 3525
rect 22281 3485 22293 3519
rect 22327 3516 22339 3519
rect 23014 3516 23020 3528
rect 22327 3488 23020 3516
rect 22327 3485 22339 3488
rect 22281 3479 22339 3485
rect 23014 3476 23020 3488
rect 23072 3516 23078 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 23072 3488 23213 3516
rect 23072 3476 23078 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 23201 3479 23259 3485
rect 3082 3420 3648 3448
rect 3620 3380 3648 3420
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 4304 3420 4349 3448
rect 4304 3408 4310 3420
rect 4706 3408 4712 3460
rect 4764 3408 4770 3460
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3448 6055 3451
rect 6638 3448 6644 3460
rect 6043 3420 6644 3448
rect 6043 3417 6055 3420
rect 5997 3411 6055 3417
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 7374 3408 7380 3460
rect 7432 3408 7438 3460
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 8481 3451 8539 3457
rect 8481 3448 8493 3451
rect 8076 3420 8493 3448
rect 8076 3408 8082 3420
rect 8481 3417 8493 3420
rect 8527 3417 8539 3451
rect 10410 3448 10416 3460
rect 8481 3411 8539 3417
rect 8956 3420 10416 3448
rect 4614 3380 4620 3392
rect 3620 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 8956 3380 8984 3420
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 11146 3408 11152 3460
rect 11204 3408 11210 3460
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 13262 3448 13268 3460
rect 12032 3420 13268 3448
rect 12032 3408 12038 3420
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 14274 3448 14280 3460
rect 13556 3420 14280 3448
rect 9122 3380 9128 3392
rect 5868 3352 8984 3380
rect 9083 3352 9128 3380
rect 5868 3340 5874 3352
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 13556 3380 13584 3420
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 16482 3448 16488 3460
rect 14599 3420 14964 3448
rect 15778 3420 16488 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 9907 3352 13584 3380
rect 13633 3383 13691 3389
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 14826 3380 14832 3392
rect 13679 3352 14832 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 14936 3380 14964 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 16758 3408 16764 3460
rect 16816 3448 16822 3460
rect 16853 3451 16911 3457
rect 16853 3448 16865 3451
rect 16816 3420 16865 3448
rect 16816 3408 16822 3420
rect 16853 3417 16865 3420
rect 16899 3448 16911 3451
rect 16942 3448 16948 3460
rect 16899 3420 16948 3448
rect 16899 3417 16911 3420
rect 16853 3411 16911 3417
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 18196 3420 20392 3448
rect 18196 3408 18202 3420
rect 15930 3380 15936 3392
rect 14936 3352 15936 3380
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 17034 3380 17040 3392
rect 16264 3352 17040 3380
rect 16264 3340 16270 3352
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 18325 3383 18383 3389
rect 18325 3380 18337 3383
rect 17184 3352 18337 3380
rect 17184 3340 17190 3352
rect 18325 3349 18337 3352
rect 18371 3349 18383 3383
rect 18325 3343 18383 3349
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 20070 3380 20076 3392
rect 18564 3352 20076 3380
rect 18564 3340 18570 3352
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 20364 3380 20392 3420
rect 20438 3408 20444 3460
rect 20496 3448 20502 3460
rect 22094 3448 22100 3460
rect 20496 3420 22100 3448
rect 20496 3408 20502 3420
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 23216 3448 23244 3479
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3516 24731 3519
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 24719 3488 25421 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 27672 3488 36093 3516
rect 27672 3476 27678 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 38289 3519 38347 3525
rect 38289 3516 38301 3519
rect 38160 3488 38301 3516
rect 38160 3476 38166 3488
rect 38289 3485 38301 3488
rect 38335 3485 38347 3519
rect 38289 3479 38347 3485
rect 37918 3448 37924 3460
rect 23216 3420 37924 3448
rect 37918 3408 37924 3420
rect 37976 3408 37982 3460
rect 24762 3380 24768 3392
rect 20364 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 36173 3383 36231 3389
rect 36173 3349 36185 3383
rect 36219 3380 36231 3383
rect 36906 3380 36912 3392
rect 36219 3352 36912 3380
rect 36219 3349 36231 3352
rect 36173 3343 36231 3349
rect 36906 3340 36912 3352
rect 36964 3340 36970 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3970 3176 3976 3188
rect 3384 3148 3976 3176
rect 3384 3136 3390 3148
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 11974 3176 11980 3188
rect 6871 3148 11980 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 15654 3136 15660 3188
rect 15712 3136 15718 3188
rect 15749 3179 15807 3185
rect 15749 3145 15761 3179
rect 15795 3176 15807 3179
rect 16758 3176 16764 3188
rect 15795 3148 16764 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 20438 3176 20444 3188
rect 16960 3148 20444 3176
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 1636 3080 3556 3108
rect 1636 3068 1642 3080
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3234 3040 3240 3052
rect 2915 3012 3240 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3528 3049 3556 3080
rect 4798 3068 4804 3120
rect 4856 3068 4862 3120
rect 5166 3068 5172 3120
rect 5224 3108 5230 3120
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 5224 3080 5549 3108
rect 5224 3068 5230 3080
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 5537 3071 5595 3077
rect 7193 3111 7251 3117
rect 7193 3077 7205 3111
rect 7239 3108 7251 3111
rect 7466 3108 7472 3120
rect 7239 3080 7472 3108
rect 7239 3077 7251 3080
rect 7193 3071 7251 3077
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 7208 3040 7236 3071
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 9214 3108 9220 3120
rect 8786 3080 9220 3108
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 9456 3080 11805 3108
rect 9456 3068 9462 3080
rect 11793 3077 11805 3080
rect 11839 3108 11851 3111
rect 11882 3108 11888 3120
rect 11839 3080 11888 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 15672 3108 15700 3136
rect 16960 3108 16988 3148
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 20588 3148 21404 3176
rect 20588 3136 20594 3148
rect 17126 3108 17132 3120
rect 15672 3080 16988 3108
rect 17087 3080 17132 3108
rect 17126 3068 17132 3080
rect 17184 3068 17190 3120
rect 21174 3108 21180 3120
rect 18354 3080 21180 3108
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 21269 3111 21327 3117
rect 21269 3077 21281 3111
rect 21315 3108 21327 3111
rect 21376 3108 21404 3148
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 23109 3179 23167 3185
rect 23109 3176 23121 3179
rect 22060 3148 23121 3176
rect 22060 3136 22066 3148
rect 23109 3145 23121 3148
rect 23155 3145 23167 3179
rect 25774 3176 25780 3188
rect 25735 3148 25780 3176
rect 23109 3139 23167 3145
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 22094 3108 22100 3120
rect 21315 3080 21404 3108
rect 21468 3080 22100 3108
rect 21315 3077 21327 3080
rect 21269 3071 21327 3077
rect 6687 3012 7236 3040
rect 9309 3043 9367 3049
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9490 3040 9496 3052
rect 9355 3012 9496 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 13170 3040 13176 3052
rect 10919 3012 13176 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1360 2944 1593 2972
rect 1360 2932 1366 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 3326 2972 3332 2984
rect 1903 2944 3332 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3476 2944 3801 2972
rect 3476 2932 3482 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 6730 2972 6736 2984
rect 6512 2944 6736 2972
rect 6512 2932 6518 2944
rect 6730 2932 6736 2944
rect 6788 2972 6794 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6788 2944 7297 2972
rect 6788 2932 6794 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 9030 2972 9036 2984
rect 7607 2944 9036 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9784 2972 9812 3003
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13998 3040 14004 3052
rect 13495 3012 14004 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 15378 3000 15384 3052
rect 15436 3000 15442 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3040 19395 3043
rect 19426 3040 19432 3052
rect 19383 3012 19432 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 20162 3040 20168 3052
rect 20027 3012 20168 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 20990 3040 20996 3052
rect 20951 3012 20996 3040
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21468 3040 21496 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 22204 3080 24716 3108
rect 22002 3040 22008 3052
rect 21100 3012 21496 3040
rect 21963 3012 22008 3040
rect 13814 2972 13820 2984
rect 9784 2944 13820 2972
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 16022 2972 16028 2984
rect 14323 2944 16028 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 21100 2972 21128 3012
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 22204 3040 22232 3080
rect 22112 3012 22232 3040
rect 19352 2944 21128 2972
rect 19352 2916 19380 2944
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 22112 2972 22140 3012
rect 22278 3000 22284 3052
rect 22336 3040 22342 3052
rect 23014 3040 23020 3052
rect 22336 3012 22381 3040
rect 22975 3012 23020 3040
rect 22336 3000 22342 3012
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23382 3000 23388 3052
rect 23440 3040 23446 3052
rect 24688 3049 24716 3080
rect 24762 3068 24768 3120
rect 24820 3108 24826 3120
rect 24820 3080 26004 3108
rect 24820 3068 24826 3080
rect 25976 3049 26004 3080
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23440 3012 23857 3040
rect 23440 3000 23446 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 24673 3043 24731 3049
rect 24673 3009 24685 3043
rect 24719 3009 24731 3043
rect 24673 3003 24731 3009
rect 25133 3043 25191 3049
rect 25133 3009 25145 3043
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25961 3043 26019 3049
rect 25961 3009 25973 3043
rect 26007 3009 26019 3043
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 25961 3003 26019 3009
rect 21324 2944 22140 2972
rect 21324 2932 21330 2944
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 22830 2972 22836 2984
rect 22244 2944 22836 2972
rect 22244 2932 22250 2944
rect 22830 2932 22836 2944
rect 22888 2932 22894 2984
rect 23937 2975 23995 2981
rect 23937 2972 23949 2975
rect 22940 2944 23949 2972
rect 9582 2904 9588 2916
rect 4816 2876 7328 2904
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 4816 2836 4844 2876
rect 3007 2808 4844 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5258 2836 5264 2848
rect 4948 2808 5264 2836
rect 4948 2796 4954 2808
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 7300 2836 7328 2876
rect 8588 2876 9588 2904
rect 8588 2836 8616 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 13630 2904 13636 2916
rect 9732 2876 13636 2904
rect 9732 2864 9738 2876
rect 13630 2864 13636 2876
rect 13688 2864 13694 2916
rect 15304 2876 15884 2904
rect 7300 2808 8616 2836
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9953 2839 10011 2845
rect 9953 2836 9965 2839
rect 9088 2808 9965 2836
rect 9088 2796 9094 2808
rect 9953 2805 9965 2808
rect 9999 2805 10011 2839
rect 9953 2799 10011 2805
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2836 11115 2839
rect 11606 2836 11612 2848
rect 11103 2808 11612 2836
rect 11103 2805 11115 2808
rect 11057 2799 11115 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 15304 2836 15332 2876
rect 12492 2808 15332 2836
rect 15856 2836 15884 2876
rect 19334 2864 19340 2916
rect 19392 2864 19398 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19484 2876 19529 2904
rect 19484 2864 19490 2876
rect 19610 2864 19616 2916
rect 19668 2904 19674 2916
rect 22940 2904 22968 2944
rect 23937 2941 23949 2944
rect 23983 2941 23995 2975
rect 25148 2972 25176 3003
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 38010 3040 38016 3052
rect 37971 3012 38016 3040
rect 38010 3000 38016 3012
rect 38068 3000 38074 3052
rect 27522 2972 27528 2984
rect 25148 2944 27528 2972
rect 23937 2935 23995 2941
rect 27522 2932 27528 2944
rect 27580 2932 27586 2984
rect 24489 2907 24547 2913
rect 24489 2904 24501 2907
rect 19668 2876 22968 2904
rect 23032 2876 24501 2904
rect 19668 2864 19674 2876
rect 18601 2839 18659 2845
rect 18601 2836 18613 2839
rect 15856 2808 18613 2836
rect 12492 2796 12498 2808
rect 18601 2805 18613 2808
rect 18647 2805 18659 2839
rect 18601 2799 18659 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19208 2808 20085 2836
rect 19208 2796 19214 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 23032 2836 23060 2876
rect 24489 2873 24501 2876
rect 24535 2873 24547 2907
rect 24489 2867 24547 2873
rect 20220 2808 23060 2836
rect 20220 2796 20226 2808
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 23164 2808 25237 2836
rect 23164 2796 23170 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 36725 2839 36783 2845
rect 36725 2805 36737 2839
rect 36771 2836 36783 2839
rect 38010 2836 38016 2848
rect 36771 2808 38016 2836
rect 36771 2805 36783 2808
rect 36725 2799 36783 2805
rect 38010 2796 38016 2808
rect 38068 2796 38074 2848
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 13446 2632 13452 2644
rect 5684 2604 13452 2632
rect 5684 2592 5690 2604
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 13998 2632 14004 2644
rect 13587 2604 14004 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16022 2632 16028 2644
rect 15983 2604 16028 2632
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 18233 2635 18291 2641
rect 18233 2601 18245 2635
rect 18279 2632 18291 2635
rect 18598 2632 18604 2644
rect 18279 2604 18604 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 18690 2592 18696 2644
rect 18748 2632 18754 2644
rect 18748 2604 18793 2632
rect 18748 2592 18754 2604
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 19116 2604 20269 2632
rect 19116 2592 19122 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 23716 2604 27169 2632
rect 23716 2592 23722 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 27157 2595 27215 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 30377 2635 30435 2641
rect 30377 2632 30389 2635
rect 29840 2604 30389 2632
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 8478 2564 8484 2576
rect 3375 2536 4108 2564
rect 8439 2536 8484 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2496 1642 2508
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 1636 2468 3985 2496
rect 1636 2456 1642 2468
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 4080 2496 4108 2536
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 19334 2564 19340 2576
rect 9180 2536 11928 2564
rect 9180 2524 9186 2536
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4080 2468 4261 2496
rect 3973 2459 4031 2465
rect 4249 2465 4261 2468
rect 4295 2496 4307 2499
rect 5994 2496 6000 2508
rect 4295 2468 5672 2496
rect 5955 2468 6000 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 3082 2332 4200 2360
rect 4172 2292 4200 2332
rect 4706 2320 4712 2372
rect 4764 2320 4770 2372
rect 5534 2292 5540 2304
rect 4172 2264 5540 2292
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 5644 2292 5672 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 10042 2496 10048 2508
rect 7055 2468 10048 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 11514 2496 11520 2508
rect 11195 2468 11520 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11514 2456 11520 2468
rect 11572 2496 11578 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11572 2468 11805 2496
rect 11572 2456 11578 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11900 2496 11928 2536
rect 13280 2536 14412 2564
rect 13280 2496 13308 2536
rect 11900 2468 13308 2496
rect 11793 2459 11851 2465
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 14148 2468 14289 2496
rect 14148 2456 14154 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14384 2496 14412 2536
rect 17604 2536 19340 2564
rect 14384 2468 17264 2496
rect 14277 2459 14335 2465
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16632 2400 16865 2428
rect 16632 2388 16638 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 8294 2360 8300 2372
rect 8234 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 8570 2360 8576 2372
rect 8404 2332 8576 2360
rect 8404 2292 8432 2332
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 12066 2360 12072 2372
rect 12027 2332 12072 2360
rect 12066 2320 12072 2332
rect 12124 2320 12130 2372
rect 14090 2360 14096 2372
rect 13294 2332 14096 2360
rect 14090 2320 14096 2332
rect 14148 2320 14154 2372
rect 14182 2320 14188 2372
rect 14240 2360 14246 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14240 2332 14565 2360
rect 14240 2320 14246 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 15562 2320 15568 2372
rect 15620 2320 15626 2372
rect 17236 2360 17264 2468
rect 17604 2437 17632 2536
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 27522 2524 27528 2576
rect 27580 2564 27586 2576
rect 29840 2564 29868 2604
rect 30377 2601 30389 2604
rect 30423 2601 30435 2635
rect 33594 2632 33600 2644
rect 33555 2604 33600 2632
rect 30377 2595 30435 2601
rect 33594 2592 33600 2604
rect 33652 2592 33658 2644
rect 27580 2536 29868 2564
rect 27580 2524 27586 2536
rect 30282 2524 30288 2576
rect 30340 2564 30346 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 30340 2536 34897 2564
rect 30340 2524 30346 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 17696 2468 18000 2496
rect 17589 2431 17647 2437
rect 17589 2397 17601 2431
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 17696 2360 17724 2468
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17972 2428 18000 2468
rect 18800 2468 24624 2496
rect 18800 2428 18828 2468
rect 17972 2400 18828 2428
rect 17773 2391 17831 2397
rect 17236 2332 17724 2360
rect 5644 2264 8432 2292
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17788 2292 17816 2391
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19429 2431 19487 2437
rect 18932 2400 18977 2428
rect 18932 2388 18938 2400
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2428 20223 2431
rect 20254 2428 20260 2440
rect 20211 2400 20260 2428
rect 20211 2397 20223 2400
rect 20165 2391 20223 2397
rect 17954 2320 17960 2372
rect 18012 2360 18018 2372
rect 19444 2360 19472 2391
rect 20254 2388 20260 2400
rect 20312 2428 20318 2440
rect 20809 2431 20867 2437
rect 20809 2428 20821 2431
rect 20312 2400 20821 2428
rect 20312 2388 20318 2400
rect 20809 2397 20821 2400
rect 20855 2397 20867 2431
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 20809 2391 20867 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23566 2428 23572 2440
rect 22971 2400 23572 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 23661 2431 23719 2437
rect 23661 2397 23673 2431
rect 23707 2428 23719 2431
rect 23750 2428 23756 2440
rect 23707 2400 23756 2428
rect 23707 2397 23719 2400
rect 23661 2391 23719 2397
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 24596 2437 24624 2468
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 33100 2468 35894 2496
rect 33100 2456 33106 2468
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24670 2388 24676 2440
rect 24728 2428 24734 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24728 2400 25881 2428
rect 24728 2388 24734 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30340 2400 30573 2428
rect 30340 2388 30346 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 30561 2391 30619 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 33560 2400 33793 2428
rect 33560 2388 33566 2400
rect 33781 2397 33793 2400
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34848 2400 35081 2428
rect 34848 2388 34854 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35866 2428 35894 2468
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35866 2400 36185 2428
rect 35069 2391 35127 2397
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 38010 2428 38016 2440
rect 37971 2400 38016 2428
rect 36173 2391 36231 2397
rect 38010 2388 38016 2400
rect 38068 2388 38074 2440
rect 22278 2360 22284 2372
rect 18012 2332 19472 2360
rect 22239 2332 22284 2360
rect 18012 2320 18018 2332
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 17862 2292 17868 2304
rect 17788 2264 17868 2292
rect 17037 2255 17095 2261
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 19613 2255 19671 2261
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22612 2264 23121 2292
rect 22612 2252 22618 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 23753 2295 23811 2301
rect 23753 2292 23765 2295
rect 23532 2264 23765 2292
rect 23532 2252 23538 2264
rect 23753 2261 23765 2264
rect 23799 2261 23811 2295
rect 23753 2255 23811 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 23900 2264 24777 2292
rect 23900 2252 23906 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 31628 2264 32505 2292
rect 31628 2252 31634 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 38197 2295 38255 2301
rect 38197 2261 38209 2295
rect 38243 2292 38255 2295
rect 39298 2292 39304 2304
rect 38243 2264 39304 2292
rect 38243 2261 38255 2264
rect 38197 2255 38255 2261
rect 39298 2252 39304 2264
rect 39356 2252 39362 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 5224 2060 17356 2088
rect 5224 2048 5230 2060
rect 1854 1980 1860 2032
rect 1912 2020 1918 2032
rect 7926 2020 7932 2032
rect 1912 1992 7932 2020
rect 1912 1980 1918 1992
rect 7926 1980 7932 1992
rect 7984 1980 7990 2032
rect 8478 1980 8484 2032
rect 8536 2020 8542 2032
rect 8536 1992 13308 2020
rect 8536 1980 8542 1992
rect 13280 1952 13308 1992
rect 14090 1980 14096 2032
rect 14148 2020 14154 2032
rect 17328 2020 17356 2060
rect 17862 2048 17868 2100
rect 17920 2088 17926 2100
rect 19426 2088 19432 2100
rect 17920 2060 19432 2088
rect 17920 2048 17926 2060
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 25222 2020 25228 2032
rect 14148 1992 16068 2020
rect 17328 1992 25228 2020
rect 14148 1980 14154 1992
rect 14458 1952 14464 1964
rect 13280 1924 14464 1952
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 12066 1844 12072 1896
rect 12124 1884 12130 1896
rect 15930 1884 15936 1896
rect 12124 1856 15936 1884
rect 12124 1844 12130 1856
rect 15930 1844 15936 1856
rect 15988 1844 15994 1896
rect 16040 1884 16068 1992
rect 25222 1980 25228 1992
rect 25280 1980 25286 2032
rect 20898 1952 20904 1964
rect 17328 1924 20904 1952
rect 17328 1884 17356 1924
rect 20898 1912 20904 1924
rect 20956 1912 20962 1964
rect 16040 1856 17356 1884
rect 18966 1844 18972 1896
rect 19024 1884 19030 1896
rect 24026 1884 24032 1896
rect 19024 1856 24032 1884
rect 19024 1844 19030 1856
rect 24026 1844 24032 1856
rect 24084 1844 24090 1896
rect 10962 1708 10968 1760
rect 11020 1748 11026 1760
rect 22278 1748 22284 1760
rect 11020 1720 22284 1748
rect 11020 1708 11026 1720
rect 22278 1708 22284 1720
rect 22336 1708 22342 1760
rect 15562 1640 15568 1692
rect 15620 1680 15626 1692
rect 21910 1680 21916 1692
rect 15620 1652 21916 1680
rect 15620 1640 15626 1652
rect 21910 1640 21916 1652
rect 21968 1640 21974 1692
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20 37272 72 37324
rect 1308 37204 1360 37256
rect 2780 37204 2832 37256
rect 3240 37204 3292 37256
rect 5448 37204 5500 37256
rect 6552 37247 6604 37256
rect 6552 37213 6561 37247
rect 6561 37213 6595 37247
rect 6595 37213 6604 37247
rect 6552 37204 6604 37213
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9036 37204 9088 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 12440 37204 12492 37256
rect 14280 37247 14332 37256
rect 14280 37213 14289 37247
rect 14289 37213 14323 37247
rect 14323 37213 14332 37247
rect 14280 37204 14332 37213
rect 15752 37204 15804 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18052 37204 18104 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 21272 37204 21324 37256
rect 22560 37204 22612 37256
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25780 37204 25832 37256
rect 27712 37204 27764 37256
rect 29000 37204 29052 37256
rect 30380 37204 30432 37256
rect 32220 37204 32272 37256
rect 33508 37204 33560 37256
rect 33968 37204 34020 37256
rect 34796 37204 34848 37256
rect 1584 37111 1636 37120
rect 1584 37077 1593 37111
rect 1593 37077 1627 37111
rect 1627 37077 1636 37111
rect 1584 37068 1636 37077
rect 5356 37136 5408 37188
rect 20352 37136 20404 37188
rect 2872 37111 2924 37120
rect 2872 37077 2881 37111
rect 2881 37077 2915 37111
rect 2915 37077 2924 37111
rect 2872 37068 2924 37077
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 4620 37068 4672 37120
rect 5816 37068 5868 37120
rect 7748 37068 7800 37120
rect 9312 37068 9364 37120
rect 10324 37068 10376 37120
rect 12348 37111 12400 37120
rect 12348 37077 12357 37111
rect 12357 37077 12391 37111
rect 12391 37077 12400 37111
rect 12348 37068 12400 37077
rect 13544 37068 13596 37120
rect 15476 37068 15528 37120
rect 16764 37068 16816 37120
rect 17132 37068 17184 37120
rect 19984 37068 20036 37120
rect 20444 37068 20496 37120
rect 23388 37136 23440 37188
rect 24492 37068 24544 37120
rect 29644 37136 29696 37188
rect 27620 37068 27672 37120
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 29828 37068 29880 37120
rect 32588 37136 32640 37188
rect 36728 37204 36780 37256
rect 32404 37068 32456 37120
rect 35348 37068 35400 37120
rect 38200 37111 38252 37120
rect 38200 37077 38209 37111
rect 38209 37077 38243 37111
rect 38243 37077 38252 37111
rect 38200 37068 38252 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1584 36864 1636 36916
rect 6460 36864 6512 36916
rect 6552 36864 6604 36916
rect 3976 36796 4028 36848
rect 9404 36796 9456 36848
rect 24860 36796 24912 36848
rect 29736 36796 29788 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 10692 36728 10744 36780
rect 39304 36796 39356 36848
rect 38016 36728 38068 36780
rect 2688 36524 2740 36576
rect 29276 36524 29328 36576
rect 38108 36567 38160 36576
rect 38108 36533 38117 36567
rect 38117 36533 38151 36567
rect 38151 36533 38160 36567
rect 38108 36524 38160 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 15752 36363 15804 36372
rect 15752 36329 15761 36363
rect 15761 36329 15795 36363
rect 15795 36329 15804 36363
rect 15752 36320 15804 36329
rect 15936 36159 15988 36168
rect 15936 36125 15945 36159
rect 15945 36125 15979 36159
rect 15979 36125 15988 36159
rect 15936 36116 15988 36125
rect 37188 36116 37240 36168
rect 35900 35980 35952 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 10692 35275 10744 35284
rect 10692 35241 10701 35275
rect 10701 35241 10735 35275
rect 10735 35241 10744 35275
rect 10692 35232 10744 35241
rect 12256 35028 12308 35080
rect 33876 35028 33928 35080
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 16856 34731 16908 34740
rect 16856 34697 16865 34731
rect 16865 34697 16899 34731
rect 16899 34697 16908 34731
rect 16856 34688 16908 34697
rect 24584 34688 24636 34740
rect 17040 34595 17092 34604
rect 17040 34561 17049 34595
rect 17049 34561 17083 34595
rect 17083 34561 17092 34595
rect 17040 34552 17092 34561
rect 23020 34595 23072 34604
rect 23020 34561 23029 34595
rect 23029 34561 23063 34595
rect 23063 34561 23072 34595
rect 23020 34552 23072 34561
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5448 34144 5500 34196
rect 10416 34144 10468 34196
rect 14280 34187 14332 34196
rect 14280 34153 14289 34187
rect 14289 34153 14323 34187
rect 14323 34153 14332 34187
rect 14280 34144 14332 34153
rect 8760 33940 8812 33992
rect 13636 33940 13688 33992
rect 14556 33872 14608 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 20076 33600 20128 33652
rect 3424 33464 3476 33516
rect 12348 33464 12400 33516
rect 19432 33464 19484 33516
rect 23388 33507 23440 33516
rect 23388 33473 23397 33507
rect 23397 33473 23431 33507
rect 23431 33473 23440 33507
rect 23388 33464 23440 33473
rect 24860 33507 24912 33516
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 37832 33464 37884 33516
rect 1768 33371 1820 33380
rect 1768 33337 1777 33371
rect 1777 33337 1811 33371
rect 1811 33337 1820 33371
rect 1768 33328 1820 33337
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 15660 33260 15712 33312
rect 22192 33260 22244 33312
rect 24952 33303 25004 33312
rect 24952 33269 24961 33303
rect 24961 33269 24995 33303
rect 24995 33269 25004 33303
rect 24952 33260 25004 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7840 33056 7892 33108
rect 11796 32852 11848 32904
rect 17132 32852 17184 32904
rect 32404 32988 32456 33040
rect 35348 32920 35400 32972
rect 38108 32852 38160 32904
rect 15108 32716 15160 32768
rect 28264 32759 28316 32768
rect 28264 32725 28273 32759
rect 28273 32725 28307 32759
rect 28307 32725 28316 32759
rect 28264 32716 28316 32725
rect 31116 32759 31168 32768
rect 31116 32725 31125 32759
rect 31125 32725 31159 32759
rect 31159 32725 31168 32759
rect 31116 32716 31168 32725
rect 31852 32716 31904 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15936 32512 15988 32564
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 5356 32376 5408 32428
rect 16948 32376 17000 32428
rect 20444 32444 20496 32496
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 38292 32419 38344 32428
rect 38292 32385 38301 32419
rect 38301 32385 38335 32419
rect 38335 32385 38344 32419
rect 38292 32376 38344 32385
rect 6736 32172 6788 32224
rect 7472 32215 7524 32224
rect 7472 32181 7481 32215
rect 7481 32181 7515 32215
rect 7515 32181 7524 32215
rect 7472 32172 7524 32181
rect 18052 32172 18104 32224
rect 20444 32215 20496 32224
rect 20444 32181 20453 32215
rect 20453 32181 20487 32215
rect 20487 32181 20496 32215
rect 20444 32172 20496 32181
rect 33232 32172 33284 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 33968 31968 34020 32020
rect 12256 31764 12308 31816
rect 12808 31764 12860 31816
rect 29000 31764 29052 31816
rect 35900 31832 35952 31884
rect 32220 31807 32272 31816
rect 32220 31773 32229 31807
rect 32229 31773 32263 31807
rect 32263 31773 32272 31807
rect 32220 31764 32272 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 5540 30812 5592 30864
rect 11336 30812 11388 30864
rect 19248 30812 19300 30864
rect 27620 30880 27672 30932
rect 33876 30923 33928 30932
rect 33876 30889 33885 30923
rect 33885 30889 33919 30923
rect 33919 30889 33928 30923
rect 33876 30880 33928 30889
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 2688 30676 2740 30728
rect 9312 30719 9364 30728
rect 9312 30685 9321 30719
rect 9321 30685 9355 30719
rect 9355 30685 9364 30719
rect 9312 30676 9364 30685
rect 9404 30676 9456 30728
rect 29828 30812 29880 30864
rect 32588 30744 32640 30796
rect 31760 30676 31812 30728
rect 29644 30608 29696 30660
rect 6092 30583 6144 30592
rect 6092 30549 6101 30583
rect 6101 30549 6135 30583
rect 6135 30549 6144 30583
rect 6092 30540 6144 30549
rect 11980 30540 12032 30592
rect 19984 30540 20036 30592
rect 25964 30583 26016 30592
rect 25964 30549 25973 30583
rect 25973 30549 26007 30583
rect 26007 30549 26016 30583
rect 25964 30540 26016 30549
rect 27804 30583 27856 30592
rect 27804 30549 27813 30583
rect 27813 30549 27847 30583
rect 27847 30549 27856 30583
rect 27804 30540 27856 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6460 30200 6512 30252
rect 29276 30243 29328 30252
rect 29276 30209 29285 30243
rect 29285 30209 29319 30243
rect 29319 30209 29328 30243
rect 29276 30200 29328 30209
rect 38292 30243 38344 30252
rect 38292 30209 38301 30243
rect 38301 30209 38335 30243
rect 38335 30209 38344 30243
rect 38292 30200 38344 30209
rect 11612 29996 11664 30048
rect 29368 30039 29420 30048
rect 29368 30005 29377 30039
rect 29377 30005 29411 30039
rect 29411 30005 29420 30039
rect 29368 29996 29420 30005
rect 36544 29996 36596 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 3424 29248 3476 29300
rect 23020 29248 23072 29300
rect 9312 29180 9364 29232
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 10140 29112 10192 29164
rect 22560 29155 22612 29164
rect 2872 29044 2924 29096
rect 22560 29121 22569 29155
rect 22569 29121 22603 29155
rect 22603 29121 22612 29155
rect 22560 29112 22612 29121
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 16856 28976 16908 29028
rect 38108 29019 38160 29028
rect 38108 28985 38117 29019
rect 38117 28985 38151 29019
rect 38151 28985 38160 29019
rect 38108 28976 38160 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 14556 28704 14608 28756
rect 17040 28704 17092 28756
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 17408 28432 17460 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8760 28203 8812 28212
rect 8760 28169 8769 28203
rect 8769 28169 8803 28203
rect 8803 28169 8812 28203
rect 8760 28160 8812 28169
rect 11796 28203 11848 28212
rect 11796 28169 11805 28203
rect 11805 28169 11839 28203
rect 11839 28169 11848 28203
rect 11796 28160 11848 28169
rect 13636 28203 13688 28212
rect 13636 28169 13645 28203
rect 13645 28169 13679 28203
rect 13679 28169 13688 28203
rect 13636 28160 13688 28169
rect 29000 28203 29052 28212
rect 29000 28169 29009 28203
rect 29009 28169 29043 28203
rect 29043 28169 29052 28203
rect 29000 28160 29052 28169
rect 11060 28024 11112 28076
rect 12716 28024 12768 28076
rect 13820 28024 13872 28076
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19432 27548 19484 27600
rect 3976 27412 4028 27464
rect 20076 27412 20128 27464
rect 33232 27455 33284 27464
rect 33232 27421 33241 27455
rect 33241 27421 33275 27455
rect 33275 27421 33284 27455
rect 33232 27412 33284 27421
rect 33508 27412 33560 27464
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 33324 27319 33376 27328
rect 33324 27285 33333 27319
rect 33333 27285 33367 27319
rect 33367 27285 33376 27319
rect 33324 27276 33376 27285
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 31760 27072 31812 27124
rect 6736 26936 6788 26988
rect 24768 26936 24820 26988
rect 8944 26732 8996 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5540 25848 5592 25900
rect 15568 25848 15620 25900
rect 17960 25848 18012 25900
rect 9588 25644 9640 25696
rect 17684 25687 17736 25696
rect 17684 25653 17693 25687
rect 17693 25653 17727 25687
rect 17727 25653 17736 25687
rect 17684 25644 17736 25653
rect 18972 25644 19024 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 12348 25236 12400 25288
rect 15292 25236 15344 25288
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 38108 25372 38160 25424
rect 36544 25304 36596 25356
rect 36912 25236 36964 25288
rect 4068 25100 4120 25152
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 18236 25100 18288 25152
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 19340 25100 19392 25152
rect 31760 25143 31812 25152
rect 31760 25109 31769 25143
rect 31769 25109 31803 25143
rect 31803 25109 31812 25143
rect 31760 25100 31812 25109
rect 32404 25143 32456 25152
rect 32404 25109 32413 25143
rect 32413 25109 32447 25143
rect 32447 25109 32456 25143
rect 32404 25100 32456 25109
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 6092 24760 6144 24812
rect 9772 24760 9824 24812
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 16304 24803 16356 24812
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 16304 24760 16356 24769
rect 18328 24803 18380 24812
rect 16580 24692 16632 24744
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 18972 24803 19024 24812
rect 17776 24692 17828 24744
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20812 24760 20864 24812
rect 22008 24760 22060 24812
rect 20628 24692 20680 24744
rect 27804 24692 27856 24744
rect 17960 24624 18012 24676
rect 19616 24624 19668 24676
rect 15844 24556 15896 24608
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 17500 24599 17552 24608
rect 17500 24565 17509 24599
rect 17509 24565 17543 24599
rect 17543 24565 17552 24599
rect 17500 24556 17552 24565
rect 19156 24599 19208 24608
rect 19156 24565 19165 24599
rect 19165 24565 19199 24599
rect 19199 24565 19208 24599
rect 19156 24556 19208 24565
rect 20352 24599 20404 24608
rect 20352 24565 20361 24599
rect 20361 24565 20395 24599
rect 20395 24565 20404 24599
rect 20352 24556 20404 24565
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 16304 24352 16356 24404
rect 16764 24352 16816 24404
rect 15936 24216 15988 24268
rect 6184 24148 6236 24200
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 15568 24148 15620 24157
rect 16304 24148 16356 24200
rect 19156 24352 19208 24404
rect 33508 24395 33560 24404
rect 33508 24361 33517 24395
rect 33517 24361 33551 24395
rect 33551 24361 33560 24395
rect 33508 24352 33560 24361
rect 31116 24284 31168 24336
rect 17684 24216 17736 24268
rect 18604 24216 18656 24268
rect 20352 24216 20404 24268
rect 17500 24148 17552 24200
rect 20720 24148 20772 24200
rect 30380 24148 30432 24200
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 18696 24080 18748 24132
rect 19616 24123 19668 24132
rect 19616 24089 19625 24123
rect 19625 24089 19659 24123
rect 19659 24089 19668 24123
rect 20168 24123 20220 24132
rect 19616 24080 19668 24089
rect 20168 24089 20177 24123
rect 20177 24089 20211 24123
rect 20211 24089 20220 24123
rect 20168 24080 20220 24089
rect 22376 24080 22428 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 16488 24012 16540 24064
rect 20904 24012 20956 24064
rect 37004 24012 37056 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3976 23851 4028 23860
rect 3976 23817 3985 23851
rect 3985 23817 4019 23851
rect 4019 23817 4028 23851
rect 3976 23808 4028 23817
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 19340 23783 19392 23792
rect 5540 23672 5592 23724
rect 14004 23672 14056 23724
rect 19340 23749 19349 23783
rect 19349 23749 19383 23783
rect 19383 23749 19392 23783
rect 19340 23740 19392 23749
rect 20168 23808 20220 23860
rect 24768 23808 24820 23860
rect 20904 23783 20956 23792
rect 20904 23749 20913 23783
rect 20913 23749 20947 23783
rect 20947 23749 20956 23783
rect 20904 23740 20956 23749
rect 22560 23740 22612 23792
rect 15660 23715 15712 23724
rect 12992 23647 13044 23656
rect 12992 23613 13001 23647
rect 13001 23613 13035 23647
rect 13035 23613 13044 23647
rect 12992 23604 13044 23613
rect 14096 23604 14148 23656
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 16120 23672 16172 23724
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 15292 23604 15344 23656
rect 16028 23604 16080 23656
rect 16672 23536 16724 23588
rect 16856 23647 16908 23656
rect 16856 23613 16865 23647
rect 16865 23613 16899 23647
rect 16899 23613 16908 23647
rect 16856 23604 16908 23613
rect 17132 23604 17184 23656
rect 13728 23511 13780 23520
rect 13728 23477 13737 23511
rect 13737 23477 13771 23511
rect 13771 23477 13780 23511
rect 13728 23468 13780 23477
rect 15568 23468 15620 23520
rect 16488 23468 16540 23520
rect 22100 23511 22152 23520
rect 22100 23477 22109 23511
rect 22109 23477 22143 23511
rect 22143 23477 22152 23511
rect 22100 23468 22152 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 9220 23264 9272 23316
rect 16580 23264 16632 23316
rect 16764 23264 16816 23316
rect 18696 23307 18748 23316
rect 18696 23273 18705 23307
rect 18705 23273 18739 23307
rect 18739 23273 18748 23307
rect 18696 23264 18748 23273
rect 14464 23060 14516 23112
rect 17132 23196 17184 23248
rect 17868 23196 17920 23248
rect 19432 23196 19484 23248
rect 16672 23171 16724 23180
rect 16672 23137 16681 23171
rect 16681 23137 16715 23171
rect 16715 23137 16724 23171
rect 16672 23128 16724 23137
rect 16856 23128 16908 23180
rect 17684 23128 17736 23180
rect 18236 23171 18288 23180
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 24952 23264 25004 23316
rect 21272 23196 21324 23248
rect 21088 23128 21140 23180
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 22376 23171 22428 23180
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 13452 22992 13504 23044
rect 15752 22992 15804 23044
rect 17316 23060 17368 23112
rect 22560 23060 22612 23112
rect 17592 22992 17644 23044
rect 13176 22924 13228 22976
rect 14280 22924 14332 22976
rect 19248 22924 19300 22976
rect 22100 22992 22152 23044
rect 21272 22924 21324 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 5540 22763 5592 22772
rect 5540 22729 5549 22763
rect 5549 22729 5583 22763
rect 5583 22729 5592 22763
rect 5540 22720 5592 22729
rect 18328 22720 18380 22772
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 36912 22720 36964 22772
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 10416 22652 10468 22704
rect 16764 22652 16816 22704
rect 21364 22652 21416 22704
rect 9312 22627 9364 22636
rect 9312 22593 9321 22627
rect 9321 22593 9355 22627
rect 9355 22593 9364 22627
rect 9312 22584 9364 22593
rect 9680 22584 9732 22636
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 13084 22584 13136 22593
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 14924 22584 14976 22636
rect 16304 22627 16356 22636
rect 16304 22593 16313 22627
rect 16313 22593 16347 22627
rect 16347 22593 16356 22627
rect 16304 22584 16356 22593
rect 17408 22627 17460 22636
rect 17408 22593 17417 22627
rect 17417 22593 17451 22627
rect 17451 22593 17460 22627
rect 17408 22584 17460 22593
rect 21824 22584 21876 22636
rect 21916 22584 21968 22636
rect 33140 22627 33192 22636
rect 33140 22593 33149 22627
rect 33149 22593 33183 22627
rect 33183 22593 33192 22627
rect 33140 22584 33192 22593
rect 10232 22516 10284 22568
rect 12900 22516 12952 22568
rect 17684 22516 17736 22568
rect 19524 22559 19576 22568
rect 19524 22525 19533 22559
rect 19533 22525 19567 22559
rect 19567 22525 19576 22559
rect 19524 22516 19576 22525
rect 19984 22516 20036 22568
rect 20628 22559 20680 22568
rect 20628 22525 20637 22559
rect 20637 22525 20671 22559
rect 20671 22525 20680 22559
rect 20628 22516 20680 22525
rect 10876 22448 10928 22500
rect 5540 22380 5592 22432
rect 10324 22380 10376 22432
rect 14556 22448 14608 22500
rect 13912 22380 13964 22432
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 14188 22380 14240 22389
rect 15660 22380 15712 22432
rect 18236 22448 18288 22500
rect 17040 22380 17092 22432
rect 17408 22380 17460 22432
rect 17776 22380 17828 22432
rect 18420 22380 18472 22432
rect 19248 22380 19300 22432
rect 21640 22380 21692 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 13084 22176 13136 22228
rect 17316 22219 17368 22228
rect 17316 22185 17325 22219
rect 17325 22185 17359 22219
rect 17359 22185 17368 22219
rect 17316 22176 17368 22185
rect 20720 22176 20772 22228
rect 21824 22219 21876 22228
rect 21824 22185 21833 22219
rect 21833 22185 21867 22219
rect 21867 22185 21876 22219
rect 21824 22176 21876 22185
rect 9680 21972 9732 22024
rect 10048 22108 10100 22160
rect 15936 22108 15988 22160
rect 16672 22108 16724 22160
rect 11796 22040 11848 22092
rect 12900 22040 12952 22092
rect 13268 22040 13320 22092
rect 14464 22040 14516 22092
rect 15568 22083 15620 22092
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 19524 22108 19576 22160
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18236 22040 18288 22049
rect 8484 21904 8536 21956
rect 10784 21972 10836 22024
rect 9128 21879 9180 21888
rect 9128 21845 9137 21879
rect 9137 21845 9171 21879
rect 9171 21845 9180 21879
rect 9128 21836 9180 21845
rect 11244 21904 11296 21956
rect 12072 21972 12124 22024
rect 14004 21972 14056 22024
rect 14280 21972 14332 22024
rect 15384 21972 15436 22024
rect 16856 21972 16908 22024
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 19984 21972 20036 22024
rect 28264 22040 28316 22092
rect 21456 21972 21508 22024
rect 13176 21947 13228 21956
rect 13176 21913 13185 21947
rect 13185 21913 13219 21947
rect 13219 21913 13228 21947
rect 13176 21904 13228 21913
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 11428 21836 11480 21888
rect 12348 21836 12400 21888
rect 15752 21904 15804 21956
rect 15936 21904 15988 21956
rect 18144 21904 18196 21956
rect 20076 21904 20128 21956
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 21548 21904 21600 21956
rect 30380 21972 30432 22024
rect 38108 21947 38160 21956
rect 38108 21913 38117 21947
rect 38117 21913 38151 21947
rect 38151 21913 38160 21947
rect 38108 21904 38160 21913
rect 14004 21836 14056 21888
rect 16304 21836 16356 21888
rect 21916 21836 21968 21888
rect 37924 21836 37976 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4068 21496 4120 21548
rect 9128 21496 9180 21548
rect 9312 21539 9364 21548
rect 9312 21505 9321 21539
rect 9321 21505 9355 21539
rect 9355 21505 9364 21539
rect 9312 21496 9364 21505
rect 10232 21564 10284 21616
rect 10692 21564 10744 21616
rect 13176 21632 13228 21684
rect 13084 21564 13136 21616
rect 14188 21632 14240 21684
rect 13912 21607 13964 21616
rect 13912 21573 13921 21607
rect 13921 21573 13955 21607
rect 13955 21573 13964 21607
rect 13912 21564 13964 21573
rect 18052 21632 18104 21684
rect 18144 21632 18196 21684
rect 23112 21632 23164 21684
rect 16764 21564 16816 21616
rect 17040 21607 17092 21616
rect 17040 21573 17049 21607
rect 17049 21573 17083 21607
rect 17083 21573 17092 21607
rect 17040 21564 17092 21573
rect 17592 21607 17644 21616
rect 17592 21573 17601 21607
rect 17601 21573 17635 21607
rect 17635 21573 17644 21607
rect 17592 21564 17644 21573
rect 10232 21360 10284 21412
rect 10784 21360 10836 21412
rect 11060 21403 11112 21412
rect 11060 21369 11069 21403
rect 11069 21369 11103 21403
rect 11103 21369 11112 21403
rect 11060 21360 11112 21369
rect 15660 21539 15712 21548
rect 15660 21505 15669 21539
rect 15669 21505 15703 21539
rect 15703 21505 15712 21539
rect 15660 21496 15712 21505
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 19248 21539 19300 21548
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 31760 21564 31812 21616
rect 14004 21428 14056 21480
rect 4712 21292 4764 21344
rect 9680 21292 9732 21344
rect 12164 21292 12216 21344
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12440 21292 12492 21301
rect 16764 21292 16816 21344
rect 18420 21428 18472 21480
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 20904 21292 20956 21344
rect 22652 21292 22704 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6184 21088 6236 21140
rect 9588 21088 9640 21140
rect 10692 21063 10744 21072
rect 10692 21029 10701 21063
rect 10701 21029 10735 21063
rect 10735 21029 10744 21063
rect 10692 21020 10744 21029
rect 11152 20952 11204 21004
rect 14740 21063 14792 21072
rect 14740 21029 14749 21063
rect 14749 21029 14783 21063
rect 14783 21029 14792 21063
rect 14740 21020 14792 21029
rect 17040 21088 17092 21140
rect 18328 21088 18380 21140
rect 19432 21088 19484 21140
rect 21456 21088 21508 21140
rect 21732 21088 21784 21140
rect 19984 21020 20036 21072
rect 20996 21020 21048 21072
rect 13728 20952 13780 21004
rect 14372 20995 14424 21004
rect 14372 20961 14381 20995
rect 14381 20961 14415 20995
rect 14415 20961 14424 20995
rect 14372 20952 14424 20961
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 15936 20927 15988 20936
rect 8668 20816 8720 20868
rect 11704 20816 11756 20868
rect 5816 20748 5868 20800
rect 7472 20748 7524 20800
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 18512 20884 18564 20936
rect 18788 20884 18840 20936
rect 20812 20952 20864 21004
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 21088 20884 21140 20936
rect 23112 20927 23164 20936
rect 12440 20816 12492 20868
rect 16488 20816 16540 20868
rect 12072 20748 12124 20800
rect 17040 20748 17092 20800
rect 17224 20859 17276 20868
rect 17224 20825 17233 20859
rect 17233 20825 17267 20859
rect 17267 20825 17276 20859
rect 17224 20816 17276 20825
rect 17592 20816 17644 20868
rect 21732 20816 21784 20868
rect 23112 20893 23121 20927
rect 23121 20893 23155 20927
rect 23155 20893 23164 20927
rect 23112 20884 23164 20893
rect 25504 20884 25556 20936
rect 33600 20884 33652 20936
rect 19432 20748 19484 20800
rect 22100 20748 22152 20800
rect 33140 20748 33192 20800
rect 38200 20791 38252 20800
rect 38200 20757 38209 20791
rect 38209 20757 38243 20791
rect 38243 20757 38252 20791
rect 38200 20748 38252 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 7932 20544 7984 20596
rect 11244 20544 11296 20596
rect 10324 20519 10376 20528
rect 10324 20485 10333 20519
rect 10333 20485 10367 20519
rect 10367 20485 10376 20519
rect 10324 20476 10376 20485
rect 11060 20476 11112 20528
rect 12164 20519 12216 20528
rect 12164 20485 12173 20519
rect 12173 20485 12207 20519
rect 12207 20485 12216 20519
rect 12164 20476 12216 20485
rect 12256 20476 12308 20528
rect 18604 20544 18656 20596
rect 16488 20476 16540 20528
rect 17316 20476 17368 20528
rect 18880 20519 18932 20528
rect 18880 20485 18889 20519
rect 18889 20485 18923 20519
rect 18923 20485 18932 20519
rect 19984 20519 20036 20528
rect 18880 20476 18932 20485
rect 19984 20485 19993 20519
rect 19993 20485 20027 20519
rect 20027 20485 20036 20519
rect 19984 20476 20036 20485
rect 20720 20544 20772 20596
rect 21272 20476 21324 20528
rect 21548 20476 21600 20528
rect 6920 20451 6972 20460
rect 6920 20417 6929 20451
rect 6929 20417 6963 20451
rect 6963 20417 6972 20451
rect 6920 20408 6972 20417
rect 3332 20340 3384 20392
rect 8392 20408 8444 20460
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 21088 20451 21140 20460
rect 9312 20340 9364 20392
rect 10324 20340 10376 20392
rect 10416 20340 10468 20392
rect 10600 20272 10652 20324
rect 12348 20340 12400 20392
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 12532 20272 12584 20324
rect 13820 20315 13872 20324
rect 13820 20281 13829 20315
rect 13829 20281 13863 20315
rect 13863 20281 13872 20315
rect 13820 20272 13872 20281
rect 14924 20272 14976 20324
rect 17040 20340 17092 20392
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 9404 20204 9456 20256
rect 11520 20204 11572 20256
rect 11704 20204 11756 20256
rect 12256 20204 12308 20256
rect 12440 20204 12492 20256
rect 15660 20204 15712 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 17684 20272 17736 20324
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 23020 20408 23072 20460
rect 20996 20340 21048 20392
rect 22652 20340 22704 20392
rect 19340 20315 19392 20324
rect 19340 20281 19349 20315
rect 19349 20281 19383 20315
rect 19383 20281 19392 20315
rect 19340 20272 19392 20281
rect 20168 20272 20220 20324
rect 15752 20204 15804 20213
rect 20076 20204 20128 20256
rect 20904 20204 20956 20256
rect 23204 20204 23256 20256
rect 23296 20247 23348 20256
rect 23296 20213 23305 20247
rect 23305 20213 23339 20247
rect 23339 20213 23348 20247
rect 23296 20204 23348 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 9956 20000 10008 20052
rect 10692 20000 10744 20052
rect 15292 20000 15344 20052
rect 15660 20000 15712 20052
rect 7012 19932 7064 19984
rect 17132 20000 17184 20052
rect 19432 20000 19484 20052
rect 19984 20000 20036 20052
rect 20996 20000 21048 20052
rect 9772 19864 9824 19916
rect 5540 19796 5592 19848
rect 8392 19796 8444 19848
rect 9036 19728 9088 19780
rect 8484 19660 8536 19712
rect 8576 19660 8628 19712
rect 9128 19660 9180 19712
rect 9312 19796 9364 19848
rect 12440 19864 12492 19916
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 14740 19864 14792 19916
rect 16212 19907 16264 19916
rect 16212 19873 16221 19907
rect 16221 19873 16255 19907
rect 16255 19873 16264 19907
rect 16212 19864 16264 19873
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 14280 19796 14332 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 16304 19796 16356 19848
rect 17592 19864 17644 19916
rect 19248 19864 19300 19916
rect 18420 19839 18472 19848
rect 9404 19728 9456 19780
rect 15200 19771 15252 19780
rect 15200 19737 15209 19771
rect 15209 19737 15243 19771
rect 15243 19737 15252 19771
rect 15200 19728 15252 19737
rect 15476 19728 15528 19780
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 19432 19796 19484 19848
rect 18696 19728 18748 19780
rect 10048 19660 10100 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 13544 19660 13596 19669
rect 15844 19660 15896 19712
rect 18236 19660 18288 19712
rect 32220 19932 32272 19984
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 32404 19864 32456 19916
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 37004 19796 37056 19848
rect 22008 19771 22060 19780
rect 22008 19737 22017 19771
rect 22017 19737 22051 19771
rect 22051 19737 22060 19771
rect 22008 19728 22060 19737
rect 24952 19728 25004 19780
rect 22192 19660 22244 19712
rect 27620 19660 27672 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5172 19456 5224 19508
rect 9588 19456 9640 19508
rect 12348 19499 12400 19508
rect 12348 19465 12357 19499
rect 12357 19465 12391 19499
rect 12391 19465 12400 19499
rect 12348 19456 12400 19465
rect 15936 19456 15988 19508
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 8484 19388 8536 19440
rect 6920 19320 6972 19329
rect 8576 19320 8628 19372
rect 8208 19252 8260 19304
rect 9772 19388 9824 19440
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 9864 19320 9916 19372
rect 11336 19320 11388 19372
rect 12992 19363 13044 19372
rect 8760 19184 8812 19236
rect 11612 19252 11664 19304
rect 11796 19252 11848 19304
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 10324 19227 10376 19236
rect 10324 19193 10333 19227
rect 10333 19193 10367 19227
rect 10367 19193 10376 19227
rect 10324 19184 10376 19193
rect 10600 19184 10652 19236
rect 15200 19252 15252 19304
rect 17960 19388 18012 19440
rect 16856 19320 16908 19372
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 23296 19456 23348 19508
rect 18972 19320 19024 19372
rect 20444 19320 20496 19372
rect 31852 19388 31904 19440
rect 17224 19295 17276 19304
rect 13912 19184 13964 19236
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 19248 19252 19300 19304
rect 19524 19295 19576 19304
rect 19524 19261 19533 19295
rect 19533 19261 19567 19295
rect 19567 19261 19576 19295
rect 19524 19252 19576 19261
rect 23204 19320 23256 19372
rect 22008 19295 22060 19304
rect 9312 19159 9364 19168
rect 9312 19125 9321 19159
rect 9321 19125 9355 19159
rect 9355 19125 9364 19159
rect 9312 19116 9364 19125
rect 9680 19116 9732 19168
rect 13268 19116 13320 19168
rect 13452 19116 13504 19168
rect 17592 19184 17644 19236
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 22100 19184 22152 19236
rect 15752 19116 15804 19168
rect 15936 19159 15988 19168
rect 15936 19125 15945 19159
rect 15945 19125 15979 19159
rect 15979 19125 15988 19159
rect 15936 19116 15988 19125
rect 18328 19116 18380 19168
rect 23020 19116 23072 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8760 18912 8812 18964
rect 10324 18912 10376 18964
rect 13912 18912 13964 18964
rect 14648 18912 14700 18964
rect 16120 18912 16172 18964
rect 17316 18912 17368 18964
rect 6920 18776 6972 18828
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 7288 18708 7340 18760
rect 13452 18844 13504 18896
rect 13820 18844 13872 18896
rect 15200 18844 15252 18896
rect 8484 18776 8536 18828
rect 9588 18776 9640 18828
rect 11796 18776 11848 18828
rect 9680 18708 9732 18760
rect 11336 18708 11388 18760
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12256 18708 12308 18717
rect 12624 18776 12676 18828
rect 15476 18844 15528 18896
rect 15752 18844 15804 18896
rect 17592 18887 17644 18896
rect 17592 18853 17601 18887
rect 17601 18853 17635 18887
rect 17635 18853 17644 18887
rect 17592 18844 17644 18853
rect 15108 18708 15160 18760
rect 16396 18776 16448 18828
rect 18972 18912 19024 18964
rect 20260 18912 20312 18964
rect 33600 18955 33652 18964
rect 33600 18921 33609 18955
rect 33609 18921 33643 18955
rect 33643 18921 33652 18955
rect 33600 18912 33652 18921
rect 19432 18776 19484 18828
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 16856 18708 16908 18760
rect 8300 18572 8352 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 8576 18572 8628 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12624 18572 12676 18624
rect 13360 18640 13412 18692
rect 16672 18640 16724 18692
rect 17132 18683 17184 18692
rect 17132 18649 17141 18683
rect 17141 18649 17175 18683
rect 17175 18649 17184 18683
rect 17132 18640 17184 18649
rect 17960 18640 18012 18692
rect 19340 18708 19392 18760
rect 25964 18844 26016 18896
rect 20812 18819 20864 18828
rect 20812 18785 20821 18819
rect 20821 18785 20855 18819
rect 20855 18785 20864 18819
rect 20812 18776 20864 18785
rect 22008 18776 22060 18828
rect 28908 18776 28960 18828
rect 22192 18708 22244 18760
rect 33416 18708 33468 18760
rect 13268 18572 13320 18624
rect 14280 18572 14332 18624
rect 16212 18572 16264 18624
rect 20628 18683 20680 18692
rect 20628 18649 20637 18683
rect 20637 18649 20671 18683
rect 20671 18649 20680 18683
rect 20628 18640 20680 18649
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 6644 18368 6696 18420
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 7288 18232 7340 18284
rect 8392 18232 8444 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 9036 18164 9088 18216
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 16028 18368 16080 18420
rect 18420 18411 18472 18420
rect 18420 18377 18429 18411
rect 18429 18377 18463 18411
rect 18463 18377 18472 18411
rect 18420 18368 18472 18377
rect 19984 18368 20036 18420
rect 20628 18368 20680 18420
rect 33416 18411 33468 18420
rect 12624 18300 12676 18352
rect 19248 18300 19300 18352
rect 20260 18343 20312 18352
rect 20260 18309 20269 18343
rect 20269 18309 20303 18343
rect 20303 18309 20312 18343
rect 20260 18300 20312 18309
rect 20812 18343 20864 18352
rect 20812 18309 20821 18343
rect 20821 18309 20855 18343
rect 20855 18309 20864 18343
rect 20812 18300 20864 18309
rect 16120 18275 16172 18284
rect 11704 18164 11756 18216
rect 12348 18164 12400 18216
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 13452 18164 13504 18216
rect 9588 18096 9640 18148
rect 9772 18139 9824 18148
rect 9772 18105 9781 18139
rect 9781 18105 9815 18139
rect 9815 18105 9824 18139
rect 9772 18096 9824 18105
rect 10048 18096 10100 18148
rect 11796 18096 11848 18148
rect 5540 18028 5592 18080
rect 11152 18028 11204 18080
rect 12440 18028 12492 18080
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 17040 18207 17092 18216
rect 14280 18096 14332 18148
rect 16396 18096 16448 18148
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 18880 18164 18932 18216
rect 17408 18096 17460 18148
rect 33416 18377 33425 18411
rect 33425 18377 33459 18411
rect 33459 18377 33468 18411
rect 33416 18368 33468 18377
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22652 18275 22704 18284
rect 22652 18241 22661 18275
rect 22661 18241 22695 18275
rect 22695 18241 22704 18275
rect 22652 18232 22704 18241
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 17868 18028 17920 18080
rect 18420 18028 18472 18080
rect 19708 18028 19760 18080
rect 22100 18096 22152 18148
rect 23388 18071 23440 18080
rect 23388 18037 23397 18071
rect 23397 18037 23431 18071
rect 23431 18037 23440 18071
rect 23388 18028 23440 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8668 17824 8720 17876
rect 8852 17824 8904 17876
rect 9588 17824 9640 17876
rect 10968 17824 11020 17876
rect 11704 17867 11756 17876
rect 11704 17833 11713 17867
rect 11713 17833 11747 17867
rect 11747 17833 11756 17867
rect 11704 17824 11756 17833
rect 12072 17824 12124 17876
rect 12440 17824 12492 17876
rect 17224 17824 17276 17876
rect 19432 17824 19484 17876
rect 8300 17756 8352 17808
rect 8944 17688 8996 17740
rect 9588 17688 9640 17740
rect 9956 17731 10008 17740
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 10048 17688 10100 17740
rect 18052 17756 18104 17808
rect 23388 17824 23440 17876
rect 12808 17688 12860 17740
rect 13084 17688 13136 17740
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 7656 17620 7708 17672
rect 8668 17620 8720 17672
rect 9036 17620 9088 17672
rect 11980 17620 12032 17672
rect 13820 17688 13872 17740
rect 21272 17756 21324 17808
rect 19432 17688 19484 17740
rect 9128 17552 9180 17604
rect 9220 17552 9272 17604
rect 10324 17552 10376 17604
rect 11612 17552 11664 17604
rect 12900 17552 12952 17604
rect 6920 17484 6972 17536
rect 11060 17484 11112 17536
rect 11152 17484 11204 17536
rect 16212 17620 16264 17672
rect 17960 17620 18012 17672
rect 19800 17620 19852 17672
rect 20260 17620 20312 17672
rect 16580 17552 16632 17604
rect 17868 17552 17920 17604
rect 15568 17527 15620 17536
rect 15568 17493 15577 17527
rect 15577 17493 15611 17527
rect 15611 17493 15620 17527
rect 15568 17484 15620 17493
rect 17960 17484 18012 17536
rect 21272 17620 21324 17672
rect 27620 17756 27672 17808
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 21824 17620 21876 17672
rect 22744 17527 22796 17536
rect 22744 17493 22753 17527
rect 22753 17493 22787 17527
rect 22787 17493 22796 17527
rect 22744 17484 22796 17493
rect 23480 17484 23532 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 8576 17144 8628 17196
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9772 17144 9824 17196
rect 10968 17212 11020 17264
rect 12808 17212 12860 17264
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 16856 17280 16908 17332
rect 19432 17323 19484 17332
rect 19432 17289 19441 17323
rect 19441 17289 19475 17323
rect 19475 17289 19484 17323
rect 19432 17280 19484 17289
rect 20260 17280 20312 17332
rect 15292 17255 15344 17264
rect 15292 17221 15301 17255
rect 15301 17221 15335 17255
rect 15335 17221 15344 17255
rect 15292 17212 15344 17221
rect 15568 17212 15620 17264
rect 20076 17255 20128 17264
rect 16304 17144 16356 17196
rect 20076 17221 20085 17255
rect 20085 17221 20119 17255
rect 20119 17221 20128 17255
rect 20076 17212 20128 17221
rect 8300 17076 8352 17128
rect 9404 17076 9456 17128
rect 9588 17076 9640 17128
rect 11888 17076 11940 17128
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 14832 17008 14884 17060
rect 16120 17076 16172 17128
rect 20628 17144 20680 17196
rect 21640 17144 21692 17196
rect 22744 17144 22796 17196
rect 34520 17144 34572 17196
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 20444 17076 20496 17128
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 23296 17119 23348 17128
rect 23296 17085 23305 17119
rect 23305 17085 23339 17119
rect 23339 17085 23348 17119
rect 23296 17076 23348 17085
rect 18604 17008 18656 17060
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 12532 16940 12584 16992
rect 16120 16940 16172 16992
rect 17960 16983 18012 16992
rect 17960 16949 17969 16983
rect 17969 16949 18003 16983
rect 18003 16949 18012 16983
rect 17960 16940 18012 16949
rect 23388 16940 23440 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 9220 16736 9272 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 9772 16736 9824 16788
rect 16304 16736 16356 16788
rect 17224 16736 17276 16788
rect 21272 16736 21324 16788
rect 21732 16736 21784 16788
rect 23296 16779 23348 16788
rect 23296 16745 23305 16779
rect 23305 16745 23339 16779
rect 23339 16745 23348 16779
rect 23296 16736 23348 16745
rect 8760 16668 8812 16720
rect 15200 16711 15252 16720
rect 9404 16600 9456 16652
rect 10324 16600 10376 16652
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7932 16575 7984 16584
rect 7104 16532 7156 16541
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8944 16532 8996 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 10692 16600 10744 16652
rect 10876 16600 10928 16652
rect 11612 16600 11664 16652
rect 12624 16600 12676 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 13084 16600 13136 16652
rect 15200 16677 15209 16711
rect 15209 16677 15243 16711
rect 15243 16677 15252 16711
rect 15200 16668 15252 16677
rect 17408 16711 17460 16720
rect 17408 16677 17417 16711
rect 17417 16677 17451 16711
rect 17451 16677 17460 16711
rect 17408 16668 17460 16677
rect 18880 16668 18932 16720
rect 7656 16464 7708 16516
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 14740 16532 14792 16584
rect 15016 16575 15068 16584
rect 11244 16507 11296 16516
rect 11244 16473 11253 16507
rect 11253 16473 11287 16507
rect 11287 16473 11296 16507
rect 11244 16464 11296 16473
rect 11796 16507 11848 16516
rect 11796 16473 11805 16507
rect 11805 16473 11839 16507
rect 11839 16473 11848 16507
rect 11796 16464 11848 16473
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 16764 16600 16816 16652
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16580 16532 16632 16541
rect 16948 16532 17000 16584
rect 17960 16600 18012 16652
rect 18236 16643 18288 16652
rect 18236 16609 18245 16643
rect 18245 16609 18279 16643
rect 18279 16609 18288 16643
rect 18236 16600 18288 16609
rect 18604 16643 18656 16652
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 20628 16668 20680 16720
rect 20720 16668 20772 16720
rect 22008 16668 22060 16720
rect 20996 16532 21048 16584
rect 23112 16600 23164 16652
rect 24860 16600 24912 16652
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 12440 16464 12492 16473
rect 15384 16464 15436 16516
rect 18328 16507 18380 16516
rect 18328 16473 18337 16507
rect 18337 16473 18371 16507
rect 18371 16473 18380 16507
rect 18328 16464 18380 16473
rect 19340 16464 19392 16516
rect 20352 16507 20404 16516
rect 20352 16473 20361 16507
rect 20361 16473 20395 16507
rect 20395 16473 20404 16507
rect 20352 16464 20404 16473
rect 13360 16396 13412 16448
rect 13820 16396 13872 16448
rect 15108 16396 15160 16448
rect 21548 16396 21600 16448
rect 34520 16396 34572 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 7932 16192 7984 16244
rect 8576 16192 8628 16244
rect 11428 16192 11480 16244
rect 11520 16192 11572 16244
rect 12440 16192 12492 16244
rect 15200 16235 15252 16244
rect 15200 16201 15209 16235
rect 15209 16201 15243 16235
rect 15243 16201 15252 16235
rect 15200 16192 15252 16201
rect 16672 16192 16724 16244
rect 17040 16192 17092 16244
rect 17684 16192 17736 16244
rect 20352 16192 20404 16244
rect 4804 16056 4856 16108
rect 4896 16056 4948 16108
rect 7104 16056 7156 16108
rect 7656 16056 7708 16108
rect 10416 16124 10468 16176
rect 9864 16099 9916 16108
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 10232 16056 10284 16108
rect 10784 16056 10836 16108
rect 11336 16056 11388 16108
rect 11796 16124 11848 16176
rect 12808 16124 12860 16176
rect 16948 16124 17000 16176
rect 19432 16124 19484 16176
rect 20904 16167 20956 16176
rect 20904 16133 20913 16167
rect 20913 16133 20947 16167
rect 20947 16133 20956 16167
rect 20904 16124 20956 16133
rect 16580 16056 16632 16108
rect 9772 15988 9824 16040
rect 10600 15988 10652 16040
rect 11612 15988 11664 16040
rect 11796 15988 11848 16040
rect 8024 15920 8076 15972
rect 9864 15920 9916 15972
rect 10416 15963 10468 15972
rect 10416 15929 10425 15963
rect 10425 15929 10459 15963
rect 10459 15929 10468 15963
rect 10416 15920 10468 15929
rect 11060 15920 11112 15972
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 14188 15988 14240 16040
rect 14648 15988 14700 16040
rect 15384 15988 15436 16040
rect 17040 16031 17092 16040
rect 12624 15920 12676 15972
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 18788 15988 18840 16040
rect 19984 15988 20036 16040
rect 17500 15920 17552 15972
rect 18052 15920 18104 15972
rect 24860 16124 24912 16176
rect 22836 16099 22888 16108
rect 22836 16065 22845 16099
rect 22845 16065 22879 16099
rect 22879 16065 22888 16099
rect 22836 16056 22888 16065
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 23112 15988 23164 16040
rect 24032 15988 24084 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 7840 15895 7892 15904
rect 7840 15861 7849 15895
rect 7849 15861 7883 15895
rect 7883 15861 7892 15895
rect 7840 15852 7892 15861
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 10140 15852 10192 15904
rect 10508 15852 10560 15904
rect 10876 15852 10928 15904
rect 11796 15852 11848 15904
rect 11980 15852 12032 15904
rect 12532 15895 12584 15904
rect 12532 15861 12541 15895
rect 12541 15861 12575 15895
rect 12575 15861 12584 15895
rect 12532 15852 12584 15861
rect 21548 15852 21600 15904
rect 22192 15852 22244 15904
rect 23296 15852 23348 15904
rect 37004 15852 37056 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8300 15648 8352 15700
rect 9588 15648 9640 15700
rect 13176 15648 13228 15700
rect 14188 15648 14240 15700
rect 16672 15691 16724 15700
rect 7840 15580 7892 15632
rect 10692 15512 10744 15564
rect 11520 15512 11572 15564
rect 11980 15580 12032 15632
rect 12716 15580 12768 15632
rect 14280 15580 14332 15632
rect 14372 15580 14424 15632
rect 15936 15580 15988 15632
rect 13084 15512 13136 15564
rect 13912 15512 13964 15564
rect 16672 15657 16681 15691
rect 16681 15657 16715 15691
rect 16715 15657 16724 15691
rect 16672 15648 16724 15657
rect 18972 15648 19024 15700
rect 24124 15648 24176 15700
rect 17500 15580 17552 15632
rect 19340 15512 19392 15564
rect 33324 15580 33376 15632
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 23296 15555 23348 15564
rect 23296 15521 23305 15555
rect 23305 15521 23339 15555
rect 23339 15521 23348 15555
rect 23296 15512 23348 15521
rect 5540 15444 5592 15496
rect 8208 15444 8260 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 7196 15376 7248 15428
rect 9680 15444 9732 15496
rect 9772 15444 9824 15496
rect 9864 15444 9916 15496
rect 11152 15444 11204 15496
rect 12072 15444 12124 15496
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 22100 15444 22152 15496
rect 25136 15444 25188 15496
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 9128 15308 9180 15360
rect 9772 15351 9824 15360
rect 9772 15317 9781 15351
rect 9781 15317 9815 15351
rect 9815 15317 9824 15351
rect 9772 15308 9824 15317
rect 12532 15376 12584 15428
rect 14372 15419 14424 15428
rect 11520 15308 11572 15360
rect 12164 15308 12216 15360
rect 14372 15385 14381 15419
rect 14381 15385 14415 15419
rect 14415 15385 14424 15419
rect 14372 15376 14424 15385
rect 13728 15308 13780 15360
rect 16948 15308 17000 15360
rect 17592 15376 17644 15428
rect 22560 15308 22612 15360
rect 23572 15308 23624 15360
rect 24860 15308 24912 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9772 15104 9824 15156
rect 12348 15104 12400 15156
rect 12808 15104 12860 15156
rect 3148 14900 3200 14952
rect 8116 14968 8168 15020
rect 11060 15036 11112 15088
rect 11520 15036 11572 15088
rect 9680 14968 9732 15020
rect 7748 14900 7800 14952
rect 11612 14968 11664 15020
rect 11980 14968 12032 15020
rect 13636 14900 13688 14952
rect 15384 15036 15436 15088
rect 16580 15104 16632 15156
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 19340 15104 19392 15156
rect 20352 15104 20404 15156
rect 20904 15104 20956 15156
rect 22100 15147 22152 15156
rect 22100 15113 22109 15147
rect 22109 15113 22143 15147
rect 22143 15113 22152 15147
rect 22100 15104 22152 15113
rect 25412 15104 25464 15156
rect 18788 15036 18840 15088
rect 9220 14832 9272 14884
rect 9588 14875 9640 14884
rect 9588 14841 9597 14875
rect 9597 14841 9631 14875
rect 9631 14841 9640 14875
rect 9588 14832 9640 14841
rect 12716 14875 12768 14884
rect 4988 14764 5040 14816
rect 8300 14807 8352 14816
rect 8300 14773 8309 14807
rect 8309 14773 8343 14807
rect 8343 14773 8352 14807
rect 8300 14764 8352 14773
rect 8392 14764 8444 14816
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 13452 14832 13504 14884
rect 14556 14968 14608 15020
rect 15476 15011 15528 15020
rect 12348 14764 12400 14816
rect 14280 14875 14332 14884
rect 14280 14841 14289 14875
rect 14289 14841 14323 14875
rect 14323 14841 14332 14875
rect 14280 14832 14332 14841
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 20720 15036 20772 15088
rect 20812 15011 20864 15020
rect 15384 14900 15436 14952
rect 16028 14900 16080 14952
rect 18420 14900 18472 14952
rect 19616 14900 19668 14952
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20904 14968 20956 15020
rect 24032 15011 24084 15020
rect 20996 14900 21048 14952
rect 21180 14900 21232 14952
rect 24032 14977 24041 15011
rect 24041 14977 24075 15011
rect 24075 14977 24084 15011
rect 24032 14968 24084 14977
rect 24860 14968 24912 15020
rect 25136 15011 25188 15020
rect 25136 14977 25145 15011
rect 25145 14977 25179 15011
rect 25179 14977 25188 15011
rect 25136 14968 25188 14977
rect 26056 14968 26108 15020
rect 37004 14968 37056 15020
rect 17408 14764 17460 14816
rect 23572 14807 23624 14816
rect 23572 14773 23581 14807
rect 23581 14773 23615 14807
rect 23615 14773 23624 14807
rect 23572 14764 23624 14773
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 24584 14764 24636 14816
rect 29368 14764 29420 14816
rect 33140 14807 33192 14816
rect 33140 14773 33149 14807
rect 33149 14773 33183 14807
rect 33183 14773 33192 14807
rect 33140 14764 33192 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4804 14603 4856 14612
rect 4804 14569 4813 14603
rect 4813 14569 4847 14603
rect 4847 14569 4856 14603
rect 4804 14560 4856 14569
rect 6368 14560 6420 14612
rect 8116 14560 8168 14612
rect 11244 14560 11296 14612
rect 6552 14492 6604 14544
rect 10600 14492 10652 14544
rect 10784 14492 10836 14544
rect 12256 14560 12308 14612
rect 12900 14560 12952 14612
rect 13360 14560 13412 14612
rect 15292 14560 15344 14612
rect 13820 14492 13872 14544
rect 16580 14560 16632 14612
rect 17040 14560 17092 14612
rect 17776 14560 17828 14612
rect 18328 14560 18380 14612
rect 20076 14560 20128 14612
rect 20168 14560 20220 14612
rect 24400 14560 24452 14612
rect 25872 14560 25924 14612
rect 12900 14424 12952 14476
rect 17132 14492 17184 14544
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2780 14356 2832 14408
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 8484 14356 8536 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 12072 14356 12124 14408
rect 12440 14356 12492 14408
rect 14464 14424 14516 14476
rect 15568 14424 15620 14476
rect 19616 14467 19668 14476
rect 9956 14288 10008 14340
rect 13176 14356 13228 14408
rect 14280 14356 14332 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 18420 14356 18472 14408
rect 22468 14492 22520 14544
rect 24216 14492 24268 14544
rect 24584 14467 24636 14476
rect 24584 14433 24593 14467
rect 24593 14433 24627 14467
rect 24627 14433 24636 14467
rect 24584 14424 24636 14433
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 21272 14356 21324 14408
rect 24492 14356 24544 14408
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 2596 14220 2648 14272
rect 9036 14220 9088 14272
rect 12072 14220 12124 14272
rect 12256 14220 12308 14272
rect 14004 14220 14056 14272
rect 14740 14220 14792 14272
rect 22192 14220 22244 14272
rect 26056 14220 26108 14272
rect 36452 14356 36504 14408
rect 37832 14288 37884 14340
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 9496 14016 9548 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 10692 14016 10744 14068
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 2780 13880 2832 13932
rect 5540 13948 5592 14000
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 7380 13880 7432 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 8208 13880 8260 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9956 13880 10008 13932
rect 10232 13880 10284 13932
rect 10416 13880 10468 13932
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 5632 13812 5684 13864
rect 7840 13812 7892 13864
rect 8300 13812 8352 13864
rect 10600 13880 10652 13932
rect 12440 13991 12492 14000
rect 12440 13957 12449 13991
rect 12449 13957 12483 13991
rect 12483 13957 12492 13991
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 12440 13948 12492 13957
rect 13728 13948 13780 14000
rect 16212 14016 16264 14068
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 19432 14016 19484 14068
rect 20904 14016 20956 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 15016 13948 15068 14000
rect 12900 13880 12952 13932
rect 14004 13880 14056 13932
rect 14280 13880 14332 13932
rect 21088 13948 21140 14000
rect 22008 13948 22060 14000
rect 24216 13991 24268 14000
rect 24216 13957 24225 13991
rect 24225 13957 24259 13991
rect 24259 13957 24268 13991
rect 24216 13948 24268 13957
rect 17592 13880 17644 13932
rect 18052 13880 18104 13932
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 20628 13880 20680 13932
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 26608 14016 26660 14068
rect 25504 13880 25556 13932
rect 9312 13744 9364 13796
rect 15384 13812 15436 13864
rect 15844 13812 15896 13864
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 17960 13812 18012 13864
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23112 13812 23164 13821
rect 24400 13812 24452 13864
rect 24768 13855 24820 13864
rect 24768 13821 24777 13855
rect 24777 13821 24811 13855
rect 24811 13821 24820 13855
rect 24768 13812 24820 13821
rect 10876 13744 10928 13796
rect 17132 13744 17184 13796
rect 23204 13744 23256 13796
rect 33140 13744 33192 13796
rect 2228 13676 2280 13728
rect 6368 13676 6420 13728
rect 10968 13676 11020 13728
rect 11612 13676 11664 13728
rect 12808 13676 12860 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 22652 13719 22704 13728
rect 22652 13685 22661 13719
rect 22661 13685 22695 13719
rect 22695 13685 22704 13719
rect 22652 13676 22704 13685
rect 23020 13676 23072 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7932 13472 7984 13524
rect 11336 13472 11388 13524
rect 11428 13515 11480 13524
rect 11428 13481 11437 13515
rect 11437 13481 11471 13515
rect 11471 13481 11480 13515
rect 11428 13472 11480 13481
rect 12348 13472 12400 13524
rect 5816 13404 5868 13456
rect 6828 13404 6880 13456
rect 4988 13336 5040 13388
rect 13728 13472 13780 13524
rect 9956 13336 10008 13388
rect 15844 13447 15896 13456
rect 15844 13413 15853 13447
rect 15853 13413 15887 13447
rect 15887 13413 15896 13447
rect 15844 13404 15896 13413
rect 16488 13379 16540 13388
rect 1400 13268 1452 13320
rect 2780 13268 2832 13320
rect 3608 13268 3660 13320
rect 3976 13268 4028 13320
rect 7380 13268 7432 13320
rect 7748 13268 7800 13320
rect 5080 13200 5132 13252
rect 9864 13268 9916 13320
rect 6644 13132 6696 13184
rect 8668 13200 8720 13252
rect 8024 13132 8076 13184
rect 9496 13132 9548 13184
rect 9956 13200 10008 13252
rect 10416 13268 10468 13320
rect 10876 13268 10928 13320
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 17408 13404 17460 13456
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 12900 13268 12952 13277
rect 15292 13311 15344 13320
rect 13176 13200 13228 13252
rect 13360 13200 13412 13252
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15016 13200 15068 13252
rect 17040 13268 17092 13320
rect 15936 13200 15988 13252
rect 20812 13472 20864 13524
rect 22468 13515 22520 13524
rect 22468 13481 22477 13515
rect 22477 13481 22511 13515
rect 22511 13481 22520 13515
rect 22468 13472 22520 13481
rect 22652 13472 22704 13524
rect 23296 13472 23348 13524
rect 24400 13472 24452 13524
rect 25136 13472 25188 13524
rect 25780 13472 25832 13524
rect 22836 13404 22888 13456
rect 23020 13336 23072 13388
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19064 13268 19116 13320
rect 19432 13268 19484 13320
rect 20168 13268 20220 13320
rect 23112 13268 23164 13320
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 24952 13379 25004 13388
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 23204 13268 23256 13277
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 26608 13311 26660 13320
rect 26608 13277 26617 13311
rect 26617 13277 26651 13311
rect 26651 13277 26660 13311
rect 26608 13268 26660 13277
rect 21456 13200 21508 13252
rect 24400 13200 24452 13252
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 10692 13132 10744 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 13268 13132 13320 13184
rect 16764 13132 16816 13184
rect 18052 13132 18104 13184
rect 20444 13175 20496 13184
rect 20444 13141 20453 13175
rect 20453 13141 20487 13175
rect 20487 13141 20496 13175
rect 20444 13132 20496 13141
rect 20812 13132 20864 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 8944 12928 8996 12980
rect 9128 12928 9180 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 2228 12792 2280 12844
rect 6460 12860 6512 12912
rect 6552 12860 6604 12912
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 6000 12835 6052 12844
rect 3976 12724 4028 12776
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 7104 12792 7156 12844
rect 9312 12860 9364 12912
rect 9404 12860 9456 12912
rect 9772 12860 9824 12912
rect 11888 12928 11940 12980
rect 12164 12928 12216 12980
rect 15476 12928 15528 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 17040 12928 17092 12980
rect 18788 12928 18840 12980
rect 20168 12971 20220 12980
rect 20168 12937 20177 12971
rect 20177 12937 20211 12971
rect 20211 12937 20220 12971
rect 20168 12928 20220 12937
rect 7932 12792 7984 12844
rect 8116 12792 8168 12844
rect 10968 12792 11020 12844
rect 12624 12792 12676 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14188 12792 14240 12844
rect 7656 12724 7708 12776
rect 8760 12724 8812 12776
rect 4804 12656 4856 12708
rect 14740 12724 14792 12776
rect 15844 12792 15896 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 18512 12792 18564 12844
rect 18880 12792 18932 12844
rect 21180 12928 21232 12980
rect 20444 12860 20496 12912
rect 22192 12903 22244 12912
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 22192 12869 22201 12903
rect 22201 12869 22235 12903
rect 22235 12869 22244 12903
rect 22192 12860 22244 12869
rect 36452 12928 36504 12980
rect 24492 12860 24544 12912
rect 24676 12792 24728 12844
rect 25504 12835 25556 12844
rect 25504 12801 25513 12835
rect 25513 12801 25547 12835
rect 25547 12801 25556 12835
rect 25504 12792 25556 12801
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 8024 12588 8076 12640
rect 8116 12588 8168 12640
rect 12440 12656 12492 12708
rect 12900 12656 12952 12708
rect 15384 12656 15436 12708
rect 17776 12724 17828 12776
rect 18236 12724 18288 12776
rect 21364 12724 21416 12776
rect 23388 12724 23440 12776
rect 23480 12724 23532 12776
rect 25228 12724 25280 12776
rect 18052 12699 18104 12708
rect 10600 12588 10652 12640
rect 13360 12588 13412 12640
rect 13728 12588 13780 12640
rect 14372 12588 14424 12640
rect 14740 12588 14792 12640
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 24032 12656 24084 12708
rect 29092 12792 29144 12844
rect 38016 12835 38068 12844
rect 38016 12801 38025 12835
rect 38025 12801 38059 12835
rect 38059 12801 38068 12835
rect 38016 12792 38068 12801
rect 17040 12588 17092 12640
rect 20628 12588 20680 12640
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21180 12588 21232 12597
rect 23204 12588 23256 12640
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5540 12384 5592 12436
rect 5908 12384 5960 12436
rect 8484 12384 8536 12436
rect 8576 12384 8628 12436
rect 10048 12384 10100 12436
rect 11428 12384 11480 12436
rect 12624 12384 12676 12436
rect 12808 12384 12860 12436
rect 13636 12384 13688 12436
rect 15936 12427 15988 12436
rect 15936 12393 15945 12427
rect 15945 12393 15979 12427
rect 15979 12393 15988 12427
rect 15936 12384 15988 12393
rect 17224 12384 17276 12436
rect 18236 12427 18288 12436
rect 18236 12393 18245 12427
rect 18245 12393 18279 12427
rect 18279 12393 18288 12427
rect 18236 12384 18288 12393
rect 20352 12384 20404 12436
rect 23480 12384 23532 12436
rect 8944 12316 8996 12368
rect 4620 12248 4672 12300
rect 6920 12248 6972 12300
rect 8300 12248 8352 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 10968 12248 11020 12300
rect 11336 12291 11388 12300
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 11612 12248 11664 12300
rect 11980 12248 12032 12300
rect 2780 12180 2832 12232
rect 3240 12180 3292 12232
rect 3792 12180 3844 12232
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 5908 12180 5960 12232
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 7196 12180 7248 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 8576 12223 8628 12232
rect 7748 12180 7800 12189
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 8668 12180 8720 12232
rect 9956 12180 10008 12232
rect 10876 12180 10928 12232
rect 11060 12180 11112 12232
rect 3056 12112 3108 12164
rect 13912 12248 13964 12300
rect 15384 12316 15436 12368
rect 14556 12248 14608 12300
rect 15016 12248 15068 12300
rect 16120 12248 16172 12300
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 24492 12316 24544 12368
rect 16672 12248 16724 12257
rect 13360 12180 13412 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 17132 12180 17184 12232
rect 18144 12180 18196 12232
rect 23296 12248 23348 12300
rect 23572 12248 23624 12300
rect 20260 12180 20312 12232
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 2412 12044 2464 12096
rect 3608 12044 3660 12096
rect 5540 12112 5592 12164
rect 4620 12044 4672 12096
rect 7012 12044 7064 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 8392 12087 8444 12096
rect 7104 12044 7156 12053
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 8484 12044 8536 12096
rect 10048 12044 10100 12096
rect 11980 12112 12032 12164
rect 12440 12155 12492 12164
rect 12440 12121 12449 12155
rect 12449 12121 12483 12155
rect 12483 12121 12492 12155
rect 12992 12155 13044 12164
rect 12440 12112 12492 12121
rect 12992 12121 13001 12155
rect 13001 12121 13035 12155
rect 13035 12121 13044 12155
rect 12992 12112 13044 12121
rect 13176 12112 13228 12164
rect 17224 12112 17276 12164
rect 17316 12112 17368 12164
rect 21180 12180 21232 12232
rect 24216 12180 24268 12232
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 38016 12384 38068 12436
rect 12256 12044 12308 12096
rect 12900 12044 12952 12096
rect 14280 12044 14332 12096
rect 15568 12044 15620 12096
rect 17040 12044 17092 12096
rect 17684 12044 17736 12096
rect 21916 12044 21968 12096
rect 22468 12044 22520 12096
rect 22744 12087 22796 12096
rect 22744 12053 22753 12087
rect 22753 12053 22787 12087
rect 22787 12053 22796 12087
rect 22744 12044 22796 12053
rect 22928 12112 22980 12164
rect 23756 12044 23808 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1584 11840 1636 11892
rect 5356 11772 5408 11824
rect 1492 11704 1544 11756
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 4620 11704 4672 11756
rect 8300 11840 8352 11892
rect 8484 11840 8536 11892
rect 8944 11840 8996 11892
rect 9404 11840 9456 11892
rect 11980 11840 12032 11892
rect 12072 11840 12124 11892
rect 12440 11840 12492 11892
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 18236 11840 18288 11892
rect 20260 11840 20312 11892
rect 21180 11840 21232 11892
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 22468 11840 22520 11892
rect 24952 11840 25004 11892
rect 25228 11883 25280 11892
rect 25228 11849 25237 11883
rect 25237 11849 25271 11883
rect 25271 11849 25280 11883
rect 25228 11840 25280 11849
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 5724 11636 5776 11688
rect 7196 11636 7248 11688
rect 7564 11704 7616 11756
rect 7472 11636 7524 11688
rect 1860 11500 1912 11552
rect 4160 11568 4212 11620
rect 8300 11636 8352 11688
rect 8668 11636 8720 11688
rect 7932 11568 7984 11620
rect 8208 11568 8260 11620
rect 9312 11704 9364 11756
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 11520 11704 11572 11756
rect 14188 11772 14240 11824
rect 14280 11815 14332 11824
rect 14280 11781 14289 11815
rect 14289 11781 14323 11815
rect 14323 11781 14332 11815
rect 14280 11772 14332 11781
rect 9404 11636 9456 11688
rect 9588 11636 9640 11688
rect 9772 11636 9824 11688
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 15844 11704 15896 11756
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 19892 11772 19944 11824
rect 18236 11704 18288 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18604 11704 18656 11756
rect 20168 11772 20220 11824
rect 21824 11772 21876 11824
rect 23020 11815 23072 11824
rect 23020 11781 23029 11815
rect 23029 11781 23063 11815
rect 23063 11781 23072 11815
rect 23020 11772 23072 11781
rect 25320 11772 25372 11824
rect 20628 11747 20680 11756
rect 20628 11713 20637 11747
rect 20637 11713 20671 11747
rect 20671 11713 20680 11747
rect 20628 11704 20680 11713
rect 26056 11747 26108 11756
rect 3884 11500 3936 11552
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 6184 11500 6236 11552
rect 7564 11500 7616 11552
rect 10416 11568 10468 11620
rect 12716 11636 12768 11688
rect 20444 11679 20496 11688
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 20444 11636 20496 11645
rect 16120 11568 16172 11620
rect 26056 11713 26065 11747
rect 26065 11713 26099 11747
rect 26099 11713 26108 11747
rect 26056 11704 26108 11713
rect 22928 11679 22980 11688
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 23664 11636 23716 11688
rect 23940 11636 23992 11688
rect 24860 11636 24912 11688
rect 25044 11636 25096 11688
rect 23848 11568 23900 11620
rect 24308 11568 24360 11620
rect 24676 11611 24728 11620
rect 24676 11577 24685 11611
rect 24685 11577 24719 11611
rect 24719 11577 24728 11611
rect 24676 11568 24728 11577
rect 9772 11500 9824 11552
rect 10508 11500 10560 11552
rect 11796 11500 11848 11552
rect 15476 11500 15528 11552
rect 15936 11500 15988 11552
rect 16396 11500 16448 11552
rect 18788 11500 18840 11552
rect 20352 11500 20404 11552
rect 20536 11500 20588 11552
rect 25872 11500 25924 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4068 11296 4120 11348
rect 8208 11296 8260 11348
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 9404 11296 9456 11348
rect 12072 11296 12124 11348
rect 3516 11228 3568 11280
rect 3976 11228 4028 11280
rect 5724 11271 5776 11280
rect 5724 11237 5733 11271
rect 5733 11237 5767 11271
rect 5767 11237 5776 11271
rect 5724 11228 5776 11237
rect 8300 11228 8352 11280
rect 10600 11271 10652 11280
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 3884 11160 3936 11212
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 9772 11160 9824 11212
rect 10324 11160 10376 11212
rect 10600 11237 10609 11271
rect 10609 11237 10643 11271
rect 10643 11237 10652 11271
rect 10600 11228 10652 11237
rect 11060 11228 11112 11280
rect 12440 11228 12492 11280
rect 11428 11160 11480 11212
rect 11888 11160 11940 11212
rect 6736 11092 6788 11144
rect 8392 11092 8444 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9680 11092 9732 11144
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 15752 11228 15804 11280
rect 16856 11296 16908 11348
rect 19432 11296 19484 11348
rect 20536 11296 20588 11348
rect 22192 11296 22244 11348
rect 16396 11228 16448 11280
rect 18972 11228 19024 11280
rect 20996 11228 21048 11280
rect 16212 11160 16264 11212
rect 16764 11160 16816 11212
rect 20444 11160 20496 11212
rect 14188 11092 14240 11144
rect 16396 11092 16448 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18236 11092 18288 11144
rect 4528 10956 4580 11008
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 7564 11024 7616 11076
rect 8668 10956 8720 11008
rect 10416 10956 10468 11008
rect 11796 11024 11848 11076
rect 13820 10956 13872 11008
rect 13912 10956 13964 11008
rect 14832 10956 14884 11008
rect 15844 11024 15896 11076
rect 17500 11024 17552 11076
rect 17868 11024 17920 11076
rect 19984 11092 20036 11144
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 22560 11228 22612 11280
rect 22468 11092 22520 11144
rect 24768 11296 24820 11348
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 29092 11296 29144 11348
rect 23848 11228 23900 11280
rect 25504 11228 25556 11280
rect 38200 11271 38252 11280
rect 38200 11237 38209 11271
rect 38209 11237 38243 11271
rect 38243 11237 38252 11271
rect 38200 11228 38252 11237
rect 25780 11160 25832 11212
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 25228 11135 25280 11144
rect 25228 11101 25237 11135
rect 25237 11101 25271 11135
rect 25271 11101 25280 11135
rect 25228 11092 25280 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 22100 11024 22152 11076
rect 22744 11024 22796 11076
rect 36084 11092 36136 11144
rect 28908 11024 28960 11076
rect 16120 10956 16172 11008
rect 16212 10956 16264 11008
rect 17960 10956 18012 11008
rect 18420 10956 18472 11008
rect 23296 10956 23348 11008
rect 23480 10999 23532 11008
rect 23480 10965 23489 10999
rect 23489 10965 23523 10999
rect 23523 10965 23532 10999
rect 23480 10956 23532 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3700 10752 3752 10804
rect 4160 10752 4212 10804
rect 5724 10684 5776 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 2504 10616 2556 10668
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 8392 10684 8444 10736
rect 8484 10684 8536 10736
rect 15844 10752 15896 10804
rect 16120 10752 16172 10804
rect 12348 10684 12400 10736
rect 12808 10684 12860 10736
rect 16856 10684 16908 10736
rect 17316 10684 17368 10736
rect 19892 10684 19944 10736
rect 20536 10752 20588 10804
rect 23756 10795 23808 10804
rect 23756 10761 23765 10795
rect 23765 10761 23799 10795
rect 23799 10761 23808 10795
rect 23756 10752 23808 10761
rect 25044 10795 25096 10804
rect 25044 10761 25053 10795
rect 25053 10761 25087 10795
rect 25087 10761 25096 10795
rect 25044 10752 25096 10761
rect 20628 10684 20680 10736
rect 22100 10684 22152 10736
rect 10140 10616 10192 10668
rect 10692 10616 10744 10668
rect 10784 10616 10836 10668
rect 2964 10548 3016 10600
rect 3424 10548 3476 10600
rect 7748 10548 7800 10600
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 10600 10548 10652 10600
rect 11060 10548 11112 10600
rect 20352 10659 20404 10668
rect 8116 10480 8168 10532
rect 9496 10480 9548 10532
rect 11888 10480 11940 10532
rect 1676 10412 1728 10464
rect 7472 10412 7524 10464
rect 9128 10412 9180 10464
rect 10048 10412 10100 10464
rect 10692 10412 10744 10464
rect 10876 10412 10928 10464
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 15476 10548 15528 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17224 10548 17276 10600
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 19524 10591 19576 10600
rect 13820 10480 13872 10532
rect 13912 10412 13964 10464
rect 15568 10480 15620 10532
rect 16212 10480 16264 10532
rect 19524 10557 19533 10591
rect 19533 10557 19567 10591
rect 19567 10557 19576 10591
rect 19524 10548 19576 10557
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 23388 10616 23440 10668
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24032 10616 24084 10668
rect 24124 10548 24176 10600
rect 18880 10480 18932 10532
rect 23388 10480 23440 10532
rect 25320 10548 25372 10600
rect 33692 10480 33744 10532
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 18512 10412 18564 10464
rect 20168 10412 20220 10464
rect 20996 10412 21048 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4712 10208 4764 10260
rect 5264 10208 5316 10260
rect 6920 10208 6972 10260
rect 8116 10208 8168 10260
rect 10876 10208 10928 10260
rect 4068 10140 4120 10192
rect 2964 10072 3016 10124
rect 6000 10072 6052 10124
rect 8668 10140 8720 10192
rect 10416 10140 10468 10192
rect 22192 10208 22244 10260
rect 23020 10208 23072 10260
rect 23204 10208 23256 10260
rect 24216 10208 24268 10260
rect 25320 10251 25372 10260
rect 25320 10217 25329 10251
rect 25329 10217 25363 10251
rect 25363 10217 25372 10251
rect 25320 10208 25372 10217
rect 36084 10208 36136 10260
rect 13176 10140 13228 10192
rect 13728 10140 13780 10192
rect 16856 10140 16908 10192
rect 23112 10140 23164 10192
rect 23296 10140 23348 10192
rect 8208 10072 8260 10124
rect 11060 10072 11112 10124
rect 11888 10115 11940 10124
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 3976 10004 4028 10056
rect 5632 10004 5684 10056
rect 8300 10004 8352 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 10692 10004 10744 10056
rect 6092 9868 6144 9920
rect 6276 9868 6328 9920
rect 6736 9936 6788 9988
rect 7288 9936 7340 9988
rect 8116 9936 8168 9988
rect 10968 9936 11020 9988
rect 17224 10072 17276 10124
rect 17868 10072 17920 10124
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 18880 10072 18932 10124
rect 19524 10115 19576 10124
rect 19524 10081 19533 10115
rect 19533 10081 19567 10115
rect 19567 10081 19576 10115
rect 19524 10072 19576 10081
rect 19616 10072 19668 10124
rect 20996 10115 21048 10124
rect 20996 10081 21005 10115
rect 21005 10081 21039 10115
rect 21039 10081 21048 10115
rect 20996 10072 21048 10081
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 16488 10004 16540 10056
rect 16672 10004 16724 10056
rect 17040 10004 17092 10056
rect 20812 10047 20864 10056
rect 14832 9936 14884 9988
rect 14464 9868 14516 9920
rect 17316 9936 17368 9988
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 22192 10004 22244 10056
rect 22376 10004 22428 10056
rect 23480 10004 23532 10056
rect 16212 9868 16264 9920
rect 17592 9868 17644 9920
rect 17868 9868 17920 9920
rect 19432 9868 19484 9920
rect 19892 9936 19944 9988
rect 22836 9936 22888 9988
rect 23112 9936 23164 9988
rect 24032 10004 24084 10056
rect 26056 10004 26108 10056
rect 28908 10004 28960 10056
rect 35072 10047 35124 10056
rect 35072 10013 35081 10047
rect 35081 10013 35115 10047
rect 35115 10013 35124 10047
rect 35072 10004 35124 10013
rect 21456 9911 21508 9920
rect 21456 9877 21465 9911
rect 21465 9877 21499 9911
rect 21499 9877 21508 9911
rect 21456 9868 21508 9877
rect 23940 9868 23992 9920
rect 34796 9868 34848 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4620 9664 4672 9716
rect 4896 9664 4948 9716
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 2780 9528 2832 9580
rect 2872 9460 2924 9512
rect 3424 9392 3476 9444
rect 3240 9324 3292 9376
rect 3608 9324 3660 9376
rect 4068 9596 4120 9648
rect 8484 9664 8536 9716
rect 3976 9460 4028 9512
rect 5724 9460 5776 9512
rect 7656 9596 7708 9648
rect 16856 9664 16908 9716
rect 17776 9664 17828 9716
rect 18420 9664 18472 9716
rect 12348 9596 12400 9648
rect 13820 9596 13872 9648
rect 14004 9639 14056 9648
rect 14004 9605 14013 9639
rect 14013 9605 14047 9639
rect 14047 9605 14056 9639
rect 14004 9596 14056 9605
rect 14832 9596 14884 9648
rect 16120 9596 16172 9648
rect 19248 9639 19300 9648
rect 8208 9528 8260 9580
rect 11244 9528 11296 9580
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6736 9460 6788 9512
rect 5908 9392 5960 9444
rect 6828 9392 6880 9444
rect 11060 9460 11112 9512
rect 14004 9460 14056 9512
rect 14280 9460 14332 9512
rect 11152 9392 11204 9444
rect 11704 9392 11756 9444
rect 13820 9392 13872 9444
rect 15752 9460 15804 9512
rect 16028 9460 16080 9512
rect 16580 9460 16632 9512
rect 19248 9605 19257 9639
rect 19257 9605 19291 9639
rect 19291 9605 19300 9639
rect 19248 9596 19300 9605
rect 20076 9664 20128 9716
rect 20444 9664 20496 9716
rect 20812 9664 20864 9716
rect 22192 9596 22244 9648
rect 22468 9639 22520 9648
rect 22468 9605 22477 9639
rect 22477 9605 22511 9639
rect 22511 9605 22520 9639
rect 22468 9596 22520 9605
rect 23204 9596 23256 9648
rect 20076 9528 20128 9580
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 25504 9528 25556 9580
rect 35072 9596 35124 9648
rect 23296 9503 23348 9512
rect 23296 9469 23305 9503
rect 23305 9469 23339 9503
rect 23339 9469 23348 9503
rect 23296 9460 23348 9469
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 23480 9460 23532 9469
rect 24400 9503 24452 9512
rect 24400 9469 24409 9503
rect 24409 9469 24443 9503
rect 24443 9469 24452 9503
rect 24400 9460 24452 9469
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 10876 9324 10928 9376
rect 12900 9324 12952 9376
rect 13360 9324 13412 9376
rect 17960 9324 18012 9376
rect 18236 9324 18288 9376
rect 23940 9324 23992 9376
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 30196 9324 30248 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3424 9120 3476 9172
rect 3608 9052 3660 9104
rect 6552 9052 6604 9104
rect 9680 9120 9732 9172
rect 2872 8984 2924 9036
rect 3424 8984 3476 9036
rect 2780 8916 2832 8968
rect 1308 8848 1360 8900
rect 3056 8848 3108 8900
rect 3608 8916 3660 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 2412 8780 2464 8832
rect 2872 8780 2924 8832
rect 4160 8780 4212 8832
rect 5264 8780 5316 8832
rect 10968 8984 11020 9036
rect 11060 8984 11112 9036
rect 11888 9120 11940 9172
rect 12716 9120 12768 9172
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 16396 9120 16448 9172
rect 12440 9052 12492 9104
rect 13268 9052 13320 9104
rect 14096 9052 14148 9104
rect 14372 9052 14424 9104
rect 18604 9120 18656 9172
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 20352 9120 20404 9172
rect 21640 9052 21692 9104
rect 22100 9120 22152 9172
rect 23480 9120 23532 9172
rect 5724 8916 5776 8968
rect 6552 8916 6604 8968
rect 6736 8916 6788 8968
rect 8208 8916 8260 8968
rect 9404 8916 9456 8968
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9772 8916 9824 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 13176 8916 13228 8968
rect 13544 8916 13596 8968
rect 5816 8780 5868 8832
rect 7380 8780 7432 8832
rect 8392 8780 8444 8832
rect 8760 8848 8812 8900
rect 11152 8848 11204 8900
rect 9312 8780 9364 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 13176 8780 13228 8832
rect 14280 8916 14332 8968
rect 16396 8916 16448 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 19064 8984 19116 9036
rect 17500 8848 17552 8900
rect 20076 8916 20128 8968
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 22468 8916 22520 8968
rect 22376 8848 22428 8900
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 24768 9052 24820 9104
rect 22836 8916 22888 8925
rect 24492 8916 24544 8968
rect 24676 8916 24728 8968
rect 34796 8916 34848 8968
rect 17224 8823 17276 8832
rect 17224 8789 17233 8823
rect 17233 8789 17267 8823
rect 17267 8789 17276 8823
rect 17224 8780 17276 8789
rect 17316 8780 17368 8832
rect 23480 8780 23532 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4068 8576 4120 8628
rect 4160 8576 4212 8628
rect 6460 8576 6512 8628
rect 7104 8576 7156 8628
rect 4988 8508 5040 8560
rect 5264 8508 5316 8560
rect 7656 8508 7708 8560
rect 9404 8576 9456 8628
rect 12440 8576 12492 8628
rect 17040 8576 17092 8628
rect 19248 8619 19300 8628
rect 2872 8440 2924 8492
rect 2964 8415 3016 8424
rect 1584 8304 1636 8356
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 2872 8304 2924 8356
rect 3700 8372 3752 8424
rect 5724 8440 5776 8492
rect 5448 8372 5500 8424
rect 7012 8440 7064 8492
rect 4528 8304 4580 8356
rect 6736 8372 6788 8424
rect 8116 8372 8168 8424
rect 3884 8236 3936 8288
rect 3976 8236 4028 8288
rect 5632 8304 5684 8356
rect 10968 8372 11020 8424
rect 9404 8304 9456 8356
rect 11152 8304 11204 8356
rect 12164 8440 12216 8492
rect 12532 8508 12584 8560
rect 12992 8508 13044 8560
rect 13360 8551 13412 8560
rect 13360 8517 13369 8551
rect 13369 8517 13403 8551
rect 13403 8517 13412 8551
rect 13360 8508 13412 8517
rect 14372 8508 14424 8560
rect 13728 8372 13780 8424
rect 5448 8236 5500 8288
rect 13728 8236 13780 8288
rect 14464 8372 14516 8424
rect 15568 8440 15620 8492
rect 17316 8440 17368 8492
rect 15476 8372 15528 8424
rect 16396 8372 16448 8424
rect 18236 8551 18288 8560
rect 18236 8517 18245 8551
rect 18245 8517 18279 8551
rect 18279 8517 18288 8551
rect 18236 8508 18288 8517
rect 18420 8508 18472 8560
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 23204 8619 23256 8628
rect 23204 8585 23213 8619
rect 23213 8585 23247 8619
rect 23247 8585 23256 8619
rect 23204 8576 23256 8585
rect 23296 8576 23348 8628
rect 24584 8576 24636 8628
rect 24952 8576 25004 8628
rect 33692 8619 33744 8628
rect 33692 8585 33701 8619
rect 33701 8585 33735 8619
rect 33735 8585 33744 8619
rect 33692 8576 33744 8585
rect 21824 8508 21876 8560
rect 19156 8440 19208 8492
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 24308 8440 24360 8492
rect 25504 8508 25556 8560
rect 29736 8440 29788 8492
rect 34704 8440 34756 8492
rect 19340 8372 19392 8424
rect 17316 8347 17368 8356
rect 14280 8236 14332 8288
rect 15476 8236 15528 8288
rect 16212 8236 16264 8288
rect 17040 8236 17092 8288
rect 17316 8313 17325 8347
rect 17325 8313 17359 8347
rect 17359 8313 17368 8347
rect 17316 8304 17368 8313
rect 17500 8304 17552 8356
rect 22560 8415 22612 8424
rect 22560 8381 22569 8415
rect 22569 8381 22603 8415
rect 22603 8381 22612 8415
rect 22560 8372 22612 8381
rect 23848 8372 23900 8424
rect 17960 8236 18012 8288
rect 18788 8236 18840 8288
rect 19156 8236 19208 8288
rect 20812 8236 20864 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2688 8032 2740 8084
rect 5264 8032 5316 8084
rect 10232 8032 10284 8084
rect 12900 7964 12952 8016
rect 16304 8032 16356 8084
rect 6736 7896 6788 7948
rect 6828 7896 6880 7948
rect 16764 7964 16816 8016
rect 15016 7896 15068 7948
rect 20536 8032 20588 8084
rect 21456 8032 21508 8084
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 23848 8075 23900 8084
rect 23848 8041 23857 8075
rect 23857 8041 23891 8075
rect 23891 8041 23900 8075
rect 23848 8032 23900 8041
rect 34704 8032 34756 8084
rect 17040 7964 17092 8016
rect 9864 7828 9916 7880
rect 10232 7828 10284 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 12532 7828 12584 7880
rect 14280 7871 14332 7880
rect 1676 7803 1728 7812
rect 1676 7769 1685 7803
rect 1685 7769 1719 7803
rect 1719 7769 1728 7803
rect 1676 7760 1728 7769
rect 2964 7760 3016 7812
rect 3608 7760 3660 7812
rect 4620 7760 4672 7812
rect 5540 7760 5592 7812
rect 9404 7692 9456 7744
rect 11704 7760 11756 7812
rect 12624 7760 12676 7812
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 17408 7896 17460 7948
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 18604 7964 18656 8016
rect 19248 7964 19300 8016
rect 19708 7964 19760 8016
rect 19432 7908 19484 7960
rect 20812 7939 20864 7948
rect 20812 7905 20821 7939
rect 20821 7905 20855 7939
rect 20855 7905 20864 7939
rect 20812 7896 20864 7905
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 19340 7828 19392 7880
rect 14648 7760 14700 7812
rect 17040 7803 17092 7812
rect 17040 7769 17049 7803
rect 17049 7769 17083 7803
rect 17083 7769 17092 7803
rect 17592 7803 17644 7812
rect 17040 7760 17092 7769
rect 17592 7769 17601 7803
rect 17601 7769 17635 7803
rect 17635 7769 17644 7803
rect 17592 7760 17644 7769
rect 12164 7692 12216 7744
rect 13268 7692 13320 7744
rect 16028 7692 16080 7744
rect 16120 7692 16172 7744
rect 18144 7692 18196 7744
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 19064 7760 19116 7812
rect 19340 7692 19392 7744
rect 19616 7803 19668 7812
rect 19616 7769 19625 7803
rect 19625 7769 19659 7803
rect 19659 7769 19668 7803
rect 19616 7760 19668 7769
rect 20444 7692 20496 7744
rect 20536 7692 20588 7744
rect 21916 7828 21968 7880
rect 22376 7871 22428 7880
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 24676 7964 24728 8016
rect 25412 7828 25464 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 21364 7760 21416 7812
rect 24492 7692 24544 7744
rect 24676 7735 24728 7744
rect 24676 7701 24685 7735
rect 24685 7701 24719 7735
rect 24719 7701 24728 7735
rect 24676 7692 24728 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2688 7488 2740 7540
rect 7196 7488 7248 7540
rect 1400 7420 1452 7472
rect 1860 7420 1912 7472
rect 3700 7420 3752 7472
rect 7840 7488 7892 7540
rect 12624 7488 12676 7540
rect 12716 7488 12768 7540
rect 9404 7463 9456 7472
rect 9404 7429 9413 7463
rect 9413 7429 9447 7463
rect 9447 7429 9456 7463
rect 9404 7420 9456 7429
rect 11060 7420 11112 7472
rect 2780 7352 2832 7404
rect 2964 7352 3016 7404
rect 3424 7352 3476 7404
rect 3608 7352 3660 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 10876 7352 10928 7404
rect 5172 7284 5224 7336
rect 5908 7327 5960 7336
rect 5908 7293 5917 7327
rect 5917 7293 5951 7327
rect 5951 7293 5960 7327
rect 5908 7284 5960 7293
rect 7472 7284 7524 7336
rect 9680 7284 9732 7336
rect 11704 7284 11756 7336
rect 4068 7216 4120 7268
rect 12532 7420 12584 7472
rect 12900 7352 12952 7404
rect 14004 7463 14056 7472
rect 14004 7429 14013 7463
rect 14013 7429 14047 7463
rect 14047 7429 14056 7463
rect 14004 7420 14056 7429
rect 16488 7420 16540 7472
rect 18236 7488 18288 7540
rect 20444 7488 20496 7540
rect 22284 7488 22336 7540
rect 24400 7488 24452 7540
rect 18604 7420 18656 7472
rect 18696 7420 18748 7472
rect 19616 7420 19668 7472
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 16580 7352 16632 7404
rect 18144 7352 18196 7404
rect 21456 7420 21508 7472
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 18328 7284 18380 7336
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 21180 7352 21232 7404
rect 22928 7395 22980 7404
rect 20904 7284 20956 7336
rect 21824 7284 21876 7336
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 23572 7284 23624 7336
rect 24676 7284 24728 7336
rect 35808 7352 35860 7404
rect 31944 7284 31996 7336
rect 12532 7216 12584 7268
rect 5448 7148 5500 7200
rect 6000 7148 6052 7200
rect 7564 7148 7616 7200
rect 10508 7148 10560 7200
rect 13452 7148 13504 7200
rect 19432 7216 19484 7268
rect 19616 7259 19668 7268
rect 19616 7225 19625 7259
rect 19625 7225 19659 7259
rect 19659 7225 19668 7259
rect 19616 7216 19668 7225
rect 15752 7148 15804 7200
rect 16488 7148 16540 7200
rect 20444 7148 20496 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 20996 7216 21048 7268
rect 26516 7216 26568 7268
rect 23112 7148 23164 7200
rect 23940 7148 23992 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3700 6944 3752 6996
rect 5908 6944 5960 6996
rect 10140 6944 10192 6996
rect 10324 6944 10376 6996
rect 12256 6944 12308 6996
rect 12900 6944 12952 6996
rect 13728 6944 13780 6996
rect 14280 6944 14332 6996
rect 5264 6876 5316 6928
rect 6092 6876 6144 6928
rect 12440 6876 12492 6928
rect 15108 6876 15160 6928
rect 17224 6944 17276 6996
rect 17408 6944 17460 6996
rect 22652 6944 22704 6996
rect 24492 6944 24544 6996
rect 1584 6808 1636 6860
rect 1768 6808 1820 6860
rect 3240 6808 3292 6860
rect 5724 6851 5776 6860
rect 1584 6672 1636 6724
rect 2688 6604 2740 6656
rect 4896 6672 4948 6724
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 6368 6808 6420 6860
rect 7472 6808 7524 6860
rect 6276 6740 6328 6792
rect 9220 6808 9272 6860
rect 9956 6808 10008 6860
rect 11060 6808 11112 6860
rect 11152 6808 11204 6860
rect 12348 6851 12400 6860
rect 9404 6740 9456 6792
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 14556 6808 14608 6860
rect 14648 6808 14700 6860
rect 16488 6876 16540 6928
rect 16856 6876 16908 6928
rect 17592 6876 17644 6928
rect 20996 6876 21048 6928
rect 17316 6808 17368 6860
rect 17684 6851 17736 6860
rect 17684 6817 17693 6851
rect 17693 6817 17727 6851
rect 17727 6817 17736 6851
rect 17684 6808 17736 6817
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 19432 6851 19484 6860
rect 19432 6817 19441 6851
rect 19441 6817 19475 6851
rect 19475 6817 19484 6851
rect 19432 6808 19484 6817
rect 19524 6808 19576 6860
rect 20260 6808 20312 6860
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 13728 6783 13780 6792
rect 12992 6740 13044 6749
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14004 6740 14056 6792
rect 16212 6740 16264 6792
rect 19892 6740 19944 6792
rect 22468 6808 22520 6860
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 21824 6740 21876 6792
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 23388 6740 23440 6792
rect 5264 6604 5316 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7012 6672 7064 6724
rect 7196 6672 7248 6724
rect 8392 6672 8444 6724
rect 9496 6604 9548 6656
rect 9864 6604 9916 6656
rect 11888 6672 11940 6724
rect 14924 6672 14976 6724
rect 15844 6672 15896 6724
rect 16580 6672 16632 6724
rect 10876 6604 10928 6656
rect 12256 6604 12308 6656
rect 12716 6604 12768 6656
rect 16120 6604 16172 6656
rect 18144 6604 18196 6656
rect 20168 6672 20220 6724
rect 18972 6604 19024 6656
rect 20260 6604 20312 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 20904 6604 20956 6656
rect 21364 6604 21416 6656
rect 21916 6604 21968 6656
rect 23204 6647 23256 6656
rect 23204 6613 23213 6647
rect 23213 6613 23247 6647
rect 23247 6613 23256 6647
rect 23204 6604 23256 6613
rect 23296 6604 23348 6656
rect 24032 6740 24084 6792
rect 30288 6740 30340 6792
rect 36360 6740 36412 6792
rect 38016 6604 38068 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1400 6400 1452 6452
rect 1676 6400 1728 6452
rect 2872 6400 2924 6452
rect 4712 6400 4764 6452
rect 4896 6400 4948 6452
rect 3608 6332 3660 6384
rect 1768 6264 1820 6316
rect 1492 6196 1544 6248
rect 2688 6196 2740 6248
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 3608 6196 3660 6248
rect 5264 6332 5316 6384
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 5908 6264 5960 6316
rect 7012 6400 7064 6452
rect 6736 6332 6788 6384
rect 9864 6400 9916 6452
rect 11796 6400 11848 6452
rect 11980 6400 12032 6452
rect 13728 6400 13780 6452
rect 14188 6400 14240 6452
rect 14556 6400 14608 6452
rect 9220 6375 9272 6384
rect 9220 6341 9229 6375
rect 9229 6341 9263 6375
rect 9263 6341 9272 6375
rect 9220 6332 9272 6341
rect 9772 6332 9824 6384
rect 10508 6332 10560 6384
rect 12900 6332 12952 6384
rect 13820 6332 13872 6384
rect 15752 6375 15804 6384
rect 15752 6341 15761 6375
rect 15761 6341 15795 6375
rect 15795 6341 15804 6375
rect 15752 6332 15804 6341
rect 15936 6332 15988 6384
rect 20260 6400 20312 6452
rect 21272 6400 21324 6452
rect 22560 6400 22612 6452
rect 19432 6332 19484 6384
rect 19984 6332 20036 6384
rect 11796 6264 11848 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 16488 6264 16540 6316
rect 16672 6264 16724 6316
rect 19892 6264 19944 6316
rect 24584 6332 24636 6384
rect 20628 6307 20680 6316
rect 20628 6273 20637 6307
rect 20637 6273 20671 6307
rect 20671 6273 20680 6307
rect 20628 6264 20680 6273
rect 21180 6264 21232 6316
rect 21456 6264 21508 6316
rect 23480 6264 23532 6316
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 6368 6196 6420 6248
rect 8668 6196 8720 6248
rect 9220 6196 9272 6248
rect 6552 6128 6604 6180
rect 10692 6196 10744 6248
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 13360 6196 13412 6248
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 16120 6196 16172 6248
rect 2596 6060 2648 6112
rect 4712 6060 4764 6112
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 18512 6196 18564 6248
rect 21548 6196 21600 6248
rect 24768 6196 24820 6248
rect 37464 6239 37516 6248
rect 37464 6205 37473 6239
rect 37473 6205 37507 6239
rect 37507 6205 37516 6239
rect 37464 6196 37516 6205
rect 9864 6060 9916 6112
rect 10784 6060 10836 6112
rect 11980 6060 12032 6112
rect 12440 6060 12492 6112
rect 16764 6060 16816 6112
rect 20904 6128 20956 6180
rect 21272 6060 21324 6112
rect 24676 6060 24728 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4620 5856 4672 5908
rect 2596 5720 2648 5772
rect 4988 5720 5040 5772
rect 6000 5788 6052 5840
rect 7840 5856 7892 5908
rect 10508 5856 10560 5908
rect 11428 5856 11480 5908
rect 10416 5788 10468 5840
rect 12716 5856 12768 5908
rect 15568 5856 15620 5908
rect 16488 5856 16540 5908
rect 7012 5720 7064 5772
rect 7196 5720 7248 5772
rect 1492 5652 1544 5704
rect 7932 5720 7984 5772
rect 9496 5720 9548 5772
rect 14096 5788 14148 5840
rect 15844 5788 15896 5840
rect 18420 5856 18472 5908
rect 19156 5856 19208 5908
rect 20352 5856 20404 5908
rect 12532 5720 12584 5772
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 16488 5763 16540 5772
rect 14280 5720 14332 5729
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 19892 5788 19944 5840
rect 22560 5856 22612 5908
rect 23756 5856 23808 5908
rect 18052 5720 18104 5772
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8944 5652 8996 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 10876 5652 10928 5704
rect 2320 5584 2372 5636
rect 6368 5584 6420 5636
rect 6644 5516 6696 5568
rect 8208 5584 8260 5636
rect 9496 5584 9548 5636
rect 9864 5584 9916 5636
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 8668 5516 8720 5568
rect 11796 5652 11848 5704
rect 11980 5652 12032 5704
rect 12992 5652 13044 5704
rect 13544 5652 13596 5704
rect 21364 5720 21416 5772
rect 19340 5652 19392 5704
rect 19984 5652 20036 5704
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 21180 5695 21232 5704
rect 20536 5652 20588 5661
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 12716 5516 12768 5568
rect 12900 5516 12952 5568
rect 13452 5516 13504 5568
rect 13912 5584 13964 5636
rect 15936 5516 15988 5568
rect 16304 5584 16356 5636
rect 20812 5584 20864 5636
rect 20904 5584 20956 5636
rect 23020 5652 23072 5704
rect 23480 5652 23532 5704
rect 30196 5652 30248 5704
rect 20352 5516 20404 5568
rect 20720 5516 20772 5568
rect 21088 5516 21140 5568
rect 22008 5516 22060 5568
rect 33048 5516 33100 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 5724 5312 5776 5364
rect 7288 5312 7340 5364
rect 7748 5312 7800 5364
rect 8208 5312 8260 5364
rect 9036 5355 9088 5364
rect 9036 5321 9045 5355
rect 9045 5321 9079 5355
rect 9079 5321 9088 5355
rect 9036 5312 9088 5321
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 9864 5312 9916 5364
rect 10692 5312 10744 5364
rect 10968 5312 11020 5364
rect 12164 5312 12216 5364
rect 7196 5244 7248 5296
rect 7840 5244 7892 5296
rect 1676 5176 1728 5228
rect 2228 5176 2280 5228
rect 2688 5176 2740 5228
rect 4988 5176 5040 5228
rect 4620 5108 4672 5160
rect 6828 5176 6880 5228
rect 7012 5176 7064 5228
rect 5724 5108 5776 5160
rect 11152 5244 11204 5296
rect 12808 5287 12860 5296
rect 12808 5253 12817 5287
rect 12817 5253 12851 5287
rect 12851 5253 12860 5287
rect 12808 5244 12860 5253
rect 12992 5244 13044 5296
rect 14004 5312 14056 5364
rect 15108 5355 15160 5364
rect 15108 5321 15117 5355
rect 15117 5321 15151 5355
rect 15151 5321 15160 5355
rect 15108 5312 15160 5321
rect 17040 5312 17092 5364
rect 14096 5244 14148 5296
rect 18880 5312 18932 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19432 5312 19484 5364
rect 20444 5312 20496 5364
rect 20720 5312 20772 5364
rect 24124 5312 24176 5364
rect 10140 5176 10192 5228
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10416 5176 10468 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11520 5176 11572 5228
rect 12164 5176 12216 5228
rect 12900 5176 12952 5228
rect 15016 5176 15068 5228
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 2044 5040 2096 5092
rect 9496 5108 9548 5160
rect 12440 5108 12492 5160
rect 12532 5108 12584 5160
rect 21916 5244 21968 5296
rect 22192 5244 22244 5296
rect 24492 5244 24544 5296
rect 19708 5219 19760 5228
rect 16856 5151 16908 5160
rect 20 4972 72 5024
rect 2780 4972 2832 5024
rect 6368 4972 6420 5024
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 10324 4972 10376 5024
rect 14832 5040 14884 5092
rect 18604 5108 18656 5160
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 20536 5176 20588 5228
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 22008 5217 22060 5228
rect 22008 5183 22017 5217
rect 22017 5183 22051 5217
rect 22051 5183 22060 5217
rect 22008 5176 22060 5183
rect 23756 5176 23808 5228
rect 26516 5219 26568 5228
rect 21824 5108 21876 5160
rect 21916 5108 21968 5160
rect 23480 5108 23532 5160
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 38016 5219 38068 5228
rect 38016 5185 38025 5219
rect 38025 5185 38059 5219
rect 38059 5185 38068 5219
rect 38016 5176 38068 5185
rect 12624 4972 12676 5024
rect 16488 4972 16540 5024
rect 16672 4972 16724 5024
rect 23940 5040 23992 5092
rect 19248 4972 19300 5024
rect 19708 4972 19760 5024
rect 21088 5015 21140 5024
rect 21088 4981 21097 5015
rect 21097 4981 21131 5015
rect 21131 4981 21140 5015
rect 21088 4972 21140 4981
rect 21640 4972 21692 5024
rect 21916 4972 21968 5024
rect 22100 5015 22152 5024
rect 22100 4981 22109 5015
rect 22109 4981 22143 5015
rect 22143 4981 22152 5015
rect 22744 5015 22796 5024
rect 22100 4972 22152 4981
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 32312 4972 32364 5024
rect 38016 4972 38068 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 6092 4768 6144 4820
rect 3056 4700 3108 4752
rect 3148 4700 3200 4752
rect 7932 4700 7984 4752
rect 9312 4768 9364 4820
rect 13268 4811 13320 4820
rect 13268 4777 13277 4811
rect 13277 4777 13311 4811
rect 13311 4777 13320 4811
rect 13268 4768 13320 4777
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 16396 4768 16448 4820
rect 18052 4768 18104 4820
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 18604 4768 18656 4820
rect 11428 4700 11480 4752
rect 20628 4700 20680 4752
rect 21456 4768 21508 4820
rect 23388 4768 23440 4820
rect 24768 4768 24820 4820
rect 31944 4811 31996 4820
rect 31944 4777 31953 4811
rect 31953 4777 31987 4811
rect 31987 4777 31996 4811
rect 31944 4768 31996 4777
rect 35808 4768 35860 4820
rect 3240 4632 3292 4684
rect 3424 4632 3476 4684
rect 6460 4632 6512 4684
rect 7012 4632 7064 4684
rect 9128 4632 9180 4684
rect 10140 4632 10192 4684
rect 11796 4632 11848 4684
rect 12164 4632 12216 4684
rect 1492 4564 1544 4616
rect 4620 4607 4672 4616
rect 3516 4496 3568 4548
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 7840 4564 7892 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 11336 4564 11388 4616
rect 14004 4632 14056 4684
rect 14280 4675 14332 4684
rect 14280 4641 14289 4675
rect 14289 4641 14323 4675
rect 14323 4641 14332 4675
rect 14280 4632 14332 4641
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 16672 4675 16724 4684
rect 16672 4641 16681 4675
rect 16681 4641 16715 4675
rect 16715 4641 16724 4675
rect 16672 4632 16724 4641
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 23848 4700 23900 4752
rect 27620 4700 27672 4752
rect 14188 4564 14240 4616
rect 18880 4564 18932 4616
rect 20168 4564 20220 4616
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22008 4564 22060 4616
rect 23940 4607 23992 4616
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 4620 4428 4672 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 6368 4539 6420 4548
rect 6368 4505 6377 4539
rect 6377 4505 6411 4539
rect 6411 4505 6420 4539
rect 6368 4496 6420 4505
rect 6920 4496 6972 4548
rect 8208 4428 8260 4480
rect 8668 4428 8720 4480
rect 9588 4539 9640 4548
rect 9588 4505 9597 4539
rect 9597 4505 9631 4539
rect 9631 4505 9640 4539
rect 9588 4496 9640 4505
rect 10876 4496 10928 4548
rect 10324 4428 10376 4480
rect 11520 4496 11572 4548
rect 12256 4496 12308 4548
rect 11336 4428 11388 4480
rect 13912 4428 13964 4480
rect 14832 4428 14884 4480
rect 15476 4428 15528 4480
rect 16764 4539 16816 4548
rect 16764 4505 16773 4539
rect 16773 4505 16807 4539
rect 16807 4505 16816 4539
rect 16764 4496 16816 4505
rect 17960 4496 18012 4548
rect 33876 4564 33928 4616
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 33600 4496 33652 4548
rect 19156 4428 19208 4480
rect 20076 4471 20128 4480
rect 20076 4437 20085 4471
rect 20085 4437 20119 4471
rect 20119 4437 20128 4471
rect 20076 4428 20128 4437
rect 21916 4471 21968 4480
rect 21916 4437 21925 4471
rect 21925 4437 21959 4471
rect 21959 4437 21968 4471
rect 21916 4428 21968 4437
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2412 4224 2464 4276
rect 1584 4199 1636 4208
rect 1584 4165 1593 4199
rect 1593 4165 1627 4199
rect 1627 4165 1636 4199
rect 1584 4156 1636 4165
rect 4068 4224 4120 4276
rect 7656 4224 7708 4276
rect 6000 4156 6052 4208
rect 6368 4156 6420 4208
rect 8668 4156 8720 4208
rect 9588 4224 9640 4276
rect 12164 4224 12216 4276
rect 12256 4224 12308 4276
rect 14096 4224 14148 4276
rect 11336 4156 11388 4208
rect 11520 4156 11572 4208
rect 12348 4156 12400 4208
rect 22744 4224 22796 4276
rect 23940 4224 23992 4276
rect 24492 4224 24544 4276
rect 22560 4156 22612 4208
rect 23388 4156 23440 4208
rect 2688 4088 2740 4140
rect 7196 4088 7248 4140
rect 7840 4088 7892 4140
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11244 4088 11296 4140
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 3700 4020 3752 4072
rect 5908 4020 5960 4072
rect 1860 3884 1912 3936
rect 6092 3884 6144 3936
rect 7932 3952 7984 4004
rect 9588 4020 9640 4072
rect 11704 4020 11756 4072
rect 9956 3952 10008 4004
rect 9772 3884 9824 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 11520 3884 11572 3936
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 17224 4088 17276 4140
rect 18052 4088 18104 4140
rect 19984 4088 20036 4140
rect 20076 4088 20128 4140
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 20996 4088 21048 4140
rect 23020 4088 23072 4140
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23756 4156 23808 4208
rect 23296 4088 23348 4097
rect 13636 4020 13688 4072
rect 14096 3884 14148 3936
rect 20536 4020 20588 4072
rect 20720 4020 20772 4072
rect 23756 4020 23808 4072
rect 15384 3952 15436 4004
rect 15936 3952 15988 4004
rect 18788 3952 18840 4004
rect 21272 3952 21324 4004
rect 21548 3952 21600 4004
rect 37188 4088 37240 4140
rect 36360 3952 36412 4004
rect 15476 3884 15528 3936
rect 21088 3884 21140 3936
rect 21180 3884 21232 3936
rect 25228 3927 25280 3936
rect 25228 3893 25237 3927
rect 25237 3893 25271 3927
rect 25271 3893 25280 3927
rect 25228 3884 25280 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 5356 3680 5408 3732
rect 5724 3680 5776 3732
rect 7932 3680 7984 3732
rect 9588 3680 9640 3732
rect 13268 3680 13320 3732
rect 16580 3680 16632 3732
rect 11980 3612 12032 3664
rect 14096 3612 14148 3664
rect 15936 3612 15988 3664
rect 16488 3612 16540 3664
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20352 3680 20404 3732
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3332 3544 3384 3596
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 8484 3544 8536 3596
rect 10140 3544 10192 3596
rect 12256 3544 12308 3596
rect 12348 3544 12400 3596
rect 14004 3544 14056 3596
rect 16856 3544 16908 3596
rect 17224 3544 17276 3596
rect 22284 3612 22336 3664
rect 21548 3587 21600 3596
rect 21548 3553 21557 3587
rect 21557 3553 21591 3587
rect 21591 3553 21600 3587
rect 21548 3544 21600 3553
rect 23480 3680 23532 3732
rect 33876 3680 33928 3732
rect 23204 3612 23256 3664
rect 23572 3612 23624 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 9680 3476 9732 3528
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 12716 3476 12768 3528
rect 17960 3476 18012 3528
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 20720 3476 20772 3528
rect 20996 3476 21048 3528
rect 22008 3476 22060 3528
rect 23020 3476 23072 3528
rect 24584 3519 24636 3528
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 4712 3408 4764 3460
rect 6644 3408 6696 3460
rect 7380 3408 7432 3460
rect 8024 3408 8076 3460
rect 4620 3340 4672 3392
rect 5816 3340 5868 3392
rect 10416 3408 10468 3460
rect 11152 3408 11204 3460
rect 11980 3408 12032 3460
rect 13268 3408 13320 3460
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 14280 3408 14332 3460
rect 14832 3340 14884 3392
rect 16488 3408 16540 3460
rect 16764 3408 16816 3460
rect 16948 3408 17000 3460
rect 18144 3408 18196 3460
rect 15936 3340 15988 3392
rect 16212 3340 16264 3392
rect 17040 3340 17092 3392
rect 17132 3340 17184 3392
rect 18512 3340 18564 3392
rect 20076 3340 20128 3392
rect 20444 3408 20496 3460
rect 22100 3408 22152 3460
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 27620 3476 27672 3528
rect 38108 3476 38160 3528
rect 37924 3408 37976 3460
rect 24768 3340 24820 3392
rect 36912 3340 36964 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3332 3136 3384 3188
rect 3976 3136 4028 3188
rect 11980 3136 12032 3188
rect 15660 3136 15712 3188
rect 16764 3136 16816 3188
rect 1584 3068 1636 3120
rect 3240 3000 3292 3052
rect 4804 3068 4856 3120
rect 5172 3068 5224 3120
rect 7472 3068 7524 3120
rect 9220 3068 9272 3120
rect 9404 3068 9456 3120
rect 11888 3068 11940 3120
rect 20444 3136 20496 3188
rect 20536 3136 20588 3188
rect 17132 3111 17184 3120
rect 17132 3077 17141 3111
rect 17141 3077 17175 3111
rect 17175 3077 17184 3111
rect 17132 3068 17184 3077
rect 21180 3068 21232 3120
rect 22008 3136 22060 3188
rect 25780 3179 25832 3188
rect 25780 3145 25789 3179
rect 25789 3145 25823 3179
rect 25823 3145 25832 3179
rect 25780 3136 25832 3145
rect 9496 3000 9548 3052
rect 1308 2932 1360 2984
rect 3332 2932 3384 2984
rect 3424 2932 3476 2984
rect 6460 2932 6512 2984
rect 6736 2932 6788 2984
rect 9036 2932 9088 2984
rect 13176 3000 13228 3052
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 15384 3000 15436 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 19432 3000 19484 3052
rect 20168 3000 20220 3052
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 22100 3068 22152 3120
rect 22008 3043 22060 3052
rect 13820 2932 13872 2984
rect 16028 2932 16080 2984
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 21272 2932 21324 2984
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 23020 3043 23072 3052
rect 22284 3000 22336 3009
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 23388 3000 23440 3052
rect 24768 3068 24820 3120
rect 36912 3043 36964 3052
rect 22192 2932 22244 2984
rect 22836 2932 22888 2984
rect 4896 2796 4948 2848
rect 5264 2796 5316 2848
rect 9588 2864 9640 2916
rect 9680 2864 9732 2916
rect 13636 2864 13688 2916
rect 9036 2796 9088 2848
rect 11612 2796 11664 2848
rect 12440 2796 12492 2848
rect 19340 2864 19392 2916
rect 19432 2907 19484 2916
rect 19432 2873 19441 2907
rect 19441 2873 19475 2907
rect 19475 2873 19484 2907
rect 19432 2864 19484 2873
rect 19616 2864 19668 2916
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 38016 3043 38068 3052
rect 38016 3009 38025 3043
rect 38025 3009 38059 3043
rect 38059 3009 38068 3043
rect 38016 3000 38068 3009
rect 27528 2932 27580 2984
rect 19156 2796 19208 2848
rect 20168 2796 20220 2848
rect 23112 2796 23164 2848
rect 38016 2796 38068 2848
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5632 2592 5684 2644
rect 13452 2592 13504 2644
rect 14004 2592 14056 2644
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 18604 2592 18656 2644
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 19064 2592 19116 2644
rect 23664 2592 23716 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 8484 2567 8536 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 8484 2533 8493 2567
rect 8493 2533 8527 2567
rect 8527 2533 8536 2567
rect 8484 2524 8536 2533
rect 9128 2524 9180 2576
rect 6000 2499 6052 2508
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 4712 2320 4764 2372
rect 5540 2252 5592 2304
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 10048 2456 10100 2508
rect 11520 2456 11572 2508
rect 14096 2456 14148 2508
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 16580 2388 16632 2440
rect 8300 2320 8352 2372
rect 8576 2320 8628 2372
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 14096 2320 14148 2372
rect 14188 2320 14240 2372
rect 15568 2320 15620 2372
rect 19340 2524 19392 2576
rect 27528 2524 27580 2576
rect 33600 2635 33652 2644
rect 33600 2601 33609 2635
rect 33609 2601 33643 2635
rect 33643 2601 33652 2635
rect 33600 2592 33652 2601
rect 30288 2524 30340 2576
rect 16764 2252 16816 2304
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 17960 2320 18012 2372
rect 20260 2388 20312 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 23572 2388 23624 2440
rect 23756 2388 23808 2440
rect 33048 2456 33100 2508
rect 24676 2388 24728 2440
rect 27068 2388 27120 2440
rect 29000 2388 29052 2440
rect 30288 2388 30340 2440
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33508 2388 33560 2440
rect 34796 2388 34848 2440
rect 38016 2431 38068 2440
rect 38016 2397 38025 2431
rect 38025 2397 38059 2431
rect 38059 2397 38068 2431
rect 38016 2388 38068 2397
rect 22284 2363 22336 2372
rect 22284 2329 22293 2363
rect 22293 2329 22327 2363
rect 22327 2329 22336 2363
rect 22284 2320 22336 2329
rect 17868 2252 17920 2304
rect 19340 2252 19392 2304
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 22560 2252 22612 2304
rect 23480 2252 23532 2304
rect 23848 2252 23900 2304
rect 25780 2252 25832 2304
rect 31576 2252 31628 2304
rect 36084 2252 36136 2304
rect 39304 2252 39356 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 5172 2048 5224 2100
rect 1860 1980 1912 2032
rect 7932 1980 7984 2032
rect 8484 1980 8536 2032
rect 14096 1980 14148 2032
rect 17868 2048 17920 2100
rect 19432 2048 19484 2100
rect 14464 1912 14516 1964
rect 12072 1844 12124 1896
rect 15936 1844 15988 1896
rect 25228 1980 25280 2032
rect 20904 1912 20956 1964
rect 18972 1844 19024 1896
rect 24032 1844 24084 1896
rect 10968 1708 11020 1760
rect 22284 1708 22336 1760
rect 15568 1640 15620 1692
rect 21916 1640 21968 1692
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 32 37330 60 39200
rect 20 37324 72 37330
rect 20 37266 72 37272
rect 1320 37262 1348 39200
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2792 37262 2820 38111
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 1308 37256 1360 37262
rect 1308 37198 1360 37204
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4632 37126 4660 37726
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 5356 37188 5408 37194
rect 5356 37130 5408 37136
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 2872 37120 2924 37126
rect 2872 37062 2924 37068
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 1596 36922 1624 37062
rect 1584 36916 1636 36922
rect 1584 36858 1636 36864
rect 1766 36816 1822 36825
rect 1766 36751 1768 36760
rect 1820 36751 1822 36760
rect 1768 36722 1820 36728
rect 2688 36576 2740 36582
rect 2688 36518 2740 36524
rect 1766 33416 1822 33425
rect 1766 33351 1768 33360
rect 1820 33351 1822 33360
rect 1768 33322 1820 33328
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1780 32065 1808 32370
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 2700 30734 2728 36518
rect 1768 30728 1820 30734
rect 1766 30696 1768 30705
rect 2688 30728 2740 30734
rect 1820 30696 1822 30705
rect 2688 30670 2740 30676
rect 1766 30631 1822 30640
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28665 1808 29106
rect 2884 29102 2912 37062
rect 3988 36854 4016 37062
rect 3976 36848 4028 36854
rect 3976 36790 4028 36796
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3436 29306 3464 33458
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 5368 32434 5396 37130
rect 5460 34202 5488 37198
rect 5828 37126 5856 39200
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 6564 36922 6592 37198
rect 7760 37126 7788 39200
rect 9048 37262 9076 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 6460 36916 6512 36922
rect 6460 36858 6512 36864
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 5448 34196 5500 34202
rect 5448 34138 5500 34144
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5540 30864 5592 30870
rect 5540 30806 5592 30812
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 2872 29096 2924 29102
rect 2872 29038 2924 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 25288 1820 25294
rect 1766 25256 1768 25265
rect 1820 25256 1822 25265
rect 1766 25191 1822 25200
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 3988 23866 4016 27406
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5552 25906 5580 30806
rect 6092 30592 6144 30598
rect 6092 30534 6144 30540
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 1766 23831 1822 23840
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 4080 21554 4108 25094
rect 6104 24818 6132 30534
rect 6472 30258 6500 36858
rect 7852 33114 7880 37198
rect 10336 37126 10364 39200
rect 10416 37256 10468 37262
rect 12268 37244 12296 39200
rect 12440 37256 12492 37262
rect 12268 37216 12440 37244
rect 10416 37198 10468 37204
rect 12440 37198 12492 37204
rect 9312 37120 9364 37126
rect 9312 37062 9364 37068
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6748 26994 6776 32166
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6092 24812 6144 24818
rect 6092 24754 6144 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5552 22778 5580 23666
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 19145 1808 19314
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 2780 14408 2832 14414
rect 1820 14376 1822 14385
rect 2780 14350 2832 14356
rect 1766 14311 1822 14320
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 1582 13968 1638 13977
rect 1582 13903 1584 13912
rect 1636 13903 1638 13912
rect 1584 13874 1636 13880
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1308 8900 1360 8906
rect 1308 8842 1360 8848
rect 20 5024 72 5030
rect 20 4966 72 4972
rect 32 800 60 4966
rect 1320 4865 1348 8842
rect 1412 7585 1440 13262
rect 2240 12850 2268 13670
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 1780 12345 1808 12786
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 11898 1624 12038
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1400 7472 1452 7478
rect 1400 7414 1452 7420
rect 1412 6458 1440 7414
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1504 6338 1532 11698
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 9586 1716 10406
rect 1780 9625 1808 10610
rect 1766 9616 1822 9625
rect 1676 9580 1728 9586
rect 1766 9551 1822 9560
rect 1676 9522 1728 9528
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 6866 1624 8298
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1584 6724 1636 6730
rect 1688 6712 1716 7754
rect 1872 7478 1900 11494
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1636 6684 1716 6712
rect 1584 6666 1636 6672
rect 1412 6310 1532 6338
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 800 1348 2926
rect 1412 2825 1440 6310
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 5710 1532 6190
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1504 4622 1532 5646
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1504 4026 1532 4558
rect 1596 4214 1624 6666
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1688 5234 1716 6394
rect 1780 6322 1808 6802
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 2056 5098 2084 8774
rect 2240 5234 2268 12582
rect 2332 5642 2360 13806
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11762 2452 12038
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 2424 4282 2452 8774
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1504 3998 1624 4026
rect 1596 3534 1624 3998
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3602 1900 3878
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3126 1624 3470
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1596 2514 1624 3062
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 2038 1900 2314
rect 1860 2032 1912 2038
rect 1860 1974 1912 1980
rect 2516 1952 2544 10610
rect 2608 6118 2636 14214
rect 2792 13938 2820 14350
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13326 2820 13874
rect 3056 13864 3108 13870
rect 3054 13832 3056 13841
rect 3108 13832 3110 13841
rect 3054 13767 3110 13776
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2792 9586 2820 12174
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2872 11688 2924 11694
rect 2924 11648 3004 11676
rect 2872 11630 2924 11636
rect 2976 10606 3004 11648
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 10130 3004 10542
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2792 8974 2820 9522
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9042 2912 9454
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2700 7546 2728 8026
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2792 7410 2820 8910
rect 3068 8906 3096 12106
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8498 2912 8774
rect 3054 8664 3110 8673
rect 3160 8650 3188 14894
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3252 12238 3280 12786
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3110 8622 3188 8650
rect 3054 8599 3110 8608
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2964 8424 3016 8430
rect 2870 8392 2926 8401
rect 2964 8366 3016 8372
rect 2870 8327 2872 8336
rect 2924 8327 2926 8336
rect 2872 8298 2924 8304
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6254 2728 6598
rect 2884 6458 2912 8298
rect 2976 7818 3004 8366
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 6769 3004 7346
rect 3252 6866 3280 9318
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 2962 6760 3018 6769
rect 2962 6695 3018 6704
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2596 5772 2648 5778
rect 2700 5760 2728 6190
rect 2648 5732 2728 5760
rect 2596 5714 2648 5720
rect 2700 5234 2728 5732
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2700 4146 2728 5170
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2516 1924 2636 1952
rect 2608 800 2636 1924
rect 2792 1465 2820 4966
rect 3160 4758 3188 6190
rect 3344 4826 3372 20334
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3620 13326 3648 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12782 4016 13262
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3988 12238 4016 12718
rect 4080 12617 4108 12786
rect 4066 12608 4122 12617
rect 4066 12543 4122 12552
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4618 12472 4674 12481
rect 4618 12407 4674 12416
rect 4632 12306 4660 12407
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 10266 3464 10542
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3436 9178 3464 9386
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3436 7410 3464 8978
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3056 4752 3108 4758
rect 3054 4720 3056 4729
rect 3148 4752 3200 4758
rect 3108 4720 3110 4729
rect 3148 4694 3200 4700
rect 3054 4655 3110 4664
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3252 3058 3280 4626
rect 3344 4162 3372 4762
rect 3436 4690 3464 7346
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3528 4554 3556 11222
rect 3620 10962 3648 12038
rect 3804 11098 3832 12174
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11762 4660 12038
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4160 11620 4212 11626
rect 3988 11580 4160 11608
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 11218 3924 11494
rect 3988 11286 4016 11580
rect 4160 11562 4212 11568
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4080 11234 4108 11290
rect 3884 11212 3936 11218
rect 4080 11206 4200 11234
rect 3884 11154 3936 11160
rect 3976 11144 4028 11150
rect 3804 11070 3924 11098
rect 3976 11086 4028 11092
rect 3620 10934 3832 10962
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9110 3648 9318
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 7818 3648 8910
rect 3712 8430 3740 10746
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3804 8276 3832 10934
rect 3896 8294 3924 11070
rect 3988 10062 4016 11086
rect 4172 10810 4200 11206
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4250 10840 4306 10849
rect 4160 10804 4212 10810
rect 4250 10775 4306 10784
rect 4160 10746 4212 10752
rect 4264 10554 4292 10775
rect 4080 10526 4292 10554
rect 4540 10554 4568 10950
rect 4632 10849 4660 11494
rect 4618 10840 4674 10849
rect 4618 10775 4674 10784
rect 4540 10526 4660 10554
rect 4080 10198 4108 10526
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9518 4016 9998
rect 4632 9874 4660 10526
rect 4724 10266 4752 21286
rect 5552 19854 5580 22374
rect 6196 21146 6224 24142
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 7484 20806 7512 32166
rect 8772 28218 8800 33934
rect 9324 30734 9352 37062
rect 9404 36848 9456 36854
rect 9404 36790 9456 36796
rect 9416 30734 9444 36790
rect 10428 34202 10456 37198
rect 13556 37126 13584 39200
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 10704 35290 10732 36722
rect 10692 35284 10744 35290
rect 10692 35226 10744 35232
rect 12256 35080 12308 35086
rect 12256 35022 12308 35028
rect 10416 34196 10468 34202
rect 10416 34138 10468 34144
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11336 30864 11388 30870
rect 11336 30806 11388 30812
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9312 29232 9364 29238
rect 9312 29174 9364 29180
rect 8760 28212 8812 28218
rect 8760 28154 8812 28160
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5184 17678 5212 19450
rect 5828 19378 5856 20742
rect 7944 20602 7972 20878
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 6932 19378 6960 20402
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7024 19990 7052 20198
rect 8404 20058 8432 20402
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19530 8432 19790
rect 8496 19718 8524 21898
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19530 8616 19654
rect 8404 19502 8616 19530
rect 8496 19446 8524 19502
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 6932 18834 6960 19314
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 6920 18828 6972 18834
rect 8220 18816 8248 19246
rect 8484 18828 8536 18834
rect 8220 18788 8484 18816
rect 6920 18770 6972 18776
rect 8484 18770 8536 18776
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 18426 6684 18702
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4816 14618 4844 16050
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4632 9846 4752 9874
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 8974 4016 9454
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4080 8634 4108 9590
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8634 4200 8774
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4526 8392 4582 8401
rect 4526 8327 4528 8336
rect 4580 8327 4582 8336
rect 4528 8298 4580 8304
rect 3712 8248 3832 8276
rect 3884 8288 3936 8294
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3620 7410 3648 7754
rect 3712 7478 3740 8248
rect 3884 8230 3936 8236
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3700 7472 3752 7478
rect 3896 7426 3924 8230
rect 3700 7414 3752 7420
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3804 7398 3924 7426
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3620 6254 3648 6326
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3344 4134 3464 4162
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3344 3602 3372 4014
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3344 2990 3372 3130
rect 3436 2990 3464 4134
rect 3712 4078 3740 6938
rect 3804 6361 3832 7398
rect 3790 6352 3846 6361
rect 3790 6287 3846 6296
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3988 3194 4016 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7818 4660 9658
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 4282 4108 7210
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 7754
rect 4724 6458 4752 9846
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4622 4660 5102
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4250 3496 4306 3505
rect 4250 3431 4252 3440
rect 4304 3431 4306 3440
rect 4252 3402 4304 3408
rect 4632 3398 4660 4422
rect 4724 3466 4752 6054
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4816 3126 4844 12650
rect 4908 9722 4936 16050
rect 5552 15502 5580 18022
rect 6932 17921 6960 18770
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7300 18290 7328 18702
rect 8588 18630 8616 19314
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 6918 17912 6974 17921
rect 6918 17847 6974 17856
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17202 6960 17478
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16114 7144 16526
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14414 5028 14758
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5000 9602 5028 13330
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4908 9574 5028 9602
rect 4908 6730 4936 9574
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 8401 5028 8502
rect 4986 8392 5042 8401
rect 4986 8327 5042 8336
rect 4986 8256 5042 8265
rect 4986 8191 5042 8200
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 4908 2854 4936 6394
rect 5000 5778 5028 8191
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4988 5228 5040 5234
rect 5092 5216 5120 13194
rect 5170 13152 5226 13161
rect 5170 13087 5226 13096
rect 5184 7342 5212 13087
rect 5552 12442 5580 13942
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5446 11792 5502 11801
rect 5368 10305 5396 11766
rect 5446 11727 5502 11736
rect 5354 10296 5410 10305
rect 5264 10260 5316 10266
rect 5354 10231 5410 10240
rect 5264 10202 5316 10208
rect 5276 8838 5304 10202
rect 5264 8832 5316 8838
rect 5316 8792 5396 8820
rect 5264 8774 5316 8780
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5276 8090 5304 8502
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5040 5188 5120 5216
rect 4988 5170 5040 5176
rect 5184 3126 5212 7278
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5276 6662 5304 6870
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5276 2938 5304 6326
rect 5368 3738 5396 8792
rect 5460 8430 5488 11727
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 7206 5488 8230
rect 5552 7818 5580 12106
rect 5644 10062 5672 13806
rect 6380 13734 6408 14554
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5736 11286 5764 11630
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5724 10736 5776 10742
rect 5722 10704 5724 10713
rect 5776 10704 5778 10713
rect 5828 10674 5856 13398
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6012 12617 6040 12786
rect 5998 12608 6054 12617
rect 5998 12543 6054 12552
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5920 12238 5948 12378
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5722 10639 5778 10648
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5920 9874 5948 12174
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6274 11520 6330 11529
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10441 6132 11086
rect 6090 10432 6146 10441
rect 6090 10367 6146 10376
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5644 9846 5948 9874
rect 5644 9330 5672 9846
rect 6012 9518 6040 10066
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5724 9512 5776 9518
rect 6000 9512 6052 9518
rect 5998 9480 6000 9489
rect 6052 9480 6054 9489
rect 5776 9460 5948 9466
rect 5724 9454 5948 9460
rect 5736 9450 5948 9454
rect 5736 9444 5960 9450
rect 5736 9438 5908 9444
rect 5998 9415 6054 9424
rect 5908 9386 5960 9392
rect 5644 9302 5764 9330
rect 5736 8974 5764 9302
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5736 8498 5764 8910
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5644 5522 5672 8298
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5552 5494 5672 5522
rect 5448 4616 5500 4622
rect 5446 4584 5448 4593
rect 5500 4584 5502 4593
rect 5446 4519 5502 4528
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5184 2910 5304 2938
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4710 2544 4766 2553
rect 4710 2479 4766 2488
rect 4724 2378 4752 2479
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 5184 2106 5212 2910
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 5276 898 5304 2790
rect 5552 2310 5580 5494
rect 5736 5370 5764 6802
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 2650 5672 4422
rect 5736 3738 5764 5102
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5828 3398 5856 8774
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5920 7002 5948 7278
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5906 6352 5962 6361
rect 5906 6287 5908 6296
rect 5960 6287 5962 6296
rect 5908 6258 5960 6264
rect 6012 5846 6040 7142
rect 6104 6934 6132 9862
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6012 4298 6040 5782
rect 6196 4842 6224 11494
rect 6274 11455 6330 11464
rect 6288 9926 6316 11455
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6380 6866 6408 13670
rect 6564 12918 6592 14486
rect 7208 14074 7236 15370
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6472 12238 6500 12854
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6458 12064 6514 12073
rect 6458 11999 6514 12008
rect 6472 8634 6500 11999
rect 6552 9104 6604 9110
rect 6550 9072 6552 9081
rect 6604 9072 6606 9081
rect 6550 9007 6606 9016
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6276 6792 6328 6798
rect 6274 6760 6276 6769
rect 6328 6760 6330 6769
rect 6274 6695 6330 6704
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 5545 6316 6598
rect 6368 6248 6420 6254
rect 6366 6216 6368 6225
rect 6420 6216 6422 6225
rect 6564 6186 6592 8910
rect 6656 7290 6684 13126
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 9994 6776 11086
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 9518 6776 9930
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 8974 6776 9454
rect 6840 9450 6868 13398
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7116 12434 7144 12786
rect 7116 12406 7236 12434
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6932 10266 6960 12242
rect 7208 12238 7236 12406
rect 7196 12232 7248 12238
rect 7010 12200 7066 12209
rect 7196 12174 7248 12180
rect 7010 12135 7066 12144
rect 7024 12102 7052 12135
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8430 6776 8910
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 7954 6776 8366
rect 6840 7954 6868 9386
rect 7024 8498 7052 11863
rect 7116 11200 7144 12038
rect 7208 11694 7236 12174
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7116 11172 7236 11200
rect 7102 11112 7158 11121
rect 7102 11047 7104 11056
rect 7156 11047 7158 11056
rect 7104 11018 7156 11024
rect 7208 10169 7236 11172
rect 7300 10985 7328 18226
rect 8312 17814 8340 18566
rect 8496 18442 8524 18566
rect 8680 18442 8708 20810
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8772 18970 8800 19178
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8496 18414 8708 18442
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 16522 7696 17614
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7668 16114 7696 16458
rect 7944 16250 7972 16526
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7392 13326 7420 13874
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7286 10976 7342 10985
rect 7286 10911 7342 10920
rect 7392 10826 7420 13262
rect 7668 13161 7696 16050
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15638 7880 15846
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14074 7788 14894
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7654 13152 7710 13161
rect 7654 13087 7710 13096
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7562 11928 7618 11937
rect 7562 11863 7618 11872
rect 7576 11762 7604 11863
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7472 11688 7524 11694
rect 7470 11656 7472 11665
rect 7524 11656 7526 11665
rect 7470 11591 7526 11600
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7470 11384 7526 11393
rect 7470 11319 7526 11328
rect 7300 10798 7420 10826
rect 7194 10160 7250 10169
rect 7300 10146 7328 10798
rect 7484 10470 7512 11319
rect 7576 11082 7604 11494
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7562 10976 7618 10985
rect 7562 10911 7618 10920
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7300 10118 7512 10146
rect 7194 10095 7250 10104
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6748 7410 6776 7890
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6656 7262 6776 7290
rect 6642 6488 6698 6497
rect 6642 6423 6698 6432
rect 6366 6151 6422 6160
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6564 5817 6592 6122
rect 6550 5808 6606 5817
rect 6550 5743 6606 5752
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6274 5536 6330 5545
rect 6274 5471 6330 5480
rect 6380 5030 6408 5578
rect 6656 5574 6684 6423
rect 6748 6390 6776 7262
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 6458 7052 6666
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6918 6216 6974 6225
rect 6918 6151 6974 6160
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6104 4826 6224 4842
rect 6092 4820 6224 4826
rect 6144 4814 6224 4820
rect 6092 4762 6144 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6012 4270 6132 4298
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5920 2774 5948 4014
rect 5828 2746 5948 2774
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 4540 870 4660 898
rect 4540 800 4568 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 4632 762 4660 870
rect 5000 870 5304 898
rect 5000 762 5028 870
rect 5828 800 5856 2746
rect 6012 2514 6040 4150
rect 6104 3942 6132 4270
rect 6380 4214 6408 4490
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6472 3602 6500 4626
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 2990 6500 3538
rect 6656 3466 6684 5510
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6840 5137 6868 5170
rect 6826 5128 6882 5137
rect 6826 5063 6882 5072
rect 6932 4554 6960 6151
rect 7024 5778 7052 6394
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5234 7052 5714
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7024 4690 7052 5170
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6748 2514 6776 2926
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7116 800 7144 8570
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7208 6730 7236 7482
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7194 5808 7250 5817
rect 7194 5743 7196 5752
rect 7248 5743 7250 5752
rect 7196 5714 7248 5720
rect 7194 5400 7250 5409
rect 7300 5370 7328 9930
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7194 5335 7250 5344
rect 7288 5364 7340 5370
rect 7208 5302 7236 5335
rect 7288 5306 7340 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7208 4146 7236 5238
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7392 3466 7420 8774
rect 7484 7342 7512 10118
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 7206 7604 10911
rect 7668 9738 7696 12718
rect 7760 12238 7788 13262
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 10606 7788 12174
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7668 9710 7788 9738
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7668 8566 7696 9590
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7484 3126 7512 6802
rect 7760 5370 7788 9710
rect 7852 7546 7880 13806
rect 7944 13530 7972 13874
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8036 13274 8064 15914
rect 8312 15706 8340 17070
rect 8404 16794 8432 18226
rect 8680 17882 8708 18226
rect 8864 17882 8892 19314
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8956 17746 8984 26726
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9140 21554 9168 21830
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 9048 18222 9076 19722
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9140 18068 9168 19654
rect 9232 18986 9260 23258
rect 9324 22642 9352 29174
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 20398 9352 21490
rect 9600 21146 9628 25638
rect 10152 25498 10180 29106
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9692 22030 9720 22578
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9692 21350 9720 21966
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19174 9352 19790
rect 9416 19786 9444 20198
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9232 18958 9352 18986
rect 9324 18290 9352 18958
rect 9600 18834 9628 19450
rect 9692 19174 9720 20402
rect 9784 19922 9812 24754
rect 10416 22704 10468 22710
rect 10416 22646 10468 22652
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9770 19544 9826 19553
rect 9770 19479 9826 19488
rect 9784 19446 9812 19479
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9862 19408 9918 19417
rect 9862 19343 9864 19352
rect 9916 19343 9918 19352
rect 9864 19314 9916 19320
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9692 18766 9720 19110
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9324 18193 9352 18226
rect 9310 18184 9366 18193
rect 9770 18184 9826 18193
rect 9310 18119 9366 18128
rect 9588 18148 9640 18154
rect 9770 18119 9772 18128
rect 9588 18090 9640 18096
rect 9824 18119 9826 18128
rect 9772 18090 9824 18096
rect 9140 18040 9352 18068
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8680 17202 8708 17614
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8588 16250 8616 17138
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 16726 8800 16934
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14618 8156 14962
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8220 13938 8248 15438
rect 8404 14822 8432 15846
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8312 13870 8340 14758
rect 8956 14498 8984 16526
rect 9048 14770 9076 17614
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9140 16590 9168 17546
rect 9232 16794 9260 17546
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9324 16538 9352 18040
rect 9600 17882 9628 18090
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9968 17746 9996 19994
rect 10060 19718 10088 22102
rect 10244 21622 10272 22510
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10232 21412 10284 21418
rect 10232 21354 10284 21360
rect 10048 19712 10100 19718
rect 10046 19680 10048 19689
rect 10100 19680 10102 19689
rect 10046 19615 10102 19624
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10060 17746 10088 18090
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9600 17134 9628 17682
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9416 16658 9444 17070
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9784 16794 9812 17138
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9324 16510 9444 16538
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 15366 9168 15438
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9048 14742 9168 14770
rect 8956 14470 9076 14498
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8300 13864 8352 13870
rect 8206 13832 8262 13841
rect 8300 13806 8352 13812
rect 8206 13767 8262 13776
rect 8036 13246 8156 13274
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12434 7972 12786
rect 8036 12646 8064 13126
rect 8128 12850 8156 13246
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 7944 12406 8064 12434
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7852 5914 7880 7482
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7944 5778 7972 11562
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7838 5536 7894 5545
rect 7838 5471 7894 5480
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7852 5302 7880 5471
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 4758 7972 5714
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7654 4312 7710 4321
rect 7654 4247 7656 4256
rect 7708 4247 7710 4256
rect 7656 4218 7708 4224
rect 7852 4146 7880 4558
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7944 3738 7972 3946
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8036 3466 8064 12406
rect 8128 10538 8156 12582
rect 8220 11626 8248 13767
rect 8298 12336 8354 12345
rect 8404 12322 8432 14350
rect 8496 12442 8524 14350
rect 9048 14278 9076 14470
rect 9140 14385 9168 14742
rect 9126 14376 9182 14385
rect 9126 14311 9182 14320
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 13161 8708 13194
rect 8666 13152 8722 13161
rect 8666 13087 8722 13096
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8574 12472 8630 12481
rect 8484 12436 8536 12442
rect 8574 12407 8576 12416
rect 8484 12378 8536 12384
rect 8628 12407 8630 12416
rect 8772 12434 8800 12718
rect 8772 12406 8892 12434
rect 8576 12378 8628 12384
rect 8404 12294 8800 12322
rect 8298 12271 8300 12280
rect 8352 12271 8354 12280
rect 8300 12242 8352 12248
rect 8576 12232 8628 12238
rect 8482 12200 8538 12209
rect 8576 12174 8628 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8482 12135 8538 12144
rect 8496 12102 8524 12135
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8300 11892 8352 11898
rect 8404 11880 8432 12038
rect 8484 11892 8536 11898
rect 8404 11852 8484 11880
rect 8300 11834 8352 11840
rect 8484 11834 8536 11840
rect 8312 11778 8340 11834
rect 8588 11778 8616 12174
rect 8680 11801 8708 12174
rect 8312 11750 8616 11778
rect 8666 11792 8722 11801
rect 8666 11727 8722 11736
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8668 11688 8720 11694
rect 8772 11665 8800 12294
rect 8668 11630 8720 11636
rect 8758 11656 8814 11665
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8220 11257 8248 11290
rect 8312 11286 8340 11630
rect 8300 11280 8352 11286
rect 8206 11248 8262 11257
rect 8300 11222 8352 11228
rect 8206 11183 8262 11192
rect 8392 11144 8444 11150
rect 8680 11121 8708 11630
rect 8758 11591 8814 11600
rect 8392 11086 8444 11092
rect 8666 11112 8722 11121
rect 8404 10742 8432 11086
rect 8666 11047 8722 11056
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8128 9994 8156 10202
rect 8220 10130 8248 10542
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8312 9738 8340 9998
rect 8220 9710 8340 9738
rect 8496 9722 8524 10678
rect 8574 10568 8630 10577
rect 8574 10503 8630 10512
rect 8588 10062 8616 10503
rect 8680 10198 8708 10950
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9716 8536 9722
rect 8220 9586 8248 9710
rect 8484 9658 8536 9664
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8114 8528 8170 8537
rect 8114 8463 8170 8472
rect 8128 8430 8156 8463
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8220 5953 8248 8910
rect 8772 8906 8800 11591
rect 8864 9081 8892 12406
rect 8956 12374 8984 12922
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8850 9072 8906 9081
rect 8850 9007 8906 9016
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 6730 8432 8774
rect 8956 7698 8984 11834
rect 8496 7670 8984 7698
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8300 6112 8352 6118
rect 8496 6100 8524 7670
rect 9048 7562 9076 14214
rect 9140 13818 9168 14311
rect 9232 13938 9260 14826
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9416 13852 9444 16510
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9600 14890 9628 15642
rect 9692 15502 9720 16730
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9784 15502 9812 15982
rect 9876 15978 9904 16050
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9876 15881 9904 15914
rect 9862 15872 9918 15881
rect 9862 15807 9918 15816
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 15162 9812 15302
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9692 14074 9720 14962
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9508 13954 9536 14010
rect 9876 13988 9904 15438
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9784 13960 9904 13988
rect 9784 13954 9812 13960
rect 9508 13926 9812 13954
rect 9968 13938 9996 14282
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9416 13824 9628 13852
rect 9140 13790 9260 13818
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9140 10470 9168 12922
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8352 6072 8524 6100
rect 8588 7534 9076 7562
rect 8300 6054 8352 6060
rect 8206 5944 8262 5953
rect 8206 5879 8262 5888
rect 8312 5817 8340 6054
rect 8298 5808 8354 5817
rect 8298 5743 8354 5752
rect 8392 5704 8444 5710
rect 8206 5672 8262 5681
rect 8392 5646 8444 5652
rect 8206 5607 8208 5616
rect 8260 5607 8262 5616
rect 8208 5578 8260 5584
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8220 4486 8248 5306
rect 8404 4622 8432 5646
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8496 4162 8524 5510
rect 8312 4134 8524 4162
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 8036 2774 8064 3402
rect 7944 2746 8064 2774
rect 7944 2038 7972 2746
rect 8312 2378 8340 4134
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8496 2582 8524 3538
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8496 2038 8524 2518
rect 8588 2378 8616 7534
rect 9232 6866 9260 13790
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9324 12918 9352 13738
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9310 12336 9366 12345
rect 9310 12271 9312 12280
rect 9364 12271 9366 12280
rect 9312 12242 9364 12248
rect 9416 11898 9444 12854
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11354 9352 11698
rect 9404 11688 9456 11694
rect 9508 11665 9536 13126
rect 9600 12753 9628 13824
rect 9770 13696 9826 13705
rect 9770 13631 9826 13640
rect 9784 12918 9812 13631
rect 9954 13424 10010 13433
rect 9954 13359 9956 13368
rect 10008 13359 10010 13368
rect 9956 13330 10008 13336
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9586 12744 9642 12753
rect 9586 12679 9642 12688
rect 9588 11688 9640 11694
rect 9404 11630 9456 11636
rect 9494 11656 9550 11665
rect 9416 11354 9444 11630
rect 9588 11630 9640 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9494 11591 9550 11600
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9496 11144 9548 11150
rect 9600 11121 9628 11630
rect 9784 11558 9812 11630
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 11144 9732 11150
rect 9496 11086 9548 11092
rect 9586 11112 9642 11121
rect 9508 10538 9536 11086
rect 9680 11086 9732 11092
rect 9586 11047 9642 11056
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9600 8974 9628 10095
rect 9692 9178 9720 11086
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 8974 9812 11154
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9312 8832 9364 8838
rect 9416 8820 9444 8910
rect 9416 8792 9628 8820
rect 9312 8774 9364 8780
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9232 6390 9260 6802
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8680 5574 8708 6190
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 8956 5710 8984 5743
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 9034 5400 9090 5409
rect 9034 5335 9036 5344
rect 9088 5335 9090 5344
rect 9036 5306 9088 5312
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4214 8708 4422
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 9048 2990 9076 5306
rect 9140 4690 9168 5646
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 7932 2032 7984 2038
rect 7932 1974 7984 1980
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 9048 800 9076 2790
rect 9140 2582 9168 3334
rect 9232 3126 9260 6190
rect 9324 4826 9352 8774
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9416 8537 9444 8570
rect 9402 8528 9458 8537
rect 9402 8463 9458 8472
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9416 7750 9444 8298
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 7478 9444 7686
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 5817 9444 6734
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9402 5808 9458 5817
rect 9508 5778 9536 6598
rect 9402 5743 9458 5752
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5273 9536 5578
rect 9494 5264 9550 5273
rect 9494 5199 9550 5208
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9416 2446 9444 3062
rect 9508 3058 9536 5102
rect 9600 4554 9628 8792
rect 9876 7886 9904 13262
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12238 9996 13194
rect 10060 12442 10088 17682
rect 10244 16114 10272 21354
rect 10336 20534 10364 22374
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 10428 20398 10456 22646
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10692 21616 10744 21622
rect 10520 21564 10692 21570
rect 10520 21558 10744 21564
rect 10520 21542 10732 21558
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10336 19242 10364 20334
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 10336 18970 10364 19178
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10336 16658 10364 17546
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 10470 10088 12038
rect 10152 10826 10180 15846
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 12209 10272 13874
rect 10230 12200 10286 12209
rect 10230 12135 10286 12144
rect 10244 11529 10272 12135
rect 10230 11520 10286 11529
rect 10230 11455 10286 11464
rect 10336 11218 10364 16594
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16182 10456 16390
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10414 16008 10470 16017
rect 10414 15943 10416 15952
rect 10468 15943 10470 15952
rect 10416 15914 10468 15920
rect 10520 15910 10548 21542
rect 10796 21418 10824 21966
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 19242 10640 20266
rect 10704 20058 10732 21014
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10600 18352 10652 18358
rect 10652 18312 10732 18340
rect 10600 18294 10652 18300
rect 10704 16658 10732 18312
rect 10888 16658 10916 22442
rect 11072 21418 11100 28018
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11072 20534 11100 21354
rect 11164 21010 11192 21830
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11256 20602 11284 21898
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11348 19378 11376 30806
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11440 19417 11468 21830
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 19854 11560 20198
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11426 19408 11482 19417
rect 11336 19372 11388 19378
rect 11426 19343 11482 19352
rect 11336 19314 11388 19320
rect 11348 18766 11376 19314
rect 11624 19310 11652 29990
rect 11808 28218 11836 32846
rect 12268 31822 12296 35022
rect 12360 33522 12388 37062
rect 14292 34202 14320 37198
rect 15488 37126 15516 39200
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15764 36378 15792 37198
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15936 36168 15988 36174
rect 15936 36110 15988 36116
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 13636 33992 13688 33998
rect 13636 33934 13688 33940
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11716 20262 11744 20810
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11808 19310 11836 22034
rect 11992 19961 12020 30534
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12084 20806 12112 21966
rect 12360 21894 12388 25230
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12072 20800 12124 20806
rect 12070 20768 12072 20777
rect 12124 20768 12126 20777
rect 12070 20703 12126 20712
rect 12176 20534 12204 21286
rect 12452 20874 12480 21286
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12268 20262 12296 20470
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11978 19952 12034 19961
rect 11978 19887 12034 19896
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10980 17270 11008 17818
rect 11164 17542 11192 18022
rect 11624 17610 11652 19246
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18222 11744 18566
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11716 17882 11744 18158
rect 11808 18154 11836 18770
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11808 17762 11836 18090
rect 11716 17734 11836 17762
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11060 17536 11112 17542
rect 11058 17504 11060 17513
rect 11152 17536 11204 17542
rect 11112 17504 11114 17513
rect 11152 17478 11204 17484
rect 11058 17439 11114 17448
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10612 14550 10640 15982
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10704 14074 10732 15506
rect 10796 14550 10824 16050
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10416 13932 10468 13938
rect 10600 13932 10652 13938
rect 10416 13874 10468 13880
rect 10520 13892 10600 13920
rect 10428 13326 10456 13874
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10414 11928 10470 11937
rect 10414 11863 10470 11872
rect 10428 11626 10456 11863
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10520 11558 10548 13892
rect 10600 13874 10652 13880
rect 10796 13818 10824 14486
rect 10612 13790 10824 13818
rect 10888 13802 10916 15846
rect 11072 15094 11100 15914
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10876 13796 10928 13802
rect 10612 13002 10640 13790
rect 10876 13738 10928 13744
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10876 13320 10928 13326
rect 10704 13268 10876 13274
rect 10704 13262 10928 13268
rect 10704 13246 10916 13262
rect 10704 13190 10732 13246
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 13025 10916 13126
rect 10874 13016 10930 13025
rect 10612 12974 10732 13002
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10152 10798 10364 10826
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9586 4312 9642 4321
rect 9586 4247 9588 4256
rect 9640 4247 9642 4256
rect 9588 4218 9640 4224
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3738 9628 4014
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9692 3618 9720 7278
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9968 6866 9996 7103
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9876 6458 9904 6598
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9784 5370 9812 6326
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9954 6080 10010 6089
rect 9876 5642 9904 6054
rect 9954 6015 10010 6024
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9770 5264 9826 5273
rect 9770 5199 9826 5208
rect 9784 4185 9812 5199
rect 9876 4729 9904 5306
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9770 4176 9826 4185
rect 9770 4111 9826 4120
rect 9784 3942 9812 4111
rect 9968 4010 9996 6015
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9600 3590 9720 3618
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9600 2922 9628 3590
rect 9680 3528 9732 3534
rect 9772 3528 9824 3534
rect 9680 3470 9732 3476
rect 9770 3496 9772 3505
rect 9824 3496 9826 3505
rect 9692 2922 9720 3470
rect 9770 3431 9826 3440
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 10060 2514 10088 9823
rect 10152 7002 10180 10610
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8090 10272 8910
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10138 6760 10194 6769
rect 10138 6695 10194 6704
rect 10152 5273 10180 6695
rect 10138 5264 10194 5273
rect 10138 5199 10140 5208
rect 10192 5199 10194 5208
rect 10140 5170 10192 5176
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 3602 10180 4626
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10244 3233 10272 7822
rect 10336 7002 10364 10798
rect 10428 10198 10456 10950
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10520 10010 10548 11494
rect 10612 11393 10640 12582
rect 10598 11384 10654 11393
rect 10598 11319 10654 11328
rect 10612 11286 10640 11319
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10704 10674 10732 12974
rect 10874 12951 10930 12960
rect 10980 12850 11008 13670
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11164 12434 11192 15438
rect 11256 14618 11284 16458
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11348 13841 11376 16050
rect 11334 13832 11390 13841
rect 11334 13767 11390 13776
rect 11440 13530 11468 16186
rect 11532 15570 11560 16186
rect 11624 16046 11652 16594
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 15094 11560 15302
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 13734 11652 14962
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11072 12406 11192 12434
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11529 10916 12174
rect 10980 11762 11008 12242
rect 11072 12238 11100 12406
rect 11348 12306 11376 13466
rect 11518 13288 11574 13297
rect 11518 13223 11574 13232
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10874 11520 10930 11529
rect 10874 11455 10930 11464
rect 10782 10840 10838 10849
rect 10782 10775 10838 10784
rect 10796 10674 10824 10775
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 10033 10640 10542
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10062 10732 10406
rect 10692 10056 10744 10062
rect 10428 9982 10548 10010
rect 10598 10024 10654 10033
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10428 6225 10456 9982
rect 10692 9998 10744 10004
rect 10598 9959 10654 9968
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7206 10548 7822
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10690 6896 10746 6905
rect 10690 6831 10746 6840
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10414 6216 10470 6225
rect 10414 6151 10470 6160
rect 10520 5914 10548 6326
rect 10704 6254 10732 6831
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10416 5840 10468 5846
rect 10414 5808 10416 5817
rect 10468 5808 10470 5817
rect 10414 5743 10470 5752
rect 10704 5370 10732 6190
rect 10796 6118 10824 10610
rect 10888 10470 10916 11455
rect 11072 11286 11100 12174
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11440 11218 11468 12378
rect 11532 11762 11560 13223
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11518 11520 11574 11529
rect 11518 11455 11574 11464
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10606 11100 11086
rect 11426 10704 11482 10713
rect 11426 10639 11482 10648
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9382 10916 10202
rect 11072 10130 11100 10542
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10980 9897 11008 9930
rect 10966 9888 11022 9897
rect 10966 9823 11022 9832
rect 11072 9518 11100 10066
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10966 9072 11022 9081
rect 11072 9042 11100 9454
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10966 9007 10968 9016
rect 11020 9007 11022 9016
rect 11060 9036 11112 9042
rect 10968 8978 11020 8984
rect 11060 8978 11112 8984
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10888 6662 10916 7346
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5710 10916 5743
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10980 5370 11008 8366
rect 11072 7478 11100 8978
rect 11164 8906 11192 9386
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 6866 11100 7414
rect 11164 6866 11192 8298
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 11072 5817 11100 6151
rect 11058 5808 11114 5817
rect 11058 5743 11114 5752
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10336 5030 10364 5170
rect 10428 5137 10456 5170
rect 10414 5128 10470 5137
rect 10414 5063 10470 5072
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4486 10364 4966
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10324 4480 10376 4486
rect 10888 4457 10916 4490
rect 10324 4422 10376 4428
rect 10874 4448 10930 4457
rect 10336 4146 10364 4422
rect 10874 4383 10930 4392
rect 10980 4146 11008 5170
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10322 4040 10378 4049
rect 10322 3975 10378 3984
rect 10230 3224 10286 3233
rect 10230 3159 10286 3168
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 10336 800 10364 3975
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3466 10456 3878
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10980 1766 11008 4082
rect 11164 3466 11192 5238
rect 11256 4146 11284 9522
rect 11440 5914 11468 10639
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11532 5234 11560 11455
rect 11520 5228 11572 5234
rect 11348 5188 11520 5216
rect 11348 4622 11376 5188
rect 11520 5170 11572 5176
rect 11426 4992 11482 5001
rect 11426 4927 11482 4936
rect 11440 4758 11468 4927
rect 11428 4752 11480 4758
rect 11624 4706 11652 12242
rect 11716 9450 11744 17734
rect 11992 17678 12020 19887
rect 12360 19514 12388 20334
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 19922 12480 20198
rect 12544 19922 12572 20266
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12256 18760 12308 18766
rect 12254 18728 12256 18737
rect 12636 18737 12664 18770
rect 12308 18728 12310 18737
rect 12254 18663 12310 18672
rect 12622 18728 12678 18737
rect 12622 18663 12678 18672
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18358 12664 18566
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11808 16182 11836 16458
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15910 11836 15982
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11794 14512 11850 14521
rect 11794 14447 11850 14456
rect 11808 14414 11836 14447
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11900 12986 11928 17070
rect 11992 15910 12020 17614
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11992 15026 12020 15574
rect 12084 15502 12112 17818
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11978 14920 12034 14929
rect 11978 14855 12034 14864
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12306 12020 14855
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 14278 12112 14350
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12176 12986 12204 15302
rect 12360 15162 12388 18158
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17882 12480 18022
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 16250 12480 16458
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12544 16130 12572 16934
rect 12728 16658 12756 28018
rect 12820 17746 12848 31758
rect 13648 28218 13676 33934
rect 14556 33924 14608 33930
rect 14556 33866 14608 33872
rect 14568 28762 14596 33866
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 13636 28212 13688 28218
rect 13636 28154 13688 28160
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 12912 22098 12940 22510
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 13004 19378 13032 23598
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13464 23050 13584 23066
rect 13452 23044 13584 23050
rect 13504 23038 13584 23044
rect 13452 22986 13504 22992
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13096 22234 13124 22578
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 13188 21962 13216 22918
rect 13556 22642 13584 23038
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22409 13584 22578
rect 13542 22400 13598 22409
rect 13542 22335 13598 22344
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 13280 21706 13308 22034
rect 13188 21690 13308 21706
rect 13176 21684 13308 21690
rect 13228 21678 13308 21684
rect 13176 21626 13228 21632
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13096 17746 13124 21558
rect 13740 21010 13768 23462
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13832 20330 13860 28018
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13924 21622 13952 22374
rect 14016 22030 14044 23666
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 14016 21486 14044 21830
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19417 13584 19654
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13280 18630 13308 19110
rect 13464 18902 13492 19110
rect 13832 18902 13860 20266
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13924 18970 13952 19178
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13372 18222 13400 18634
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12820 17270 12848 17682
rect 12900 17604 12952 17610
rect 13464 17592 13492 18158
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 12900 17546 12952 17552
rect 13280 17564 13492 17592
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12452 16102 12572 16130
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12268 14278 12296 14554
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12360 13530 12388 14758
rect 12452 14414 12480 16102
rect 12636 15978 12664 16594
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12544 15434 12572 15846
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12452 14006 12480 14350
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12162 12744 12218 12753
rect 12452 12714 12480 13262
rect 12162 12679 12218 12688
rect 12440 12708 12492 12714
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11992 11898 12020 12106
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11558 11836 11630
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 12084 11354 12112 11834
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7342 11744 7754
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11702 6760 11758 6769
rect 11702 6695 11758 6704
rect 11428 4694 11480 4700
rect 11532 4678 11652 4706
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11532 4554 11560 4678
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 4214 11376 4422
rect 11532 4214 11560 4490
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11716 4078 11744 6695
rect 11808 6458 11836 11018
rect 11900 10538 11928 11154
rect 12176 11098 12204 12679
rect 12440 12650 12492 12656
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12256 12096 12308 12102
rect 12308 12056 12388 12084
rect 12256 12038 12308 12044
rect 12360 11506 12388 12056
rect 12452 11898 12480 12106
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12360 11478 12480 11506
rect 12452 11286 12480 11478
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12084 11070 12204 11098
rect 12346 11112 12402 11121
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 10130 11928 10474
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11886 9208 11942 9217
rect 11886 9143 11888 9152
rect 11940 9143 11942 9152
rect 11888 9114 11940 9120
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 5710 11836 6258
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11808 4146 11836 4626
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11532 2514 11560 3878
rect 11900 3126 11928 6666
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 6118 12020 6394
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5273 12020 5646
rect 11978 5264 12034 5273
rect 11978 5199 12034 5208
rect 11992 3670 12020 5199
rect 12084 4078 12112 11070
rect 12346 11047 12402 11056
rect 12162 10976 12218 10985
rect 12162 10911 12218 10920
rect 12176 8498 12204 10911
rect 12360 10742 12388 11047
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12346 9888 12402 9897
rect 12346 9823 12402 9832
rect 12360 9654 12388 9823
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12452 8634 12480 9046
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12452 7868 12480 8570
rect 12544 8566 12572 15370
rect 12728 14890 12756 15574
rect 12820 15162 12848 16118
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12714 14512 12770 14521
rect 12714 14447 12770 14456
rect 12728 13920 12756 14447
rect 12636 13892 12756 13920
rect 12636 12850 12664 13892
rect 12820 13818 12848 15098
rect 12912 14618 12940 17546
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13004 14498 13032 15982
rect 13096 15570 13124 16594
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 15706 13216 15982
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12912 14482 13032 14498
rect 12900 14476 13032 14482
rect 12952 14470 13032 14476
rect 12900 14418 12952 14424
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12728 13790 12848 13818
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12636 12442 12664 12786
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 11694 12756 13790
rect 12808 13728 12860 13734
rect 12912 13716 12940 13874
rect 12860 13688 12940 13716
rect 13188 13682 13216 14350
rect 12808 13670 12860 13676
rect 12820 12442 12848 13670
rect 13004 13654 13216 13682
rect 12898 13424 12954 13433
rect 12898 13359 12954 13368
rect 12912 13326 12940 13359
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12912 12102 12940 12650
rect 13004 12322 13032 13654
rect 13082 13560 13138 13569
rect 13082 13495 13138 13504
rect 13096 12481 13124 13495
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13082 12472 13138 12481
rect 13082 12407 13138 12416
rect 13004 12294 13124 12322
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12900 12096 12952 12102
rect 13004 12073 13032 12106
rect 12900 12038 12952 12044
rect 12990 12064 13046 12073
rect 12990 11999 13046 12008
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12714 10024 12770 10033
rect 12714 9959 12770 9968
rect 12728 9178 12756 9959
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12532 7880 12584 7886
rect 12162 7848 12218 7857
rect 12452 7840 12532 7868
rect 12532 7822 12584 7828
rect 12162 7783 12218 7792
rect 12624 7812 12676 7818
rect 12176 7750 12204 7783
rect 12624 7754 12676 7760
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12636 7546 12664 7754
rect 12728 7546 12756 9114
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12544 7274 12572 7414
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12346 7032 12402 7041
rect 12256 6996 12308 7002
rect 12346 6967 12402 6976
rect 12256 6938 12308 6944
rect 12268 6905 12296 6938
rect 12254 6896 12310 6905
rect 12360 6866 12388 6967
rect 12440 6928 12492 6934
rect 12438 6896 12440 6905
rect 12492 6896 12494 6905
rect 12254 6831 12310 6840
rect 12348 6860 12400 6866
rect 12438 6831 12494 6840
rect 12348 6802 12400 6808
rect 12256 6656 12308 6662
rect 12254 6624 12256 6633
rect 12716 6656 12768 6662
rect 12308 6624 12310 6633
rect 12254 6559 12310 6568
rect 12438 6624 12494 6633
rect 12716 6598 12768 6604
rect 12438 6559 12494 6568
rect 12452 6118 12480 6559
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12544 5778 12572 6190
rect 12622 5944 12678 5953
rect 12728 5914 12756 6598
rect 12622 5879 12678 5888
rect 12716 5908 12768 5914
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12162 5400 12218 5409
rect 12162 5335 12164 5344
rect 12216 5335 12218 5344
rect 12164 5306 12216 5312
rect 12438 5264 12494 5273
rect 12164 5228 12216 5234
rect 12438 5199 12494 5208
rect 12164 5170 12216 5176
rect 12176 4690 12204 5170
rect 12452 5166 12480 5199
rect 12544 5166 12572 5714
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12636 5030 12664 5879
rect 12716 5850 12768 5856
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12268 4434 12296 4490
rect 12176 4406 12296 4434
rect 12176 4282 12204 4406
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11992 3194 12020 3402
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11612 2848 11664 2854
rect 12084 2825 12112 4014
rect 12268 3602 12296 4218
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12360 3602 12388 4150
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12728 3534 12756 5510
rect 12820 5302 12848 10678
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8838 12940 9318
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8022 12940 8774
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12912 7002 12940 7346
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13004 6798 13032 8502
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12992 6792 13044 6798
rect 13096 6769 13124 12294
rect 13188 12170 13216 13194
rect 13280 13190 13308 17564
rect 13450 17504 13506 17513
rect 13450 17439 13506 17448
rect 13464 17202 13492 17439
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13832 16454 13860 17682
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13372 14618 13400 16390
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13372 13258 13400 14010
rect 13464 13569 13492 14826
rect 13450 13560 13506 13569
rect 13450 13495 13506 13504
rect 13648 13410 13676 14894
rect 13740 14006 13768 15302
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13464 13382 13676 13410
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13372 12434 13400 12582
rect 13280 12406 13400 12434
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9217 13216 10134
rect 13174 9208 13230 9217
rect 13174 9143 13230 9152
rect 13188 8974 13216 9143
rect 13280 9110 13308 12406
rect 13360 12232 13412 12238
rect 13358 12200 13360 12209
rect 13412 12200 13414 12209
rect 13358 12135 13414 12144
rect 13464 11121 13492 13382
rect 13740 12646 13768 13466
rect 13832 12850 13860 14486
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13450 11112 13506 11121
rect 13450 11047 13506 11056
rect 13450 10024 13506 10033
rect 13450 9959 13506 9968
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12992 6734 13044 6740
rect 13082 6760 13138 6769
rect 12912 6610 12940 6734
rect 13082 6695 13138 6704
rect 12912 6582 13032 6610
rect 12900 6384 12952 6390
rect 13004 6338 13032 6582
rect 12952 6332 13032 6338
rect 12900 6326 13032 6332
rect 12912 6310 13032 6326
rect 13004 5710 13032 6310
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12912 5234 12940 5510
rect 12992 5296 13044 5302
rect 12990 5264 12992 5273
rect 13044 5264 13046 5273
rect 12900 5228 12952 5234
rect 12990 5199 13046 5208
rect 12900 5170 12952 5176
rect 12912 3641 12940 5170
rect 12898 3632 12954 3641
rect 12898 3567 12954 3576
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 13188 3058 13216 8774
rect 13372 8566 13400 9318
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 4826 13308 7686
rect 13464 7290 13492 9959
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13372 7262 13492 7290
rect 13372 6254 13400 7262
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13464 5574 13492 7142
rect 13556 5710 13584 8910
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13648 4078 13676 12378
rect 13924 12306 13952 15506
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13938 14044 14214
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13726 11792 13782 11801
rect 13726 11727 13782 11736
rect 13740 10198 13768 11727
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13832 10538 13860 10950
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13924 10470 13952 10950
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 9450 13860 9590
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13728 8424 13780 8430
rect 13780 8401 13860 8412
rect 13780 8392 13874 8401
rect 13780 8384 13818 8392
rect 13728 8366 13780 8372
rect 13818 8327 13874 8336
rect 13728 8288 13780 8294
rect 13780 8236 13860 8242
rect 13728 8230 13860 8236
rect 13740 8214 13860 8230
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 7002 13768 7346
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6458 13768 6734
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13832 6390 13860 8214
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13924 5642 13952 10406
rect 14004 9648 14056 9654
rect 14002 9616 14004 9625
rect 14056 9616 14058 9625
rect 14002 9551 14058 9560
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 7585 14044 9454
rect 14108 9194 14136 23598
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 21690 14228 22374
rect 14292 22094 14320 22918
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14384 22545 14412 22578
rect 14370 22536 14426 22545
rect 14370 22471 14426 22480
rect 14476 22098 14504 23054
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14292 22066 14412 22094
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14292 19854 14320 21966
rect 14384 21010 14412 22066
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14568 21010 14596 22442
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 14372 21004 14424 21010
rect 14372 20946 14424 20952
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18154 14320 18566
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15706 14228 15982
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 13297 14228 15642
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14292 14890 14320 15574
rect 14384 15434 14412 15574
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14568 15026 14596 19790
rect 14660 18970 14688 20402
rect 14752 19922 14780 21014
rect 14936 20330 14964 22578
rect 15120 20466 15148 32710
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15304 23662 15332 25230
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15384 22024 15436 22030
rect 15488 22012 15516 24754
rect 15580 24206 15608 25842
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15580 23610 15608 24142
rect 15672 23730 15700 33254
rect 15948 32570 15976 36110
rect 16868 34746 16896 37198
rect 19996 37126 20024 39200
rect 21284 37262 21312 39200
rect 22572 37262 22600 39200
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 17132 37120 17184 37126
rect 17132 37062 17184 37068
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16856 29028 16908 29034
rect 16856 28970 16908 28976
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 23730 15884 24550
rect 15948 24274 15976 25094
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 15936 24268 15988 24274
rect 15936 24210 15988 24216
rect 16132 23730 16160 24550
rect 16316 24410 16344 24754
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16316 23866 16344 24142
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16028 23656 16080 23662
rect 15580 23582 15884 23610
rect 16028 23598 16080 23604
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15580 22098 15608 23462
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15436 21984 15516 22012
rect 15384 21966 15436 21972
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14648 18216 14700 18222
rect 14646 18184 14648 18193
rect 14700 18184 14702 18193
rect 14646 18119 14702 18128
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14648 16040 14700 16046
rect 14646 16008 14648 16017
rect 14700 16008 14702 16017
rect 14646 15943 14702 15952
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14292 14498 14320 14826
rect 14292 14470 14412 14498
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13938 14320 14350
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14186 13288 14242 13297
rect 14186 13223 14242 13232
rect 14186 13016 14242 13025
rect 14186 12951 14242 12960
rect 14200 12850 14228 12951
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14384 12646 14412 14470
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14476 12434 14504 14418
rect 14648 14408 14700 14414
rect 14646 14376 14648 14385
rect 14700 14376 14702 14385
rect 14646 14311 14702 14320
rect 14752 14278 14780 16526
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 12646 14780 12718
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14844 12434 14872 17002
rect 14384 12406 14504 12434
rect 14752 12406 14872 12434
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11830 14320 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14200 11150 14228 11766
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14200 10606 14228 11086
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 10044 14228 10542
rect 14280 10056 14332 10062
rect 14200 10016 14280 10044
rect 14280 9998 14332 10004
rect 14292 9518 14320 9998
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14108 9166 14228 9194
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14002 7576 14058 7585
rect 14002 7511 14058 7520
rect 14004 7472 14056 7478
rect 14002 7440 14004 7449
rect 14056 7440 14058 7449
rect 14002 7375 14058 7384
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6497 14044 6734
rect 14002 6488 14058 6497
rect 14002 6423 14058 6432
rect 14108 5930 14136 9046
rect 14200 6458 14228 9166
rect 14292 8974 14320 9454
rect 14384 9110 14412 12406
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 9926 14504 10542
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8294 14320 8910
rect 14476 8650 14504 9862
rect 14384 8622 14504 8650
rect 14384 8566 14412 8622
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14464 8424 14516 8430
rect 14370 8392 14426 8401
rect 14464 8366 14516 8372
rect 14370 8327 14426 8336
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7886 14320 8230
rect 14384 8106 14412 8327
rect 14476 8265 14504 8366
rect 14462 8256 14518 8265
rect 14462 8191 14518 8200
rect 14384 8078 14504 8106
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7002 14320 7822
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14016 5902 14136 5930
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 14016 5370 14044 5902
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14108 5302 14136 5782
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14200 4706 14228 6394
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14108 4678 14228 4706
rect 14292 4690 14320 5714
rect 14280 4684 14332 4690
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13542 3768 13598 3777
rect 13268 3732 13320 3738
rect 13542 3703 13598 3712
rect 13268 3674 13320 3680
rect 13280 3466 13308 3674
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12440 2848 12492 2854
rect 11612 2790 11664 2796
rect 12070 2816 12126 2825
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 11624 800 11652 2790
rect 12070 2751 12126 2760
rect 12438 2816 12440 2825
rect 12492 2816 12494 2825
rect 12438 2751 12494 2760
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 12084 1902 12112 2314
rect 13464 2281 13492 2586
rect 13450 2272 13506 2281
rect 13450 2207 13506 2216
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 13556 800 13584 3703
rect 13818 3360 13874 3369
rect 13818 3295 13874 3304
rect 13832 2990 13860 3295
rect 13820 2984 13872 2990
rect 13634 2952 13690 2961
rect 13820 2926 13872 2932
rect 13634 2887 13636 2896
rect 13688 2887 13690 2896
rect 13636 2858 13688 2864
rect 13924 2774 13952 4422
rect 14016 3602 14044 4626
rect 14108 4282 14136 4678
rect 14280 4626 14332 4632
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3670 14136 3878
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14016 3058 14044 3538
rect 14004 3052 14056 3058
rect 14056 3012 14136 3040
rect 14004 2994 14056 3000
rect 13924 2746 14044 2774
rect 14016 2650 14044 2746
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 2514 14136 3012
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14200 2378 14228 4558
rect 14278 3904 14334 3913
rect 14278 3839 14334 3848
rect 14292 3466 14320 3839
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14476 3097 14504 8078
rect 14568 6866 14596 12242
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 6866 14688 7754
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14568 5817 14596 6394
rect 14554 5808 14610 5817
rect 14554 5743 14610 5752
rect 14568 4690 14596 5743
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14462 3088 14518 3097
rect 14462 3023 14518 3032
rect 14752 2774 14780 12406
rect 14832 11008 14884 11014
rect 14936 10996 14964 20266
rect 15304 20058 15332 20334
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15488 19786 15516 21984
rect 15672 21554 15700 22374
rect 15764 21962 15792 22986
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15856 20346 15884 23582
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15948 21962 15976 22102
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15580 20318 15884 20346
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15212 19553 15240 19722
rect 15198 19544 15254 19553
rect 15198 19479 15254 19488
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 18902 15240 19246
rect 15488 18902 15516 19722
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15108 18760 15160 18766
rect 15580 18748 15608 20318
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15672 20058 15700 20198
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15764 19174 15792 20198
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15160 18720 15608 18748
rect 15108 18702 15160 18708
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15212 16726 15240 17070
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15028 14006 15056 16526
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12306 15056 13194
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14884 10968 14964 10996
rect 14832 10950 14884 10956
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14844 9897 14872 9930
rect 14830 9888 14886 9897
rect 14830 9823 14886 9832
rect 15120 9674 15148 16390
rect 15212 16250 15240 16662
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15304 14618 15332 17206
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 16046 15424 16458
rect 15488 16266 15516 18720
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17270 15608 17478
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15488 16238 15608 16266
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15094 15424 15982
rect 15474 15872 15530 15881
rect 15474 15807 15530 15816
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15488 15026 15516 15807
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15396 14521 15424 14894
rect 15382 14512 15438 14521
rect 15382 14447 15438 14456
rect 15488 14414 15516 14962
rect 15580 14482 15608 16238
rect 15764 15314 15792 18838
rect 15856 18766 15884 19654
rect 15948 19514 15976 20878
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15948 15638 15976 19110
rect 16040 18426 16068 23598
rect 16500 23526 16528 24006
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16592 23322 16620 24686
rect 16776 24410 16804 28494
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16684 23186 16712 23530
rect 16776 23322 16804 24346
rect 16868 23662 16896 28970
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16868 23186 16896 23598
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16316 21894 16344 22578
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16132 18970 16160 20878
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16500 20534 16528 20810
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16210 19952 16266 19961
rect 16210 19887 16212 19896
rect 16264 19887 16266 19896
rect 16212 19858 16264 19864
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16132 17134 16160 18226
rect 16224 17678 16252 18566
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16316 17202 16344 19790
rect 16396 18828 16448 18834
rect 16448 18788 16528 18816
rect 16396 18770 16448 18776
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15672 15286 15792 15314
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 13320 15344 13326
rect 15290 13288 15292 13297
rect 15344 13288 15346 13297
rect 15290 13223 15346 13232
rect 15396 12714 15424 13806
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12986 15516 13262
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 14832 9648 14884 9654
rect 15120 9646 15332 9674
rect 14832 9590 14884 9596
rect 14844 6361 14872 9590
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14830 6352 14886 6361
rect 14936 6322 14964 6666
rect 14830 6287 14886 6296
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15028 5234 15056 7890
rect 15304 7426 15332 9646
rect 15396 8106 15424 12310
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 10606 15516 11494
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15580 10538 15608 12038
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15672 10033 15700 15286
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 13864 15896 13870
rect 15948 13841 15976 14350
rect 15844 13806 15896 13812
rect 15934 13832 15990 13841
rect 15856 13462 15884 13806
rect 15934 13767 15990 13776
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15856 12850 15884 13398
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15948 12442 15976 13194
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15856 11801 15884 12174
rect 15842 11792 15898 11801
rect 15842 11727 15844 11736
rect 15896 11727 15898 11736
rect 15844 11698 15896 11704
rect 15856 11667 15884 11698
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15764 11286 15792 11317
rect 15752 11280 15804 11286
rect 15750 11248 15752 11257
rect 15804 11248 15806 11257
rect 15750 11183 15806 11192
rect 15658 10024 15714 10033
rect 15658 9959 15714 9968
rect 15474 9888 15530 9897
rect 15474 9823 15530 9832
rect 15488 8430 15516 9823
rect 15764 9674 15792 11183
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10810 15884 11018
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15764 9646 15884 9674
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 8294 15516 8366
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15396 8078 15516 8106
rect 15382 7440 15438 7449
rect 15304 7398 15382 7426
rect 15382 7375 15438 7384
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15120 5370 15148 6870
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14844 4486 14872 5034
rect 15198 4720 15254 4729
rect 15198 4655 15254 4664
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14476 2746 14780 2774
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14108 2038 14136 2314
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 14476 1970 14504 2746
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14844 800 14872 3334
rect 15212 2961 15240 4655
rect 15396 4010 15424 7375
rect 15488 4486 15516 8078
rect 15580 5914 15608 8434
rect 15764 8401 15792 9454
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 15750 7576 15806 7585
rect 15750 7511 15806 7520
rect 15764 7342 15792 7511
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6390 15792 7142
rect 15856 7041 15884 9646
rect 15842 7032 15898 7041
rect 15842 6967 15898 6976
rect 15856 6730 15884 6967
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15948 6390 15976 11494
rect 16040 9518 16068 14894
rect 16132 12306 16160 16934
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14074 16252 15438
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 11014 16160 11562
rect 16210 11384 16266 11393
rect 16210 11319 16266 11328
rect 16224 11218 16252 11319
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16120 11008 16172 11014
rect 16212 11008 16264 11014
rect 16120 10950 16172 10956
rect 16210 10976 16212 10985
rect 16264 10976 16266 10985
rect 16132 10810 16160 10950
rect 16210 10911 16266 10920
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16224 9926 16252 10474
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16132 9330 16160 9590
rect 16040 9302 16160 9330
rect 16040 7750 16068 9302
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16132 7750 16160 9114
rect 16224 8294 16252 9862
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16316 8090 16344 16730
rect 16408 11558 16436 18090
rect 16500 13394 16528 18788
rect 16684 18698 16712 22102
rect 16776 21622 16804 22646
rect 16960 22094 16988 32370
rect 17052 28762 17080 34546
rect 17144 32910 17172 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20088 33658 20116 37198
rect 20352 37188 20404 37194
rect 20352 37130 20404 37136
rect 23388 37188 23440 37194
rect 23388 37130 23440 37136
rect 20076 33652 20128 33658
rect 20076 33594 20128 33600
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 18052 32224 18104 32230
rect 18052 32166 18104 32172
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17144 23254 17172 23598
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16868 22066 16988 22094
rect 16868 22030 16896 22066
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 20913 16804 21286
rect 16762 20904 16818 20913
rect 16762 20839 16818 20848
rect 16960 20380 16988 22066
rect 17052 21622 17080 22374
rect 17328 22234 17356 23054
rect 17420 22930 17448 28426
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24206 17540 24550
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17604 23050 17632 25230
rect 17696 24274 17724 25638
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 17420 22902 17632 22930
rect 17406 22672 17462 22681
rect 17406 22607 17408 22616
rect 17460 22607 17462 22616
rect 17408 22578 17460 22584
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17052 20806 17080 21082
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17040 20392 17092 20398
rect 16960 20352 17040 20380
rect 17040 20334 17092 20340
rect 17144 20058 17172 21966
rect 17222 20904 17278 20913
rect 17222 20839 17224 20848
rect 17276 20839 17278 20848
rect 17224 20810 17276 20816
rect 17420 20618 17448 22374
rect 17604 21622 17632 22902
rect 17696 22574 17724 23122
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17788 22438 17816 24686
rect 17972 24682 18000 25842
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 18064 23730 18092 32166
rect 19248 30864 19300 30870
rect 19248 30806 19300 30812
rect 18972 25696 19024 25702
rect 18972 25638 19024 25644
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17880 22681 17908 23190
rect 18248 23186 18276 25094
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18340 22778 18368 24754
rect 18616 24274 18644 25094
rect 18984 24818 19012 25638
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19168 24410 19196 24550
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18708 23322 18736 24074
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 19260 23066 19288 30806
rect 19444 27606 19472 33458
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20364 32434 20392 37130
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20456 32502 20484 37062
rect 23020 34604 23072 34610
rect 23020 34546 23072 34552
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 20444 32496 20496 32502
rect 20444 32438 20496 32444
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 30592 20036 30598
rect 19984 30534 20036 30540
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 23798 19380 25094
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19444 23254 19472 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19628 24138 19656 24618
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19168 23038 19288 23066
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 17866 22672 17922 22681
rect 17866 22607 17922 22616
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 18248 22098 18276 22442
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18064 21690 18092 21966
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18156 21690 18184 21898
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17604 21010 17632 21558
rect 18432 21486 18460 22374
rect 19168 22094 19196 23038
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 22438 19288 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22574 20024 30534
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19536 22166 19564 22510
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 20088 22094 20116 27406
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20364 24274 20392 24550
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 20180 23866 20208 24074
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20456 22094 20484 32166
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20640 22574 20668 24686
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20732 22234 20760 24142
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 19168 22066 19288 22094
rect 20088 22066 20208 22094
rect 19260 21554 19288 22066
rect 19984 22024 20036 22030
rect 19982 21992 19984 22001
rect 20036 21992 20038 22001
rect 19982 21927 20038 21936
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17592 20868 17644 20874
rect 17592 20810 17644 20816
rect 17236 20590 17448 20618
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16854 19408 16910 19417
rect 17236 19394 17264 20590
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 16854 19343 16856 19352
rect 16908 19343 16910 19352
rect 16960 19366 17264 19394
rect 16856 19314 16908 19320
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16592 16590 16620 17546
rect 16868 17338 16896 18702
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16960 17218 16988 19366
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16868 17190 16988 17218
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 15162 16620 16050
rect 16684 15706 16712 16186
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16408 11150 16436 11222
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16486 10160 16542 10169
rect 16486 10095 16542 10104
rect 16500 10062 16528 10095
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16592 9518 16620 14554
rect 16776 13190 16804 16594
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16868 12434 16896 17190
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 16182 16988 16526
rect 17052 16250 17080 18158
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16960 12986 16988 15302
rect 17052 14618 17080 15982
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17144 14550 17172 18634
rect 17236 17882 17264 19246
rect 17328 18970 17356 20470
rect 17604 19922 17632 20810
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17696 19378 17724 20266
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17604 18902 17632 19178
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17236 14362 17264 16730
rect 17420 16726 17448 18090
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15638 17540 15914
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 14414 17448 14758
rect 17052 14334 17264 14362
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17052 13870 17080 14334
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12986 17080 13262
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12850 17172 13738
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16868 12406 16988 12434
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16684 11937 16712 12242
rect 16670 11928 16726 11937
rect 16670 11863 16726 11872
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16408 8974 16436 9114
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16132 6254 16160 6598
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15672 5409 15700 6190
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15658 5400 15714 5409
rect 15658 5335 15714 5344
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3369 15516 3878
rect 15474 3360 15530 3369
rect 15474 3295 15530 3304
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15384 3052 15436 3058
rect 15672 3040 15700 3130
rect 15436 3012 15700 3040
rect 15384 2994 15436 3000
rect 15198 2952 15254 2961
rect 15198 2887 15254 2896
rect 15856 2774 15884 5782
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 4010 15976 5510
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16026 4856 16082 4865
rect 16026 4791 16028 4800
rect 16080 4791 16082 4800
rect 16028 4762 16080 4768
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15934 3768 15990 3777
rect 15934 3703 15990 3712
rect 15948 3670 15976 3703
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15936 3392 15988 3398
rect 16040 3380 16068 4762
rect 15988 3352 16068 3380
rect 15936 3334 15988 3340
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15856 2746 15976 2774
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15580 1698 15608 2314
rect 15948 1902 15976 2746
rect 16040 2689 16068 2926
rect 16026 2680 16082 2689
rect 16026 2615 16028 2624
rect 16080 2615 16082 2624
rect 16028 2586 16080 2592
rect 16040 2555 16068 2586
rect 16132 2553 16160 5170
rect 16224 3398 16252 6734
rect 16316 5642 16344 8026
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16408 4826 16436 8366
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16500 7206 16528 7414
rect 16592 7410 16620 8910
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16500 6322 16528 6870
rect 16578 6760 16634 6769
rect 16578 6695 16580 6704
rect 16632 6695 16634 6704
rect 16580 6666 16632 6672
rect 16684 6497 16712 9998
rect 16776 9058 16804 11154
rect 16868 10742 16896 11290
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16868 9722 16896 10134
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16776 9030 16896 9058
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8022 16804 8910
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16868 6934 16896 9030
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16500 5914 16528 6258
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16488 5772 16540 5778
rect 16684 5760 16712 6258
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16540 5732 16712 5760
rect 16488 5714 16540 5720
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 3670 16528 4966
rect 16684 4690 16712 4966
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16776 4554 16804 6054
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16486 3496 16542 3505
rect 16486 3431 16488 3440
rect 16540 3431 16542 3440
rect 16488 3402 16540 3408
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16118 2544 16174 2553
rect 16118 2479 16174 2488
rect 16592 2446 16620 3674
rect 16868 3602 16896 5102
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16776 3194 16804 3402
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16868 3058 16896 3538
rect 16960 3466 16988 12406
rect 17052 12102 17080 12582
rect 17236 12442 17264 13806
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13462 17448 13670
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17144 11898 17172 12174
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17236 11778 17264 12106
rect 17144 11750 17264 11778
rect 17328 11762 17356 12106
rect 17316 11756 17368 11762
rect 17144 10606 17172 11750
rect 17316 11698 17368 11704
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 8634 17080 9998
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17052 8022 17080 8230
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 17052 5370 17080 7754
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17144 4146 17172 10542
rect 17236 10130 17264 10542
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17328 9994 17356 10678
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17236 8378 17264 8774
rect 17328 8498 17356 8774
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17236 8362 17356 8378
rect 17236 8356 17368 8362
rect 17236 8350 17316 8356
rect 17316 8298 17368 8304
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17236 4146 17264 6938
rect 17328 6866 17356 8298
rect 17420 7954 17448 13398
rect 17512 12434 17540 15574
rect 17604 15434 17632 18838
rect 17696 16250 17724 19314
rect 17972 18698 18000 19382
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 17610 17908 18022
rect 17972 17678 18000 18634
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17788 14618 17816 17070
rect 17972 16998 18000 17478
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17604 13394 17632 13874
rect 17972 13870 18000 16594
rect 18064 15978 18092 17750
rect 18248 16658 18276 19654
rect 18340 19174 18368 21082
rect 18800 20942 18828 21490
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18290 18368 19110
rect 18432 18426 18460 19790
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 18340 14618 18368 16458
rect 18432 14958 18460 18022
rect 18524 16561 18552 20878
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18616 20482 18644 20538
rect 18880 20528 18932 20534
rect 18616 20476 18880 20482
rect 18616 20470 18932 20476
rect 18616 20454 18920 20470
rect 19260 19922 19288 21490
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19444 21146 19472 21422
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18708 19514 18736 19722
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18984 18970 19012 19314
rect 19260 19310 19288 19858
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 19352 18850 19380 20266
rect 19444 20058 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20534 20024 21014
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 20088 20262 20116 21898
rect 20180 20330 20208 22066
rect 20364 22066 20484 22094
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19260 18822 19380 18850
rect 19444 18834 19472 19790
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19432 18828 19484 18834
rect 19260 18358 19288 18822
rect 19432 18770 19484 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18616 16658 18644 17002
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18510 16552 18566 16561
rect 18510 16487 18566 16496
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18064 13938 18092 14350
rect 18432 14074 18460 14350
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17512 12406 17632 12434
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17512 8906 17540 11018
rect 17604 9926 17632 12406
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11150 17724 12038
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17788 10996 17816 12718
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17696 10968 17816 10996
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17512 7177 17540 8298
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17498 7168 17554 7177
rect 17498 7103 17554 7112
rect 17406 7032 17462 7041
rect 17406 6967 17408 6976
rect 17460 6967 17462 6976
rect 17408 6938 17460 6944
rect 17604 6934 17632 7754
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17696 6866 17724 10968
rect 17880 10130 17908 11018
rect 17972 11014 18000 13806
rect 18064 13705 18092 13874
rect 18050 13696 18106 13705
rect 18050 13631 18106 13640
rect 18326 13424 18382 13433
rect 18326 13359 18382 13368
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12714 18092 13126
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 7585 17816 9658
rect 17774 7576 17830 7585
rect 17774 7511 17830 7520
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17880 4690 17908 9862
rect 17972 9382 18000 10066
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 5953 18000 8230
rect 18064 7954 18092 12650
rect 18248 12442 18276 12718
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 11898 18184 12174
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 11762 18276 11834
rect 18340 11762 18368 13359
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18524 11529 18552 12786
rect 18616 11762 18644 16594
rect 18800 16046 18828 17070
rect 18892 16726 18920 18158
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18984 15706 19012 17070
rect 19352 16522 19380 18702
rect 19536 18612 19564 19246
rect 19444 18584 19564 18612
rect 19444 17882 19472 18584
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 19994
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20272 18358 20300 18906
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20364 18204 20392 22066
rect 20824 21332 20852 24754
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20916 23798 20944 24006
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 21100 23186 21128 24550
rect 22020 23730 22048 24754
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21272 23248 21324 23254
rect 21272 23190 21324 23196
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21284 22982 21312 23190
rect 22112 23050 22140 23462
rect 22204 23186 22232 33254
rect 23032 29306 23060 34546
rect 23400 33522 23428 37130
rect 24504 37126 24532 39200
rect 25792 37262 25820 39200
rect 27724 37262 27752 39200
rect 29012 37262 29040 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 29000 37256 29052 37262
rect 30300 37244 30328 39200
rect 32232 37262 32260 39200
rect 33520 37262 33548 39200
rect 34808 37262 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36740 37262 36768 39200
rect 37186 38176 37242 38185
rect 37186 38111 37242 38120
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 29000 37198 29052 37204
rect 30380 37198 30432 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33968 37256 34020 37262
rect 33968 37198 34020 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24596 34746 24624 37198
rect 29644 37188 29696 37194
rect 29644 37130 29696 37136
rect 32588 37188 32640 37194
rect 32588 37130 32640 37136
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 24860 36848 24912 36854
rect 24860 36790 24912 36796
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 24872 33522 24900 36790
rect 23388 33516 23440 33522
rect 23388 33458 23440 33464
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 23020 29300 23072 29306
rect 23020 29242 23072 29248
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22388 23186 22416 24074
rect 22572 23798 22600 29106
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24780 23866 24808 26930
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22572 23118 22600 23734
rect 24964 23322 24992 33254
rect 27632 30938 27660 37062
rect 29276 36576 29328 36582
rect 29276 36518 29328 36524
rect 28264 32768 28316 32774
rect 28264 32710 28316 32716
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 25964 30592 26016 30598
rect 25964 30534 26016 30540
rect 27804 30592 27856 30598
rect 27804 30534 27856 30540
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21284 22778 21312 22918
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21376 21962 21404 22646
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 20904 21344 20956 21350
rect 20824 21304 20904 21332
rect 20824 21010 20852 21304
rect 20904 21286 20956 21292
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20602 20760 20878
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 21008 20398 21036 21014
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 20466 21128 20878
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 19922 20944 20198
rect 21008 20058 21036 20334
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 19706 18184 19762 18193
rect 19706 18119 19762 18128
rect 19812 18176 20392 18204
rect 19720 18086 19748 18119
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19444 17338 19472 17682
rect 19812 17678 19840 18176
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20272 17338 20300 17614
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 15162 18920 15438
rect 19352 15162 19380 15506
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18800 12986 18828 15030
rect 19444 14074 19472 16118
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19628 14482 19656 14894
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13326 19472 13874
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18892 12850 18920 13262
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19076 12434 19104 13262
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 18708 12406 19104 12434
rect 19996 12434 20024 15982
rect 20088 14618 20116 17206
rect 20456 17134 20484 19314
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20640 18426 20668 18634
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20824 18358 20852 18770
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20640 16726 20668 17138
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 20364 16250 20392 16458
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 14618 20208 15438
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 12986 20208 13262
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19996 12406 20116 12434
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18510 11520 18566 11529
rect 18510 11455 18566 11464
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18248 10690 18276 11086
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18156 10662 18276 10690
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18156 7834 18184 10662
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8566 18276 9318
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18064 7806 18184 7834
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 17958 5944 18014 5953
rect 17958 5879 18014 5888
rect 18064 5778 18092 7806
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7410 18184 7686
rect 18248 7546 18276 7822
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18340 7342 18368 10406
rect 18432 9722 18460 10950
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 10169 18552 10406
rect 18510 10160 18566 10169
rect 18510 10095 18566 10104
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18616 9178 18644 10542
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18420 8560 18472 8566
rect 18418 8528 18420 8537
rect 18472 8528 18474 8537
rect 18418 8463 18474 8472
rect 18418 8256 18474 8265
rect 18418 8191 18474 8200
rect 18432 8106 18460 8191
rect 18708 8106 18736 12406
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19892 11824 19944 11830
rect 19944 11772 20024 11778
rect 19892 11766 20024 11772
rect 19904 11750 20024 11766
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 8650 18828 11494
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 10532 18932 10538
rect 18880 10474 18932 10480
rect 18892 10130 18920 10474
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18800 8622 18920 8650
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18432 8078 18736 8106
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 6866 18368 7278
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18142 6760 18198 6769
rect 18142 6695 18198 6704
rect 18156 6662 18184 6695
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18432 5914 18460 8078
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18616 7478 18644 7958
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 7478 18736 7686
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18524 4826 18552 6190
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18616 4826 18644 5102
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17236 3482 17264 3538
rect 17972 3534 18000 4490
rect 18064 4146 18092 4762
rect 18524 4468 18552 4762
rect 18524 4440 18644 4468
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 17052 3454 17264 3482
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18144 3460 18196 3466
rect 17052 3398 17080 3454
rect 18144 3402 18196 3408
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17144 3233 17172 3334
rect 17130 3224 17186 3233
rect 17130 3159 17186 3168
rect 17144 3126 17172 3159
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 18156 2774 18184 3402
rect 18512 3392 18564 3398
rect 18510 3360 18512 3369
rect 18564 3360 18566 3369
rect 18510 3295 18566 3304
rect 18064 2746 18184 2774
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 17868 2304 17920 2310
rect 17972 2281 18000 2314
rect 17868 2246 17920 2252
rect 17958 2272 18014 2281
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 15568 1692 15620 1698
rect 15568 1634 15620 1640
rect 16776 800 16804 2246
rect 17880 2106 17908 2246
rect 17958 2207 18014 2216
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 18064 800 18092 2746
rect 18616 2650 18644 4440
rect 18800 4010 18828 8230
rect 18892 5522 18920 8622
rect 18984 6662 19012 11222
rect 19444 10010 19472 11290
rect 19996 11150 20024 11750
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19536 10130 19564 10542
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19628 10010 19656 10066
rect 19352 9982 19656 10010
rect 19904 9994 19932 10678
rect 19892 9988 19944 9994
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19062 9072 19118 9081
rect 19062 9007 19064 9016
rect 19116 9007 19118 9016
rect 19064 8978 19116 8984
rect 19076 7936 19104 8978
rect 19260 8634 19288 9590
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8514 19380 9982
rect 19892 9930 19944 9936
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19444 9178 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19260 8486 19380 8514
rect 19890 8528 19946 8537
rect 19168 8294 19196 8434
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19260 8022 19288 8486
rect 19996 8498 20024 11086
rect 20088 9722 20116 12406
rect 20272 12238 20300 13874
rect 20364 12442 20392 15098
rect 20640 13938 20668 16662
rect 20732 15094 20760 16662
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20916 15162 20944 16118
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20824 13530 20852 14962
rect 20916 14074 20944 14962
rect 21008 14958 21036 16526
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 21100 14006 21128 20402
rect 21284 17814 21312 20470
rect 21272 17808 21324 17814
rect 21272 17750 21324 17756
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 16794 21312 17614
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21192 14414 21220 14894
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20456 12918 20484 13126
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20824 12850 20852 13126
rect 21192 12986 21220 14350
rect 21284 14074 21312 14350
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 21376 12782 21404 21898
rect 21468 21146 21496 21966
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21560 20534 21588 21898
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21652 17202 21680 22374
rect 21836 22234 21864 22578
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21928 21894 21956 22578
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21744 20874 21772 21082
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22112 19802 22140 20742
rect 22664 20398 22692 21286
rect 23124 20942 23152 21626
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22020 19786 22140 19802
rect 22008 19780 22140 19786
rect 22060 19774 22140 19780
rect 22008 19722 22060 19728
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22008 19304 22060 19310
rect 22204 19258 22232 19654
rect 22008 19246 22060 19252
rect 22020 18834 22048 19246
rect 22112 19242 22232 19258
rect 22100 19236 22232 19242
rect 22152 19230 22232 19236
rect 22100 19178 22152 19184
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22204 18290 22232 18702
rect 22664 18290 22692 20334
rect 23032 19854 23060 20402
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 23032 19174 23060 19790
rect 23216 19378 23244 20198
rect 23308 19514 23336 20198
rect 24952 19780 25004 19786
rect 24952 19722 25004 19728
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22112 18034 22140 18090
rect 22020 18006 22140 18034
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21744 16794 21772 17614
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 15910 21588 16390
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 13258 21496 13874
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20180 10577 20208 11766
rect 20166 10568 20222 10577
rect 20166 10503 20222 10512
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20088 9178 20116 9522
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19890 8463 19946 8472
rect 19984 8492 20036 8498
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 8016 19300 8022
rect 19352 7993 19380 8366
rect 19708 8016 19760 8022
rect 19248 7958 19300 7964
rect 19338 7984 19394 7993
rect 19076 7908 19196 7936
rect 19444 7966 19708 7970
rect 19338 7919 19394 7928
rect 19432 7964 19708 7966
rect 19432 7960 19760 7964
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18892 5494 19012 5522
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18892 4622 18920 5306
rect 18880 4616 18932 4622
rect 18984 4593 19012 5494
rect 19076 5370 19104 7754
rect 19168 7426 19196 7908
rect 19484 7958 19760 7960
rect 19484 7942 19748 7958
rect 19432 7902 19484 7908
rect 19340 7880 19392 7886
rect 19392 7840 19472 7868
rect 19340 7822 19392 7828
rect 19444 7834 19472 7840
rect 19444 7818 19656 7834
rect 19444 7812 19668 7818
rect 19444 7806 19616 7812
rect 19616 7754 19668 7760
rect 19340 7744 19392 7750
rect 19904 7732 19932 8463
rect 19984 8434 20036 8440
rect 20088 8412 20116 8910
rect 20180 8537 20208 10406
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20088 8384 20208 8412
rect 20074 8256 20130 8265
rect 20074 8191 20130 8200
rect 19904 7704 20024 7732
rect 19340 7686 19392 7692
rect 19352 7562 19380 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19352 7534 19472 7562
rect 19444 7449 19472 7534
rect 19616 7472 19668 7478
rect 19430 7440 19486 7449
rect 19168 7398 19288 7426
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19168 5914 19196 7278
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19260 5030 19288 7398
rect 19616 7414 19668 7420
rect 19430 7375 19486 7384
rect 19430 7304 19486 7313
rect 19628 7274 19656 7414
rect 19430 7239 19432 7248
rect 19484 7239 19486 7248
rect 19616 7268 19668 7274
rect 19432 7210 19484 7216
rect 19616 7210 19668 7216
rect 19430 7168 19486 7177
rect 19430 7103 19486 7112
rect 19444 6866 19472 7103
rect 19890 6896 19946 6905
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19524 6860 19576 6866
rect 19890 6831 19946 6840
rect 19524 6802 19576 6808
rect 19536 6746 19564 6802
rect 19904 6798 19932 6831
rect 19352 6718 19564 6746
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19352 5710 19380 6718
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6390 20024 7704
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 18880 4558 18932 4564
rect 18970 4584 19026 4593
rect 18970 4519 19026 4528
rect 19156 4480 19208 4486
rect 19062 4448 19118 4457
rect 19156 4422 19208 4428
rect 19062 4383 19118 4392
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18708 2746 19012 2774
rect 18708 2650 18736 2746
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 18892 2446 18920 2479
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18984 1902 19012 2746
rect 19076 2650 19104 4383
rect 19168 2854 19196 4422
rect 19352 3913 19380 5646
rect 19444 5370 19472 6326
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19904 5846 19932 6258
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19720 5030 19748 5170
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4146 20024 5646
rect 20088 4486 20116 8191
rect 20180 7313 20208 8384
rect 20272 8265 20300 11834
rect 20640 11762 20668 12582
rect 21192 12238 21220 12582
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21192 11898 21220 12174
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21836 11830 21864 17614
rect 22020 16726 22048 18006
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 22204 15910 22232 18226
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22112 15162 22140 15438
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20718 11656 20774 11665
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 10674 20392 11494
rect 20456 11218 20484 11630
rect 20718 11591 20774 11600
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20548 11354 20576 11494
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20548 10810 20576 11086
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20350 10568 20406 10577
rect 20350 10503 20406 10512
rect 20364 9178 20392 10503
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20258 8256 20314 8265
rect 20258 8191 20314 8200
rect 20456 8106 20484 9658
rect 20272 8078 20484 8106
rect 20536 8084 20588 8090
rect 20166 7304 20222 7313
rect 20166 7239 20222 7248
rect 20272 6866 20300 8078
rect 20536 8026 20588 8032
rect 20548 7868 20576 8026
rect 20364 7840 20576 7868
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20166 6760 20222 6769
rect 20166 6695 20168 6704
rect 20220 6695 20222 6704
rect 20168 6666 20220 6672
rect 20260 6656 20312 6662
rect 20258 6624 20260 6633
rect 20312 6624 20314 6633
rect 20258 6559 20314 6568
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19338 3904 19394 3913
rect 19338 3839 19394 3848
rect 20088 3641 20116 4082
rect 19522 3632 19578 3641
rect 19522 3567 19578 3576
rect 20074 3632 20130 3641
rect 20074 3567 20130 3576
rect 19536 3534 19564 3567
rect 20180 3534 20208 4558
rect 20272 3738 20300 6394
rect 20364 5914 20392 7840
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20456 7546 20484 7686
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 4146 20392 5510
rect 20456 5370 20484 7142
rect 20548 6304 20576 7686
rect 20640 6662 20668 10678
rect 20732 8974 20760 11591
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21008 10674 21036 11222
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21008 10130 21036 10406
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9722 20852 9998
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20902 9480 20958 9489
rect 20902 9415 20958 9424
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20718 8528 20774 8537
rect 20718 8463 20774 8472
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20628 6316 20680 6322
rect 20548 6276 20628 6304
rect 20628 6258 20680 6264
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20548 5234 20576 5646
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20640 4758 20668 6258
rect 20732 5574 20760 8463
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7954 20852 8230
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20916 7342 20944 9415
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20996 7268 21048 7274
rect 20996 7210 21048 7216
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 5642 20852 7142
rect 21008 6934 21036 7210
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 21192 6798 21220 7346
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 20904 6656 20956 6662
rect 20902 6624 20904 6633
rect 20956 6624 20958 6633
rect 20902 6559 20958 6568
rect 21192 6322 21220 6734
rect 21284 6458 21312 8327
rect 21468 8090 21496 9862
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21376 6905 21404 7754
rect 21468 7478 21496 8026
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21362 6896 21418 6905
rect 21362 6831 21418 6840
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20916 5642 20944 6122
rect 21086 5944 21142 5953
rect 21086 5879 21142 5888
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 21100 5574 21128 5879
rect 21192 5710 21220 6258
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 20732 4570 20760 5306
rect 21284 5234 21312 6054
rect 21376 5778 21404 6598
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 20640 4542 20760 4570
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20258 3632 20314 3641
rect 20364 3618 20392 3674
rect 20314 3590 20392 3618
rect 20258 3567 20314 3576
rect 19524 3528 19576 3534
rect 19444 3488 19524 3516
rect 19444 3058 19472 3488
rect 19524 3470 19576 3476
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19430 2952 19486 2961
rect 19340 2916 19392 2922
rect 20088 2938 20116 3334
rect 20180 3058 20208 3470
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19430 2887 19432 2896
rect 19340 2858 19392 2864
rect 19484 2887 19486 2896
rect 19616 2916 19668 2922
rect 19432 2858 19484 2864
rect 20088 2910 20208 2938
rect 19616 2858 19668 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19352 2774 19380 2858
rect 19628 2774 19656 2858
rect 20180 2854 20208 2910
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19260 2746 19380 2774
rect 19444 2746 19656 2774
rect 19260 2666 19288 2746
rect 19064 2644 19116 2650
rect 19260 2638 19380 2666
rect 19064 2586 19116 2592
rect 19352 2582 19380 2638
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 18972 1896 19024 1902
rect 18972 1838 19024 1844
rect 19352 800 19380 2246
rect 19444 2106 19472 2746
rect 20272 2446 20300 3567
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20456 3194 20484 3402
rect 20548 3194 20576 4014
rect 20640 3505 20668 4542
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 3534 20760 4014
rect 21008 3534 21036 4082
rect 21100 3942 21128 4966
rect 21468 4826 21496 6258
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21284 4010 21312 4558
rect 21560 4010 21588 6190
rect 21652 5030 21680 9046
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 21836 8090 21864 8502
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21928 7886 21956 12038
rect 22020 11898 22048 13942
rect 22204 13938 22232 14214
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22480 13530 22508 14486
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22480 13274 22508 13466
rect 22296 13246 22508 13274
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22204 11354 22232 12854
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22112 10742 22140 11018
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 22112 9178 22140 10678
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22204 10062 22232 10202
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21836 6798 21864 7278
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21916 6656 21968 6662
rect 21836 6604 21916 6610
rect 21836 6598 21968 6604
rect 21836 6582 21956 6598
rect 21836 5166 21864 6582
rect 22008 5568 22060 5574
rect 21928 5516 22008 5522
rect 21928 5510 22060 5516
rect 21928 5494 22048 5510
rect 21928 5302 21956 5494
rect 22204 5302 22232 9590
rect 22296 7546 22324 13246
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22480 11898 22508 12038
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22572 11286 22600 15302
rect 22664 14929 22692 18226
rect 23308 18193 23336 18226
rect 23294 18184 23350 18193
rect 23294 18119 23350 18128
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23400 17882 23428 18022
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 22756 17202 22784 17478
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23124 16658 23152 17070
rect 23308 16794 23336 17070
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22650 14920 22706 14929
rect 22650 14855 22706 14864
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22664 13530 22692 13670
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22848 13462 22876 16050
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23124 15570 23152 15982
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15570 23336 15846
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 23032 13394 23060 13670
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23124 13326 23152 13806
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 23216 13326 23244 13738
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22388 9586 22416 9998
rect 22480 9654 22508 11086
rect 22756 11082 22784 12038
rect 22940 11694 22968 12106
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 23032 10266 23060 11766
rect 23216 10266 23244 12582
rect 23308 12306 23336 13466
rect 23400 12782 23428 16934
rect 23492 16590 23520 17478
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 24872 16182 24900 16594
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23584 14822 23612 15302
rect 24044 15026 24072 15982
rect 24136 15706 24164 16050
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24872 15026 24900 15302
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23492 12442 23520 12718
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23492 11098 23520 12378
rect 23584 12306 23612 14758
rect 24412 14618 24440 14758
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24216 14544 24268 14550
rect 24216 14486 24268 14492
rect 24228 14006 24256 14486
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24412 13870 24440 14554
rect 24596 14482 24624 14758
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24412 13258 24440 13466
rect 24400 13252 24452 13258
rect 24400 13194 24452 13200
rect 24504 12918 24532 14350
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24688 12850 24716 13194
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24032 12708 24084 12714
rect 24032 12650 24084 12656
rect 24044 12434 24072 12650
rect 24688 12434 24716 12786
rect 23952 12406 24072 12434
rect 24412 12406 24716 12434
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23400 11070 23520 11098
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23308 10198 23336 10950
rect 23400 10674 23428 11070
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23112 10192 23164 10198
rect 23112 10134 23164 10140
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 23124 9994 23152 10134
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 23112 9988 23164 9994
rect 23112 9930 23164 9936
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22848 8974 22876 9930
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22376 8900 22428 8906
rect 22376 8842 22428 8848
rect 22388 7886 22416 8842
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22480 6866 22508 8910
rect 23216 8634 23244 9590
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23308 8634 23336 9454
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22572 6458 22600 8366
rect 22926 7440 22982 7449
rect 22926 7375 22928 7384
rect 22980 7375 22982 7384
rect 22928 7346 22980 7352
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22664 6798 22692 6938
rect 23124 6798 23152 7142
rect 23400 6798 23428 10474
rect 23492 10062 23520 10950
rect 23570 10296 23626 10305
rect 23570 10231 23626 10240
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23492 9178 23520 9454
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 23112 6792 23164 6798
rect 23388 6792 23440 6798
rect 23112 6734 23164 6740
rect 23294 6760 23350 6769
rect 23388 6734 23440 6740
rect 23294 6695 23350 6704
rect 23308 6662 23336 6695
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22572 5914 22600 6394
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 23020 5704 23072 5710
rect 23072 5664 23152 5692
rect 23020 5646 23072 5652
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21928 5030 21956 5102
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 22020 4622 22048 5170
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20720 3528 20772 3534
rect 20626 3496 20682 3505
rect 20720 3470 20772 3476
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20626 3431 20682 3440
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 21008 3058 21036 3470
rect 21192 3126 21220 3878
rect 21560 3602 21588 3946
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21180 3120 21232 3126
rect 21180 3062 21232 3068
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 20916 1970 20944 2246
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 21284 800 21312 2926
rect 21928 1698 21956 4422
rect 22020 3534 22048 4558
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22020 3194 22048 3470
rect 22112 3466 22140 4966
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 4214 22600 4422
rect 22756 4282 22784 4966
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 23020 4140 23072 4146
rect 23124 4128 23152 5664
rect 23216 4729 23244 6598
rect 23492 6322 23520 8774
rect 23584 7426 23612 10231
rect 23676 7970 23704 11630
rect 23768 10810 23796 12038
rect 23952 11694 23980 12406
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23848 11620 23900 11626
rect 23848 11562 23900 11568
rect 23860 11286 23888 11562
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 23952 9926 23980 10610
rect 24044 10062 24072 10610
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23860 8090 23888 8366
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23676 7942 23888 7970
rect 23584 7398 23796 7426
rect 23572 7336 23624 7342
rect 23624 7296 23704 7324
rect 23572 7278 23624 7284
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23294 5264 23350 5273
rect 23294 5199 23350 5208
rect 23202 4720 23258 4729
rect 23202 4655 23258 4664
rect 23308 4146 23336 5199
rect 23492 5166 23520 5646
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23400 4214 23428 4762
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23204 4140 23256 4146
rect 23124 4100 23204 4128
rect 23020 4082 23072 4088
rect 23204 4082 23256 4088
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22020 3058 22048 3130
rect 22100 3120 22152 3126
rect 22152 3068 22232 3074
rect 22100 3062 22232 3068
rect 22008 3052 22060 3058
rect 22112 3046 22232 3062
rect 22296 3058 22324 3606
rect 23032 3534 23060 4082
rect 23216 3670 23244 4082
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 3058 23060 3470
rect 23400 3058 23428 4150
rect 23492 3738 23520 5102
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 22008 2994 22060 3000
rect 22020 2446 22048 2994
rect 22204 2990 22232 3046
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22836 2984 22888 2990
rect 22888 2932 23152 2938
rect 22836 2926 23152 2932
rect 22848 2910 23152 2926
rect 23124 2854 23152 2910
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23584 2446 23612 3606
rect 23676 2650 23704 7296
rect 23768 5914 23796 7398
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23768 4214 23796 5170
rect 23860 4758 23888 7942
rect 23952 7206 23980 9318
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23952 5098 23980 7142
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23848 4752 23900 4758
rect 23848 4694 23900 4700
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23952 4282 23980 4558
rect 23940 4276 23992 4282
rect 23940 4218 23992 4224
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23768 4078 23796 4150
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23768 2446 23796 4014
rect 22008 2440 22060 2446
rect 23572 2440 23624 2446
rect 22008 2382 22060 2388
rect 23478 2408 23534 2417
rect 22284 2372 22336 2378
rect 23572 2382 23624 2388
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23478 2343 23534 2352
rect 22284 2314 22336 2320
rect 22296 1766 22324 2314
rect 23492 2310 23520 2343
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 22284 1760 22336 1766
rect 22284 1702 22336 1708
rect 21916 1692 21968 1698
rect 21916 1634 21968 1640
rect 22572 800 22600 2246
rect 23860 800 23888 2246
rect 24044 1902 24072 6734
rect 24136 5370 24164 10542
rect 24228 10266 24256 12174
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24320 8498 24348 11562
rect 24412 9518 24440 12406
rect 24492 12368 24544 12374
rect 24780 12322 24808 13806
rect 24964 13394 24992 19722
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25148 15026 25176 15438
rect 25424 15162 25452 15438
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25148 13530 25176 14962
rect 25516 13938 25544 20878
rect 25976 18902 26004 30534
rect 27816 24750 27844 30534
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 28276 22098 28304 32710
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29012 28218 29040 31758
rect 29288 30258 29316 36518
rect 29656 30666 29684 37130
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 29748 36854 29776 37062
rect 29736 36848 29788 36854
rect 29736 36790 29788 36796
rect 29840 30870 29868 37062
rect 32416 33046 32444 37062
rect 32404 33040 32456 33046
rect 32404 32982 32456 32988
rect 31116 32768 31168 32774
rect 31116 32710 31168 32716
rect 31852 32768 31904 32774
rect 31852 32710 31904 32716
rect 29828 30864 29880 30870
rect 29828 30806 29880 30812
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29276 30252 29328 30258
rect 29276 30194 29328 30200
rect 29368 30048 29420 30054
rect 29368 29990 29420 29996
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 28264 22092 28316 22098
rect 28264 22034 28316 22040
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 25964 18896 26016 18902
rect 25964 18838 26016 18844
rect 27632 17814 27660 19654
rect 28920 18834 28948 28018
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25884 14414 25912 14554
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 25792 13326 25820 13466
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24492 12310 24544 12316
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24412 7546 24440 9454
rect 24504 8974 24532 12310
rect 24688 12294 24808 12322
rect 24688 11626 24716 12294
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24780 11354 24808 12174
rect 24872 11694 24900 12582
rect 25240 11898 25268 12718
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24596 8634 24624 9454
rect 24780 9110 24808 11086
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24688 8022 24716 8910
rect 24964 8634 24992 11834
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 25056 10810 25084 11630
rect 25332 11354 25360 11766
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25516 11286 25544 12786
rect 25884 12434 25912 14350
rect 26068 14278 26096 14962
rect 29380 14822 29408 29990
rect 31128 24342 31156 32710
rect 31760 30728 31812 30734
rect 31760 30670 31812 30676
rect 31772 27130 31800 30670
rect 31760 27124 31812 27130
rect 31760 27066 31812 27072
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31116 24336 31168 24342
rect 31116 24278 31168 24284
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30392 22030 30420 24142
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 31772 21622 31800 25094
rect 31760 21616 31812 21622
rect 31760 21558 31812 21564
rect 31864 19446 31892 32710
rect 32220 31816 32272 31822
rect 32220 31758 32272 31764
rect 32232 19990 32260 31758
rect 32600 30802 32628 37130
rect 33876 35080 33928 35086
rect 33876 35022 33928 35028
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 32588 30796 32640 30802
rect 32588 30738 32640 30744
rect 33244 27470 33272 32166
rect 33888 30938 33916 35022
rect 33980 32026 34008 37198
rect 35348 37120 35400 37126
rect 35348 37062 35400 37068
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 32978 35388 37062
rect 37200 36174 37228 38111
rect 38028 36786 38056 39200
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 38212 36825 38240 37062
rect 39316 36854 39344 39200
rect 39304 36848 39356 36854
rect 38198 36816 38254 36825
rect 38016 36780 38068 36786
rect 39304 36790 39356 36796
rect 38198 36751 38254 36760
rect 38016 36722 38068 36728
rect 38108 36576 38160 36582
rect 38108 36518 38160 36524
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 35900 36032 35952 36038
rect 35900 35974 35952 35980
rect 35348 32972 35400 32978
rect 35348 32914 35400 32920
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 33968 32020 34020 32026
rect 33968 31962 34020 31968
rect 35912 31890 35940 35974
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 35900 31884 35952 31890
rect 35900 31826 35952 31832
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33508 27464 33560 27470
rect 33508 27406 33560 27412
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 32404 25152 32456 25158
rect 32404 25094 32456 25100
rect 32220 19984 32272 19990
rect 32220 19926 32272 19932
rect 32416 19922 32444 25094
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33152 20806 33180 22578
rect 33140 20800 33192 20806
rect 33140 20742 33192 20748
rect 32404 19916 32456 19922
rect 32404 19858 32456 19864
rect 31852 19440 31904 19446
rect 31852 19382 31904 19388
rect 33336 15638 33364 27270
rect 33520 24410 33548 27406
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36556 25362 36584 29990
rect 36544 25356 36596 25362
rect 36544 25298 36596 25304
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33508 24404 33560 24410
rect 33508 24346 33560 24352
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 36924 22778 36952 25230
rect 37004 24064 37056 24070
rect 37004 24006 37056 24012
rect 36912 22772 36964 22778
rect 36912 22714 36964 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 33600 20936 33652 20942
rect 33600 20878 33652 20884
rect 33612 18970 33640 20878
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 37016 19854 37044 24006
rect 37004 19848 37056 19854
rect 37004 19790 37056 19796
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 33428 18426 33456 18702
rect 33416 18420 33468 18426
rect 33416 18362 33468 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34532 16454 34560 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 37004 15904 37056 15910
rect 37004 15846 37056 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33324 15632 33376 15638
rect 33324 15574 33376 15580
rect 37016 15026 37044 15846
rect 37004 15020 37056 15026
rect 37004 14962 37056 14968
rect 29368 14816 29420 14822
rect 29368 14758 29420 14764
rect 33140 14816 33192 14822
rect 33140 14758 33192 14764
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 25792 12406 25912 12434
rect 25504 11280 25556 11286
rect 25504 11222 25556 11228
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 25240 9625 25268 11086
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25332 10266 25360 10542
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25226 9616 25282 9625
rect 25516 9586 25544 11222
rect 25792 11218 25820 12406
rect 26068 11762 26096 14214
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26620 13326 26648 14010
rect 33152 13802 33180 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 33140 13796 33192 13802
rect 33140 13738 33192 13744
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 36464 12986 36492 14350
rect 37844 14346 37872 33458
rect 38120 32910 38148 36518
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 32065 38332 32370
rect 38290 32056 38346 32065
rect 38290 31991 38346 32000
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 38304 30025 38332 30194
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38108 29028 38160 29034
rect 38108 28970 38160 28976
rect 38120 25430 38148 28970
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38108 25424 38160 25430
rect 38108 25366 38160 25372
rect 38198 25256 38254 25265
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 38108 21956 38160 21962
rect 38108 21898 38160 21904
rect 37924 21888 37976 21894
rect 38120 21865 38148 21898
rect 37924 21830 37976 21836
rect 38106 21856 38162 21865
rect 37832 14340 37884 14346
rect 37832 14282 37884 14288
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25884 11150 25912 11494
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 26068 10062 26096 11698
rect 29104 11354 29132 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 29092 11348 29144 11354
rect 29092 11290 29144 11296
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 28908 11076 28960 11082
rect 28908 11018 28960 11024
rect 28920 10062 28948 11018
rect 33692 10532 33744 10538
rect 33692 10474 33744 10480
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 25226 9551 25282 9560
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25516 9466 25544 9522
rect 25424 9438 25544 9466
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 25424 7886 25452 9438
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 25516 8566 25544 9318
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24504 7002 24532 7686
rect 24688 7342 24716 7686
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 26516 7268 26568 7274
rect 26516 7210 26568 7216
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 24492 5296 24544 5302
rect 24492 5238 24544 5244
rect 24504 4282 24532 5238
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24596 3534 24624 6326
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24688 2446 24716 6054
rect 24780 4826 24808 6190
rect 26528 5234 26556 7210
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 27620 4752 27672 4758
rect 27620 4694 27672 4700
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3126 24808 3334
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 25240 2038 25268 3878
rect 27632 3534 27660 4694
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25792 3097 25820 3130
rect 25778 3088 25834 3097
rect 25778 3023 25834 3032
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27540 2582 27568 2926
rect 29748 2650 29776 8434
rect 30208 5710 30236 9318
rect 33704 8634 33732 10474
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 36096 10266 36124 11086
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 35072 10056 35124 10062
rect 35072 9998 35124 10004
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 8974 34836 9862
rect 35084 9654 35112 9998
rect 35072 9648 35124 9654
rect 35072 9590 35124 9596
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34716 8090 34744 8434
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 31944 7336 31996 7342
rect 31944 7278 31996 7284
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 30300 2582 30328 6734
rect 31956 4826 31984 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 33048 5568 33100 5574
rect 33048 5510 33100 5516
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 31944 4820 31996 4826
rect 31944 4762 31996 4768
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 32324 2446 32352 4966
rect 33060 2514 33088 5510
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35820 4826 35848 7346
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 35808 4820 35860 4826
rect 35808 4762 35860 4768
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 33600 4548 33652 4554
rect 33600 4490 33652 4496
rect 33612 2650 33640 4490
rect 33888 3738 33916 4558
rect 36372 4010 36400 6734
rect 37738 6352 37794 6361
rect 37738 6287 37740 6296
rect 37792 6287 37794 6296
rect 37740 6258 37792 6264
rect 37464 6248 37516 6254
rect 37462 6216 37464 6225
rect 37516 6216 37518 6225
rect 37462 6151 37518 6160
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 36360 4004 36412 4010
rect 36360 3946 36412 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 36912 3392 36964 3398
rect 36912 3334 36964 3340
rect 36924 3058 36952 3334
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25228 2032 25280 2038
rect 25228 1974 25280 1980
rect 24032 1896 24084 1902
rect 24032 1838 24084 1844
rect 25792 800 25820 2246
rect 27080 800 27108 2382
rect 29012 800 29040 2382
rect 30300 800 30328 2382
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 800 31616 2246
rect 33520 800 33548 2382
rect 34808 800 34836 2382
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 36096 800 36124 2246
rect 37200 1465 37228 4082
rect 37936 3466 37964 21830
rect 38106 21791 38162 21800
rect 38200 20800 38252 20806
rect 38200 20742 38252 20748
rect 38212 20505 38240 20742
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 38304 15745 38332 16050
rect 38290 15736 38346 15745
rect 38290 15671 38346 15680
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38028 12442 38056 12786
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38016 12436 38068 12442
rect 38016 12378 38068 12384
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38200 11280 38252 11286
rect 38200 11222 38252 11228
rect 38212 10985 38240 11222
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38028 5234 38056 6598
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 37924 3460 37976 3466
rect 37924 3402 37976 3408
rect 38028 3058 38056 4966
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4185 38332 4558
rect 38290 4176 38346 4185
rect 38290 4111 38346 4120
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 38028 2446 38056 2790
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38120 1986 38148 3470
rect 38200 2848 38252 2854
rect 38198 2816 38200 2825
rect 38252 2816 38254 2825
rect 38198 2751 38254 2760
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 38028 1958 38148 1986
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 38028 800 38056 1958
rect 39316 800 39344 2246
rect 4632 734 5028 762
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 2778 38120 2834 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1766 36780 1822 36816
rect 1766 36760 1768 36780
rect 1768 36760 1820 36780
rect 1820 36760 1822 36780
rect 1766 33380 1822 33416
rect 1766 33360 1768 33380
rect 1768 33360 1820 33380
rect 1820 33360 1822 33380
rect 1766 32000 1822 32056
rect 1766 30676 1768 30696
rect 1768 30676 1820 30696
rect 1820 30676 1822 30696
rect 1766 30640 1822 30676
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 1766 28600 1822 28656
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1766 25236 1768 25256
rect 1768 25236 1820 25256
rect 1820 25236 1822 25256
rect 1766 25200 1822 25236
rect 1766 23840 1822 23896
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 1766 22480 1822 22536
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1766 20440 1822 20496
rect 1766 19080 1822 19136
rect 1766 17720 1822 17776
rect 1766 15680 1822 15736
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 1582 13932 1638 13968
rect 1582 13912 1584 13932
rect 1584 13912 1636 13932
rect 1636 13912 1638 13932
rect 1766 12280 1822 12336
rect 1398 7520 1454 7576
rect 1766 10920 1822 10976
rect 1766 9560 1822 9616
rect 1306 4800 1362 4856
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1398 2760 1454 2816
rect 3054 13812 3056 13832
rect 3056 13812 3108 13832
rect 3108 13812 3110 13832
rect 3054 13776 3110 13812
rect 3054 8608 3110 8664
rect 2870 8356 2926 8392
rect 2870 8336 2872 8356
rect 2872 8336 2924 8356
rect 2924 8336 2926 8356
rect 2962 6704 3018 6760
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12552 4122 12608
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4618 12416 4674 12472
rect 3054 4700 3056 4720
rect 3056 4700 3108 4720
rect 3108 4700 3110 4720
rect 3054 4664 3110 4700
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4250 10784 4306 10840
rect 4618 10784 4674 10840
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4526 8356 4582 8392
rect 4526 8336 4528 8356
rect 4528 8336 4580 8356
rect 4580 8336 4582 8356
rect 3790 6296 3846 6352
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3460 4306 3496
rect 4250 3440 4252 3460
rect 4252 3440 4304 3460
rect 4304 3440 4306 3460
rect 6918 17856 6974 17912
rect 4986 8336 5042 8392
rect 4986 8200 5042 8256
rect 5170 13096 5226 13152
rect 5446 11736 5502 11792
rect 5354 10240 5410 10296
rect 5722 10684 5724 10704
rect 5724 10684 5776 10704
rect 5776 10684 5778 10704
rect 5722 10648 5778 10684
rect 5998 12552 6054 12608
rect 6090 10376 6146 10432
rect 5998 9460 6000 9480
rect 6000 9460 6052 9480
rect 6052 9460 6054 9480
rect 5998 9424 6054 9460
rect 5446 4564 5448 4584
rect 5448 4564 5500 4584
rect 5500 4564 5502 4584
rect 5446 4528 5502 4564
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4710 2488 4766 2544
rect 2778 1400 2834 1456
rect 5906 6316 5962 6352
rect 5906 6296 5908 6316
rect 5908 6296 5960 6316
rect 5960 6296 5962 6316
rect 6274 11464 6330 11520
rect 6458 12008 6514 12064
rect 6550 9052 6552 9072
rect 6552 9052 6604 9072
rect 6604 9052 6606 9072
rect 6550 9016 6606 9052
rect 6274 6740 6276 6760
rect 6276 6740 6328 6760
rect 6328 6740 6330 6760
rect 6274 6704 6330 6740
rect 6366 6196 6368 6216
rect 6368 6196 6420 6216
rect 6420 6196 6422 6216
rect 6366 6160 6422 6196
rect 7010 12144 7066 12200
rect 7010 11872 7066 11928
rect 7102 11076 7158 11112
rect 7102 11056 7104 11076
rect 7104 11056 7156 11076
rect 7156 11056 7158 11076
rect 7286 10920 7342 10976
rect 7654 13096 7710 13152
rect 7562 11872 7618 11928
rect 7470 11636 7472 11656
rect 7472 11636 7524 11656
rect 7524 11636 7526 11656
rect 7470 11600 7526 11636
rect 7470 11328 7526 11384
rect 7194 10104 7250 10160
rect 7562 10920 7618 10976
rect 6642 6432 6698 6488
rect 6550 5752 6606 5808
rect 6274 5480 6330 5536
rect 6918 6160 6974 6216
rect 6826 5072 6882 5128
rect 7194 5772 7250 5808
rect 7194 5752 7196 5772
rect 7196 5752 7248 5772
rect 7248 5752 7250 5772
rect 7194 5344 7250 5400
rect 9770 19488 9826 19544
rect 9862 19372 9918 19408
rect 9862 19352 9864 19372
rect 9864 19352 9916 19372
rect 9916 19352 9918 19372
rect 9310 18128 9366 18184
rect 9770 18148 9826 18184
rect 9770 18128 9772 18148
rect 9772 18128 9824 18148
rect 9824 18128 9826 18148
rect 10046 19660 10048 19680
rect 10048 19660 10100 19680
rect 10100 19660 10102 19680
rect 10046 19624 10102 19660
rect 8206 13776 8262 13832
rect 7838 5480 7894 5536
rect 7654 4276 7710 4312
rect 7654 4256 7656 4276
rect 7656 4256 7708 4276
rect 7708 4256 7710 4276
rect 8298 12300 8354 12336
rect 8298 12280 8300 12300
rect 8300 12280 8352 12300
rect 8352 12280 8354 12300
rect 9126 14320 9182 14376
rect 8666 13096 8722 13152
rect 8574 12436 8630 12472
rect 8574 12416 8576 12436
rect 8576 12416 8628 12436
rect 8628 12416 8630 12436
rect 8482 12144 8538 12200
rect 8666 11736 8722 11792
rect 8206 11192 8262 11248
rect 8758 11600 8814 11656
rect 8666 11056 8722 11112
rect 8574 10512 8630 10568
rect 8114 8472 8170 8528
rect 8850 9016 8906 9072
rect 9862 15816 9918 15872
rect 8206 5888 8262 5944
rect 8298 5752 8354 5808
rect 8206 5636 8262 5672
rect 8206 5616 8208 5636
rect 8208 5616 8260 5636
rect 8260 5616 8262 5636
rect 9310 12300 9366 12336
rect 9310 12280 9312 12300
rect 9312 12280 9364 12300
rect 9364 12280 9366 12300
rect 9770 13640 9826 13696
rect 9954 13388 10010 13424
rect 9954 13368 9956 13388
rect 9956 13368 10008 13388
rect 10008 13368 10010 13388
rect 9586 12688 9642 12744
rect 9494 11600 9550 11656
rect 9586 11056 9642 11112
rect 9586 10104 9642 10160
rect 8942 5752 8998 5808
rect 9034 5364 9090 5400
rect 9034 5344 9036 5364
rect 9036 5344 9088 5364
rect 9088 5344 9090 5364
rect 9402 8472 9458 8528
rect 9402 5752 9458 5808
rect 9494 5208 9550 5264
rect 10230 12144 10286 12200
rect 10230 11464 10286 11520
rect 10414 15972 10470 16008
rect 10414 15952 10416 15972
rect 10416 15952 10468 15972
rect 10468 15952 10470 15972
rect 11426 19352 11482 19408
rect 12070 20748 12072 20768
rect 12072 20748 12124 20768
rect 12124 20748 12126 20768
rect 12070 20712 12126 20748
rect 11978 19896 12034 19952
rect 11058 17484 11060 17504
rect 11060 17484 11112 17504
rect 11112 17484 11114 17504
rect 11058 17448 11114 17484
rect 10414 11872 10470 11928
rect 10046 9832 10102 9888
rect 9586 4276 9642 4312
rect 9586 4256 9588 4276
rect 9588 4256 9640 4276
rect 9640 4256 9642 4276
rect 9954 7112 10010 7168
rect 9954 6024 10010 6080
rect 9770 5208 9826 5264
rect 9862 4664 9918 4720
rect 9770 4120 9826 4176
rect 9770 3476 9772 3496
rect 9772 3476 9824 3496
rect 9824 3476 9826 3496
rect 9770 3440 9826 3476
rect 10138 6704 10194 6760
rect 10138 5228 10194 5264
rect 10138 5208 10140 5228
rect 10140 5208 10192 5228
rect 10192 5208 10194 5228
rect 10598 11328 10654 11384
rect 10874 12960 10930 13016
rect 11334 13776 11390 13832
rect 11518 13232 11574 13288
rect 10874 11464 10930 11520
rect 10782 10784 10838 10840
rect 10598 9968 10654 10024
rect 10690 6840 10746 6896
rect 10414 6160 10470 6216
rect 10414 5788 10416 5808
rect 10416 5788 10468 5808
rect 10468 5788 10470 5808
rect 10414 5752 10470 5788
rect 11518 11464 11574 11520
rect 11426 10648 11482 10704
rect 10966 9832 11022 9888
rect 10966 9036 11022 9072
rect 10966 9016 10968 9036
rect 10968 9016 11020 9036
rect 11020 9016 11022 9036
rect 10874 5752 10930 5808
rect 11058 6160 11114 6216
rect 11058 5752 11114 5808
rect 10414 5072 10470 5128
rect 10874 4392 10930 4448
rect 10322 3984 10378 4040
rect 10230 3168 10286 3224
rect 11426 4936 11482 4992
rect 12254 18708 12256 18728
rect 12256 18708 12308 18728
rect 12308 18708 12310 18728
rect 12254 18672 12310 18708
rect 12622 18672 12678 18728
rect 11794 14456 11850 14512
rect 11978 14864 12034 14920
rect 13542 22344 13598 22400
rect 13542 19352 13598 19408
rect 12162 12688 12218 12744
rect 11702 6704 11758 6760
rect 11886 9172 11942 9208
rect 11886 9152 11888 9172
rect 11888 9152 11940 9172
rect 11940 9152 11942 9172
rect 11978 5208 12034 5264
rect 12346 11056 12402 11112
rect 12162 10920 12218 10976
rect 12346 9832 12402 9888
rect 12714 14456 12770 14512
rect 12898 13368 12954 13424
rect 13082 13504 13138 13560
rect 13082 12416 13138 12472
rect 12990 12008 13046 12064
rect 12714 9968 12770 10024
rect 12162 7792 12218 7848
rect 12346 6976 12402 7032
rect 12254 6840 12310 6896
rect 12438 6876 12440 6896
rect 12440 6876 12492 6896
rect 12492 6876 12494 6896
rect 12438 6840 12494 6876
rect 12254 6604 12256 6624
rect 12256 6604 12308 6624
rect 12308 6604 12310 6624
rect 12254 6568 12310 6604
rect 12438 6568 12494 6624
rect 12622 5888 12678 5944
rect 12162 5364 12218 5400
rect 12162 5344 12164 5364
rect 12164 5344 12216 5364
rect 12216 5344 12218 5364
rect 12438 5208 12494 5264
rect 13450 17448 13506 17504
rect 13450 13504 13506 13560
rect 13174 9152 13230 9208
rect 13358 12180 13360 12200
rect 13360 12180 13412 12200
rect 13412 12180 13414 12200
rect 13358 12144 13414 12180
rect 13450 11056 13506 11112
rect 13450 9968 13506 10024
rect 13082 6704 13138 6760
rect 12990 5244 12992 5264
rect 12992 5244 13044 5264
rect 13044 5244 13046 5264
rect 12990 5208 13046 5244
rect 12898 3576 12954 3632
rect 13726 11736 13782 11792
rect 13818 8336 13874 8392
rect 14002 9596 14004 9616
rect 14004 9596 14056 9616
rect 14056 9596 14058 9616
rect 14002 9560 14058 9596
rect 14370 22480 14426 22536
rect 14646 18164 14648 18184
rect 14648 18164 14700 18184
rect 14700 18164 14702 18184
rect 14646 18128 14702 18164
rect 14646 15988 14648 16008
rect 14648 15988 14700 16008
rect 14700 15988 14702 16008
rect 14646 15952 14702 15988
rect 14186 13232 14242 13288
rect 14186 12960 14242 13016
rect 14646 14356 14648 14376
rect 14648 14356 14700 14376
rect 14700 14356 14702 14376
rect 14646 14320 14702 14356
rect 14002 7520 14058 7576
rect 14002 7420 14004 7440
rect 14004 7420 14056 7440
rect 14056 7420 14058 7440
rect 14002 7384 14058 7420
rect 14002 6432 14058 6488
rect 14370 8336 14426 8392
rect 14462 8200 14518 8256
rect 13542 3712 13598 3768
rect 12070 2760 12126 2816
rect 12438 2796 12440 2816
rect 12440 2796 12492 2816
rect 12492 2796 12494 2816
rect 12438 2760 12494 2796
rect 13450 2216 13506 2272
rect 13818 3304 13874 3360
rect 13634 2916 13690 2952
rect 13634 2896 13636 2916
rect 13636 2896 13688 2916
rect 13688 2896 13690 2916
rect 14278 3848 14334 3904
rect 14554 5752 14610 5808
rect 14462 3032 14518 3088
rect 15198 19488 15254 19544
rect 14830 9832 14886 9888
rect 15474 15816 15530 15872
rect 15382 14456 15438 14512
rect 16210 19916 16266 19952
rect 16210 19896 16212 19916
rect 16212 19896 16264 19916
rect 16264 19896 16266 19916
rect 15290 13268 15292 13288
rect 15292 13268 15344 13288
rect 15344 13268 15346 13288
rect 15290 13232 15346 13268
rect 14830 6296 14886 6352
rect 15934 13776 15990 13832
rect 15842 11756 15898 11792
rect 15842 11736 15844 11756
rect 15844 11736 15896 11756
rect 15896 11736 15898 11756
rect 15750 11228 15752 11248
rect 15752 11228 15804 11248
rect 15804 11228 15806 11248
rect 15750 11192 15806 11228
rect 15658 9968 15714 10024
rect 15474 9832 15530 9888
rect 15382 7384 15438 7440
rect 15198 4664 15254 4720
rect 15750 8336 15806 8392
rect 15750 7520 15806 7576
rect 15842 6976 15898 7032
rect 16210 11328 16266 11384
rect 16210 10956 16212 10976
rect 16212 10956 16264 10976
rect 16264 10956 16266 10976
rect 16210 10920 16266 10956
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 16762 20848 16818 20904
rect 17406 22636 17462 22672
rect 17406 22616 17408 22636
rect 17408 22616 17460 22636
rect 17460 22616 17462 22636
rect 17222 20868 17278 20904
rect 17222 20848 17224 20868
rect 17224 20848 17276 20868
rect 17276 20848 17278 20868
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 17866 22616 17922 22672
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19982 21972 19984 21992
rect 19984 21972 20036 21992
rect 20036 21972 20038 21992
rect 19982 21936 20038 21972
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 16854 19372 16910 19408
rect 16854 19352 16856 19372
rect 16856 19352 16908 19372
rect 16908 19352 16910 19372
rect 16486 10104 16542 10160
rect 16670 11872 16726 11928
rect 15658 5344 15714 5400
rect 15474 3304 15530 3360
rect 15198 2896 15254 2952
rect 16026 4820 16082 4856
rect 16026 4800 16028 4820
rect 16028 4800 16080 4820
rect 16080 4800 16082 4820
rect 15934 3712 15990 3768
rect 16026 2644 16082 2680
rect 16026 2624 16028 2644
rect 16028 2624 16080 2644
rect 16080 2624 16082 2644
rect 16578 6724 16634 6760
rect 16578 6704 16580 6724
rect 16580 6704 16632 6724
rect 16632 6704 16634 6724
rect 16670 6432 16726 6488
rect 16486 3460 16542 3496
rect 16486 3440 16488 3460
rect 16488 3440 16540 3460
rect 16540 3440 16542 3460
rect 16118 2488 16174 2544
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 18510 16496 18566 16552
rect 17498 7112 17554 7168
rect 17406 6996 17462 7032
rect 17406 6976 17408 6996
rect 17408 6976 17460 6996
rect 17460 6976 17462 6996
rect 18050 13640 18106 13696
rect 18326 13368 18382 13424
rect 17774 7520 17830 7576
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38120 37242 38176
rect 19706 18128 19762 18184
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 18510 11464 18566 11520
rect 17958 5888 18014 5944
rect 18510 10104 18566 10160
rect 18418 8508 18420 8528
rect 18420 8508 18472 8528
rect 18472 8508 18474 8528
rect 18418 8472 18474 8508
rect 18418 8200 18474 8256
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18142 6704 18198 6760
rect 17130 3168 17186 3224
rect 18510 3340 18512 3360
rect 18512 3340 18564 3360
rect 18564 3340 18566 3360
rect 18510 3304 18566 3340
rect 17958 2216 18014 2272
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19062 9036 19118 9072
rect 19062 9016 19064 9036
rect 19064 9016 19116 9036
rect 19116 9016 19118 9036
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19890 8472 19946 8528
rect 20166 10512 20222 10568
rect 19338 7928 19394 7984
rect 20166 8472 20222 8528
rect 20074 8200 20130 8256
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7384 19486 7440
rect 19430 7268 19486 7304
rect 19430 7248 19432 7268
rect 19432 7248 19484 7268
rect 19484 7248 19486 7268
rect 19430 7112 19486 7168
rect 19890 6840 19946 6896
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 18970 4528 19026 4584
rect 19062 4392 19118 4448
rect 18878 2488 18934 2544
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20718 11600 20774 11656
rect 20350 10512 20406 10568
rect 20258 8200 20314 8256
rect 20166 7248 20222 7304
rect 20166 6724 20222 6760
rect 20166 6704 20168 6724
rect 20168 6704 20220 6724
rect 20220 6704 20222 6724
rect 20258 6604 20260 6624
rect 20260 6604 20312 6624
rect 20312 6604 20314 6624
rect 20258 6568 20314 6604
rect 19338 3848 19394 3904
rect 19522 3576 19578 3632
rect 20074 3576 20130 3632
rect 20902 9424 20958 9480
rect 20718 8472 20774 8528
rect 21270 8336 21326 8392
rect 20902 6604 20904 6624
rect 20904 6604 20956 6624
rect 20956 6604 20958 6624
rect 20902 6568 20958 6604
rect 21362 6840 21418 6896
rect 21086 5888 21142 5944
rect 20258 3576 20314 3632
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19430 2916 19486 2952
rect 19430 2896 19432 2916
rect 19432 2896 19484 2916
rect 19484 2896 19486 2916
rect 23294 18128 23350 18184
rect 22650 14864 22706 14920
rect 22926 7404 22982 7440
rect 22926 7384 22928 7404
rect 22928 7384 22980 7404
rect 22980 7384 22982 7404
rect 23570 10240 23626 10296
rect 23294 6704 23350 6760
rect 20626 3440 20682 3496
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 23294 5208 23350 5264
rect 23202 4664 23258 4720
rect 23478 2352 23534 2408
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 38198 36760 38254 36816
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 25226 9560 25282 9616
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 38198 34720 38254 34776
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 32000 38346 32056
rect 38290 29960 38346 30016
rect 38290 28600 38346 28656
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38198 25200 38254 25256
rect 38290 23840 38346 23896
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 25778 3032 25834 3088
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37738 6316 37794 6352
rect 37738 6296 37740 6316
rect 37740 6296 37792 6316
rect 37792 6296 37794 6316
rect 37462 6196 37464 6216
rect 37464 6196 37516 6216
rect 37516 6196 37518 6216
rect 37462 6160 37518 6196
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38106 21800 38162 21856
rect 38198 20440 38254 20496
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 38290 15680 38346 15736
rect 38198 14320 38254 14376
rect 38198 12280 38254 12336
rect 38198 10920 38254 10976
rect 38198 8880 38254 8936
rect 38290 7520 38346 7576
rect 38290 4120 38346 4176
rect 38198 2796 38200 2816
rect 38200 2796 38252 2816
rect 38252 2796 38254 2816
rect 38198 2760 38254 2796
rect 37186 1400 37242 1456
<< metal3 >>
rect 200 38178 800 38208
rect 2773 38178 2839 38181
rect 200 38176 2839 38178
rect 200 38120 2778 38176
rect 2834 38120 2839 38176
rect 200 38118 2839 38120
rect 200 38088 800 38118
rect 2773 38115 2839 38118
rect 37181 38178 37247 38181
rect 39200 38178 39800 38208
rect 37181 38176 39800 38178
rect 37181 38120 37186 38176
rect 37242 38120 39800 38176
rect 37181 38118 39800 38120
rect 37181 38115 37247 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1761 36818 1827 36821
rect 200 36816 1827 36818
rect 200 36760 1766 36816
rect 1822 36760 1827 36816
rect 200 36758 1827 36760
rect 200 36728 800 36758
rect 1761 36755 1827 36758
rect 38193 36818 38259 36821
rect 39200 36818 39800 36848
rect 38193 36816 39800 36818
rect 38193 36760 38198 36816
rect 38254 36760 39800 36816
rect 38193 36758 39800 36760
rect 38193 36755 38259 36758
rect 39200 36728 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 9070 22612 9076 22676
rect 9140 22674 9146 22676
rect 17401 22674 17467 22677
rect 17861 22674 17927 22677
rect 9140 22672 17927 22674
rect 9140 22616 17406 22672
rect 17462 22616 17866 22672
rect 17922 22616 17927 22672
rect 9140 22614 17927 22616
rect 9140 22612 9146 22614
rect 17401 22611 17467 22614
rect 17861 22611 17927 22614
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 11278 22476 11284 22540
rect 11348 22538 11354 22540
rect 14365 22538 14431 22541
rect 11348 22536 14431 22538
rect 11348 22480 14370 22536
rect 14426 22480 14431 22536
rect 11348 22478 14431 22480
rect 11348 22476 11354 22478
rect 14365 22475 14431 22478
rect 13537 22402 13603 22405
rect 16062 22402 16068 22404
rect 13537 22400 16068 22402
rect 13537 22344 13542 22400
rect 13598 22344 16068 22400
rect 13537 22342 16068 22344
rect 13537 22339 13603 22342
rect 16062 22340 16068 22342
rect 16132 22340 16138 22404
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 17166 21932 17172 21996
rect 17236 21994 17242 21996
rect 19977 21994 20043 21997
rect 17236 21992 20043 21994
rect 17236 21936 19982 21992
rect 20038 21936 20043 21992
rect 17236 21934 20043 21936
rect 17236 21932 17242 21934
rect 19977 21931 20043 21934
rect 38101 21858 38167 21861
rect 39200 21858 39800 21888
rect 38101 21856 39800 21858
rect 38101 21800 38106 21856
rect 38162 21800 39800 21856
rect 38101 21798 39800 21800
rect 38101 21795 38167 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 16757 20906 16823 20909
rect 17217 20906 17283 20909
rect 16757 20904 17283 20906
rect 16757 20848 16762 20904
rect 16818 20848 17222 20904
rect 17278 20848 17283 20904
rect 16757 20846 17283 20848
rect 16757 20843 16823 20846
rect 17217 20843 17283 20846
rect 10910 20708 10916 20772
rect 10980 20770 10986 20772
rect 12065 20770 12131 20773
rect 10980 20768 12131 20770
rect 10980 20712 12070 20768
rect 12126 20712 12131 20768
rect 10980 20710 12131 20712
rect 10980 20708 10986 20710
rect 12065 20707 12131 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 11973 19954 12039 19957
rect 16205 19954 16271 19957
rect 11973 19952 16271 19954
rect 11973 19896 11978 19952
rect 12034 19896 16210 19952
rect 16266 19896 16271 19952
rect 11973 19894 16271 19896
rect 11973 19891 12039 19894
rect 16205 19891 16271 19894
rect 10041 19682 10107 19685
rect 10726 19682 10732 19684
rect 10041 19680 10732 19682
rect 10041 19624 10046 19680
rect 10102 19624 10732 19680
rect 10041 19622 10732 19624
rect 10041 19619 10107 19622
rect 10726 19620 10732 19622
rect 10796 19620 10802 19684
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 9765 19546 9831 19549
rect 15193 19546 15259 19549
rect 9765 19544 15259 19546
rect 9765 19488 9770 19544
rect 9826 19488 15198 19544
rect 15254 19488 15259 19544
rect 9765 19486 15259 19488
rect 9765 19483 9831 19486
rect 15193 19483 15259 19486
rect 9857 19410 9923 19413
rect 11421 19410 11487 19413
rect 9857 19408 11487 19410
rect 9857 19352 9862 19408
rect 9918 19352 11426 19408
rect 11482 19352 11487 19408
rect 9857 19350 11487 19352
rect 9857 19347 9923 19350
rect 11421 19347 11487 19350
rect 13537 19410 13603 19413
rect 16849 19410 16915 19413
rect 13537 19408 16915 19410
rect 13537 19352 13542 19408
rect 13598 19352 16854 19408
rect 16910 19352 16915 19408
rect 13537 19350 16915 19352
rect 13537 19347 13603 19350
rect 16849 19347 16915 19350
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19168
rect 34930 19007 35246 19008
rect 12249 18732 12315 18733
rect 12198 18730 12204 18732
rect 12122 18670 12204 18730
rect 12268 18730 12315 18732
rect 12617 18730 12683 18733
rect 12268 18728 12683 18730
rect 12310 18672 12622 18728
rect 12678 18672 12683 18728
rect 12198 18668 12204 18670
rect 12268 18670 12683 18672
rect 12268 18668 12315 18670
rect 12249 18667 12315 18668
rect 12617 18667 12683 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 7598 18124 7604 18188
rect 7668 18186 7674 18188
rect 9305 18186 9371 18189
rect 7668 18184 9371 18186
rect 7668 18128 9310 18184
rect 9366 18128 9371 18184
rect 7668 18126 9371 18128
rect 7668 18124 7674 18126
rect 9305 18123 9371 18126
rect 9765 18186 9831 18189
rect 14641 18186 14707 18189
rect 9765 18184 14707 18186
rect 9765 18128 9770 18184
rect 9826 18128 14646 18184
rect 14702 18128 14707 18184
rect 9765 18126 14707 18128
rect 9765 18123 9831 18126
rect 14641 18123 14707 18126
rect 19701 18186 19767 18189
rect 23289 18186 23355 18189
rect 19701 18184 23355 18186
rect 19701 18128 19706 18184
rect 19762 18128 23294 18184
rect 23350 18128 23355 18184
rect 19701 18126 23355 18128
rect 19701 18123 19767 18126
rect 23289 18123 23355 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 6678 17852 6684 17916
rect 6748 17914 6754 17916
rect 6913 17914 6979 17917
rect 6748 17912 6979 17914
rect 6748 17856 6918 17912
rect 6974 17856 6979 17912
rect 6748 17854 6979 17856
rect 6748 17852 6754 17854
rect 6913 17851 6979 17854
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 11053 17506 11119 17509
rect 13445 17506 13511 17509
rect 11053 17504 13511 17506
rect 11053 17448 11058 17504
rect 11114 17448 13450 17504
rect 13506 17448 13511 17504
rect 11053 17446 13511 17448
rect 11053 17443 11119 17446
rect 13445 17443 13511 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 16246 16492 16252 16556
rect 16316 16554 16322 16556
rect 18505 16554 18571 16557
rect 16316 16552 18571 16554
rect 16316 16496 18510 16552
rect 18566 16496 18571 16552
rect 16316 16494 18571 16496
rect 16316 16492 16322 16494
rect 18505 16491 18571 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 10409 16010 10475 16013
rect 14641 16010 14707 16013
rect 10409 16008 14707 16010
rect 10409 15952 10414 16008
rect 10470 15952 14646 16008
rect 14702 15952 14707 16008
rect 10409 15950 14707 15952
rect 10409 15947 10475 15950
rect 14641 15947 14707 15950
rect 9857 15874 9923 15877
rect 15469 15874 15535 15877
rect 9857 15872 15535 15874
rect 9857 15816 9862 15872
rect 9918 15816 15474 15872
rect 15530 15816 15535 15872
rect 9857 15814 15535 15816
rect 9857 15811 9923 15814
rect 15469 15811 15535 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 11973 14922 12039 14925
rect 22645 14922 22711 14925
rect 11973 14920 22711 14922
rect 11973 14864 11978 14920
rect 12034 14864 22650 14920
rect 22706 14864 22711 14920
rect 11973 14862 22711 14864
rect 11973 14859 12039 14862
rect 22645 14859 22711 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 11789 14514 11855 14517
rect 12709 14514 12775 14517
rect 15377 14514 15443 14517
rect 11789 14512 15443 14514
rect 11789 14456 11794 14512
rect 11850 14456 12714 14512
rect 12770 14456 15382 14512
rect 15438 14456 15443 14512
rect 11789 14454 15443 14456
rect 11789 14451 11855 14454
rect 12709 14451 12775 14454
rect 15377 14451 15443 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 9121 14378 9187 14381
rect 14641 14378 14707 14381
rect 9121 14376 14707 14378
rect 9121 14320 9126 14376
rect 9182 14320 14646 14376
rect 14702 14320 14707 14376
rect 9121 14318 14707 14320
rect 9121 14315 9187 14318
rect 14641 14315 14707 14318
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 1577 13970 1643 13973
rect 9622 13970 9628 13972
rect 1577 13968 9628 13970
rect 1577 13912 1582 13968
rect 1638 13912 9628 13968
rect 1577 13910 9628 13912
rect 1577 13907 1643 13910
rect 9622 13908 9628 13910
rect 9692 13908 9698 13972
rect 3049 13834 3115 13837
rect 3182 13834 3188 13836
rect 3049 13832 3188 13834
rect 3049 13776 3054 13832
rect 3110 13776 3188 13832
rect 3049 13774 3188 13776
rect 3049 13771 3115 13774
rect 3182 13772 3188 13774
rect 3252 13772 3258 13836
rect 8201 13834 8267 13837
rect 11329 13834 11395 13837
rect 15929 13834 15995 13837
rect 8201 13832 15995 13834
rect 8201 13776 8206 13832
rect 8262 13776 11334 13832
rect 11390 13776 15934 13832
rect 15990 13776 15995 13832
rect 8201 13774 15995 13776
rect 8201 13771 8267 13774
rect 11329 13771 11395 13774
rect 15929 13771 15995 13774
rect 9765 13698 9831 13701
rect 18045 13698 18111 13701
rect 9765 13696 18111 13698
rect 9765 13640 9770 13696
rect 9826 13640 18050 13696
rect 18106 13640 18111 13696
rect 9765 13638 18111 13640
rect 9765 13635 9831 13638
rect 18045 13635 18111 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 13077 13562 13143 13565
rect 13445 13562 13511 13565
rect 13077 13560 13511 13562
rect 13077 13504 13082 13560
rect 13138 13504 13450 13560
rect 13506 13504 13511 13560
rect 13077 13502 13511 13504
rect 13077 13499 13143 13502
rect 13445 13499 13511 13502
rect 9949 13426 10015 13429
rect 12893 13426 12959 13429
rect 18321 13426 18387 13429
rect 9949 13424 18387 13426
rect 9949 13368 9954 13424
rect 10010 13368 12898 13424
rect 12954 13368 18326 13424
rect 18382 13368 18387 13424
rect 9949 13366 18387 13368
rect 9949 13363 10015 13366
rect 12893 13363 12959 13366
rect 18321 13363 18387 13366
rect 11513 13290 11579 13293
rect 14181 13290 14247 13293
rect 15285 13290 15351 13293
rect 11513 13288 15351 13290
rect 11513 13232 11518 13288
rect 11574 13232 14186 13288
rect 14242 13232 15290 13288
rect 15346 13232 15351 13288
rect 11513 13230 15351 13232
rect 11513 13227 11579 13230
rect 14181 13227 14247 13230
rect 15285 13227 15351 13230
rect 5165 13154 5231 13157
rect 7649 13154 7715 13157
rect 8661 13154 8727 13157
rect 5165 13152 8727 13154
rect 5165 13096 5170 13152
rect 5226 13096 7654 13152
rect 7710 13096 8666 13152
rect 8722 13096 8727 13152
rect 5165 13094 8727 13096
rect 5165 13091 5231 13094
rect 7649 13091 7715 13094
rect 8661 13091 8727 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 10869 13018 10935 13021
rect 14181 13018 14247 13021
rect 10869 13016 14247 13018
rect 10869 12960 10874 13016
rect 10930 12960 14186 13016
rect 14242 12960 14247 13016
rect 10869 12958 14247 12960
rect 10869 12955 10935 12958
rect 14181 12955 14247 12958
rect 9581 12746 9647 12749
rect 12157 12746 12223 12749
rect 9581 12744 12223 12746
rect 9581 12688 9586 12744
rect 9642 12688 12162 12744
rect 12218 12688 12223 12744
rect 9581 12686 12223 12688
rect 9581 12683 9647 12686
rect 12157 12683 12223 12686
rect 3918 12548 3924 12612
rect 3988 12610 3994 12612
rect 4061 12610 4127 12613
rect 3988 12608 4127 12610
rect 3988 12552 4066 12608
rect 4122 12552 4127 12608
rect 3988 12550 4127 12552
rect 3988 12548 3994 12550
rect 4061 12547 4127 12550
rect 5993 12610 6059 12613
rect 6126 12610 6132 12612
rect 5993 12608 6132 12610
rect 5993 12552 5998 12608
rect 6054 12552 6132 12608
rect 5993 12550 6132 12552
rect 5993 12547 6059 12550
rect 6126 12548 6132 12550
rect 6196 12548 6202 12612
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4613 12474 4679 12477
rect 8569 12474 8635 12477
rect 4613 12472 8635 12474
rect 4613 12416 4618 12472
rect 4674 12416 8574 12472
rect 8630 12416 8635 12472
rect 4613 12414 8635 12416
rect 4613 12411 4679 12414
rect 8569 12411 8635 12414
rect 10542 12412 10548 12476
rect 10612 12474 10618 12476
rect 13077 12474 13143 12477
rect 10612 12472 13143 12474
rect 10612 12416 13082 12472
rect 13138 12416 13143 12472
rect 10612 12414 13143 12416
rect 10612 12412 10618 12414
rect 13077 12411 13143 12414
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 8293 12338 8359 12341
rect 9305 12338 9371 12341
rect 8293 12336 9371 12338
rect 8293 12280 8298 12336
rect 8354 12280 9310 12336
rect 9366 12280 9371 12336
rect 8293 12278 9371 12280
rect 8293 12275 8359 12278
rect 9305 12275 9371 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 7005 12202 7071 12205
rect 8477 12202 8543 12205
rect 7005 12200 8543 12202
rect 7005 12144 7010 12200
rect 7066 12144 8482 12200
rect 8538 12144 8543 12200
rect 7005 12142 8543 12144
rect 7005 12139 7071 12142
rect 8477 12139 8543 12142
rect 10225 12202 10291 12205
rect 13353 12202 13419 12205
rect 10225 12200 13419 12202
rect 10225 12144 10230 12200
rect 10286 12144 13358 12200
rect 13414 12144 13419 12200
rect 10225 12142 13419 12144
rect 10225 12139 10291 12142
rect 13353 12139 13419 12142
rect 6453 12066 6519 12069
rect 12985 12066 13051 12069
rect 6453 12064 13051 12066
rect 6453 12008 6458 12064
rect 6514 12008 12990 12064
rect 13046 12008 13051 12064
rect 6453 12006 13051 12008
rect 6453 12003 6519 12006
rect 12985 12003 13051 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 7005 11930 7071 11933
rect 7557 11930 7623 11933
rect 7005 11928 7623 11930
rect 7005 11872 7010 11928
rect 7066 11872 7562 11928
rect 7618 11872 7623 11928
rect 7005 11870 7623 11872
rect 7005 11867 7071 11870
rect 7557 11867 7623 11870
rect 10409 11930 10475 11933
rect 16665 11930 16731 11933
rect 10409 11928 16731 11930
rect 10409 11872 10414 11928
rect 10470 11872 16670 11928
rect 16726 11872 16731 11928
rect 10409 11870 16731 11872
rect 10409 11867 10475 11870
rect 16665 11867 16731 11870
rect 5441 11794 5507 11797
rect 8661 11794 8727 11797
rect 5441 11792 8727 11794
rect 5441 11736 5446 11792
rect 5502 11736 8666 11792
rect 8722 11736 8727 11792
rect 5441 11734 8727 11736
rect 5441 11731 5507 11734
rect 8661 11731 8727 11734
rect 13721 11794 13787 11797
rect 15837 11794 15903 11797
rect 13721 11792 15903 11794
rect 13721 11736 13726 11792
rect 13782 11736 15842 11792
rect 15898 11736 15903 11792
rect 13721 11734 15903 11736
rect 13721 11731 13787 11734
rect 15837 11731 15903 11734
rect 7465 11658 7531 11661
rect 8753 11658 8819 11661
rect 7465 11656 8819 11658
rect 7465 11600 7470 11656
rect 7526 11600 8758 11656
rect 8814 11600 8819 11656
rect 7465 11598 8819 11600
rect 7465 11595 7531 11598
rect 8753 11595 8819 11598
rect 9489 11658 9555 11661
rect 20713 11658 20779 11661
rect 9489 11656 20779 11658
rect 9489 11600 9494 11656
rect 9550 11600 20718 11656
rect 20774 11600 20779 11656
rect 9489 11598 20779 11600
rect 9489 11595 9555 11598
rect 20713 11595 20779 11598
rect 6269 11522 6335 11525
rect 10225 11522 10291 11525
rect 10869 11522 10935 11525
rect 6269 11520 10291 11522
rect 6269 11464 6274 11520
rect 6330 11464 10230 11520
rect 10286 11464 10291 11520
rect 6269 11462 10291 11464
rect 6269 11459 6335 11462
rect 10225 11459 10291 11462
rect 10366 11520 10935 11522
rect 10366 11464 10874 11520
rect 10930 11464 10935 11520
rect 10366 11462 10935 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 7465 11386 7531 11389
rect 10366 11386 10426 11462
rect 10869 11459 10935 11462
rect 11513 11522 11579 11525
rect 18505 11522 18571 11525
rect 11513 11520 18571 11522
rect 11513 11464 11518 11520
rect 11574 11464 18510 11520
rect 18566 11464 18571 11520
rect 11513 11462 18571 11464
rect 11513 11459 11579 11462
rect 18505 11459 18571 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 7465 11384 10426 11386
rect 7465 11328 7470 11384
rect 7526 11328 10426 11384
rect 7465 11326 10426 11328
rect 10593 11386 10659 11389
rect 16205 11386 16271 11389
rect 10593 11384 16271 11386
rect 10593 11328 10598 11384
rect 10654 11328 16210 11384
rect 16266 11328 16271 11384
rect 10593 11326 16271 11328
rect 7465 11323 7531 11326
rect 10593 11323 10659 11326
rect 16205 11323 16271 11326
rect 8201 11250 8267 11253
rect 15745 11250 15811 11253
rect 8201 11248 15811 11250
rect 8201 11192 8206 11248
rect 8262 11192 15750 11248
rect 15806 11192 15811 11248
rect 8201 11190 15811 11192
rect 8201 11187 8267 11190
rect 15745 11187 15811 11190
rect 7097 11114 7163 11117
rect 8150 11114 8156 11116
rect 7097 11112 8156 11114
rect 7097 11056 7102 11112
rect 7158 11056 8156 11112
rect 7097 11054 8156 11056
rect 7097 11051 7163 11054
rect 8150 11052 8156 11054
rect 8220 11052 8226 11116
rect 8661 11114 8727 11117
rect 9581 11114 9647 11117
rect 8661 11112 9647 11114
rect 8661 11056 8666 11112
rect 8722 11056 9586 11112
rect 9642 11056 9647 11112
rect 8661 11054 9647 11056
rect 8661 11051 8727 11054
rect 9581 11051 9647 11054
rect 12341 11114 12407 11117
rect 13445 11114 13511 11117
rect 12341 11112 13511 11114
rect 12341 11056 12346 11112
rect 12402 11056 13450 11112
rect 13506 11056 13511 11112
rect 12341 11054 13511 11056
rect 12341 11051 12407 11054
rect 13445 11051 13511 11054
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 7281 10978 7347 10981
rect 7557 10978 7623 10981
rect 7281 10976 7623 10978
rect 7281 10920 7286 10976
rect 7342 10920 7562 10976
rect 7618 10920 7623 10976
rect 7281 10918 7623 10920
rect 7281 10915 7347 10918
rect 7557 10915 7623 10918
rect 12157 10978 12223 10981
rect 16205 10978 16271 10981
rect 12157 10976 16271 10978
rect 12157 10920 12162 10976
rect 12218 10920 16210 10976
rect 16266 10920 16271 10976
rect 12157 10918 16271 10920
rect 12157 10915 12223 10918
rect 16205 10915 16271 10918
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4245 10842 4311 10845
rect 4613 10842 4679 10845
rect 10777 10842 10843 10845
rect 4245 10840 10843 10842
rect 4245 10784 4250 10840
rect 4306 10784 4618 10840
rect 4674 10784 10782 10840
rect 10838 10784 10843 10840
rect 4245 10782 10843 10784
rect 4245 10779 4311 10782
rect 4613 10779 4679 10782
rect 10777 10779 10843 10782
rect 5717 10706 5783 10709
rect 11421 10706 11487 10709
rect 5717 10704 11487 10706
rect 5717 10648 5722 10704
rect 5778 10648 11426 10704
rect 11482 10648 11487 10704
rect 5717 10646 11487 10648
rect 5717 10643 5783 10646
rect 11421 10643 11487 10646
rect 8569 10570 8635 10573
rect 20161 10570 20227 10573
rect 20345 10570 20411 10573
rect 8569 10568 20411 10570
rect 8569 10512 8574 10568
rect 8630 10512 20166 10568
rect 20222 10512 20350 10568
rect 20406 10512 20411 10568
rect 8569 10510 20411 10512
rect 8569 10507 8635 10510
rect 20161 10507 20227 10510
rect 20345 10507 20411 10510
rect 6085 10434 6151 10437
rect 19374 10434 19380 10436
rect 6085 10432 19380 10434
rect 6085 10376 6090 10432
rect 6146 10376 19380 10432
rect 6085 10374 19380 10376
rect 6085 10371 6151 10374
rect 19374 10372 19380 10374
rect 19444 10372 19450 10436
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 5349 10298 5415 10301
rect 23565 10298 23631 10301
rect 5349 10296 23631 10298
rect 5349 10240 5354 10296
rect 5410 10240 23570 10296
rect 23626 10240 23631 10296
rect 5349 10238 23631 10240
rect 5349 10235 5415 10238
rect 23565 10235 23631 10238
rect 7189 10162 7255 10165
rect 9581 10162 9647 10165
rect 7189 10160 9647 10162
rect 7189 10104 7194 10160
rect 7250 10104 9586 10160
rect 9642 10104 9647 10160
rect 7189 10102 9647 10104
rect 7189 10099 7255 10102
rect 9581 10099 9647 10102
rect 16481 10162 16547 10165
rect 18505 10162 18571 10165
rect 16481 10160 18571 10162
rect 16481 10104 16486 10160
rect 16542 10104 18510 10160
rect 18566 10104 18571 10160
rect 16481 10102 18571 10104
rect 16481 10099 16547 10102
rect 18505 10099 18571 10102
rect 10593 10026 10659 10029
rect 12709 10026 12775 10029
rect 13445 10026 13511 10029
rect 15653 10026 15719 10029
rect 10593 10024 12775 10026
rect 10593 9968 10598 10024
rect 10654 9968 12714 10024
rect 12770 9968 12775 10024
rect 10593 9966 12775 9968
rect 10593 9963 10659 9966
rect 12709 9963 12775 9966
rect 13080 10024 15719 10026
rect 13080 9968 13450 10024
rect 13506 9968 15658 10024
rect 15714 9968 15719 10024
rect 13080 9966 15719 9968
rect 10041 9890 10107 9893
rect 10542 9890 10548 9892
rect 10041 9888 10548 9890
rect 10041 9832 10046 9888
rect 10102 9832 10548 9888
rect 10041 9830 10548 9832
rect 10041 9827 10107 9830
rect 10542 9828 10548 9830
rect 10612 9890 10618 9892
rect 10961 9890 11027 9893
rect 10612 9888 11027 9890
rect 10612 9832 10966 9888
rect 11022 9832 11027 9888
rect 10612 9830 11027 9832
rect 10612 9828 10618 9830
rect 10961 9827 11027 9830
rect 12341 9890 12407 9893
rect 13080 9890 13140 9966
rect 13445 9963 13511 9966
rect 15653 9963 15719 9966
rect 12341 9888 13140 9890
rect 12341 9832 12346 9888
rect 12402 9832 13140 9888
rect 12341 9830 13140 9832
rect 14825 9890 14891 9893
rect 15469 9890 15535 9893
rect 14825 9888 15535 9890
rect 14825 9832 14830 9888
rect 14886 9832 15474 9888
rect 15530 9832 15535 9888
rect 14825 9830 15535 9832
rect 12341 9827 12407 9830
rect 14825 9827 14891 9830
rect 15469 9827 15535 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 13997 9618 14063 9621
rect 25221 9618 25287 9621
rect 13997 9616 25287 9618
rect 13997 9560 14002 9616
rect 14058 9560 25226 9616
rect 25282 9560 25287 9616
rect 13997 9558 25287 9560
rect 13997 9555 14063 9558
rect 25221 9555 25287 9558
rect 5993 9482 6059 9485
rect 20897 9482 20963 9485
rect 5993 9480 20963 9482
rect 5993 9424 5998 9480
rect 6054 9424 20902 9480
rect 20958 9424 20963 9480
rect 5993 9422 20963 9424
rect 5993 9419 6059 9422
rect 20897 9419 20963 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 11881 9210 11947 9213
rect 13169 9210 13235 9213
rect 11881 9208 13235 9210
rect 11881 9152 11886 9208
rect 11942 9152 13174 9208
rect 13230 9152 13235 9208
rect 11881 9150 13235 9152
rect 11881 9147 11947 9150
rect 13169 9147 13235 9150
rect 6545 9074 6611 9077
rect 8845 9074 8911 9077
rect 6545 9072 8911 9074
rect 6545 9016 6550 9072
rect 6606 9016 8850 9072
rect 8906 9016 8911 9072
rect 6545 9014 8911 9016
rect 6545 9011 6611 9014
rect 8845 9011 8911 9014
rect 10961 9074 11027 9077
rect 19057 9074 19123 9077
rect 10961 9072 19123 9074
rect 10961 9016 10966 9072
rect 11022 9016 19062 9072
rect 19118 9016 19123 9072
rect 10961 9014 19123 9016
rect 10961 9011 11027 9014
rect 19057 9011 19123 9014
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 3049 8664 3115 8669
rect 3049 8608 3054 8664
rect 3110 8608 3115 8664
rect 3049 8603 3115 8608
rect 2865 8394 2931 8397
rect 3052 8394 3112 8603
rect 8109 8530 8175 8533
rect 9397 8530 9463 8533
rect 8109 8528 9463 8530
rect 8109 8472 8114 8528
rect 8170 8472 9402 8528
rect 9458 8472 9463 8528
rect 8109 8470 9463 8472
rect 8109 8467 8175 8470
rect 9397 8467 9463 8470
rect 9622 8468 9628 8532
rect 9692 8530 9698 8532
rect 18413 8530 18479 8533
rect 19885 8530 19951 8533
rect 9692 8528 19951 8530
rect 9692 8472 18418 8528
rect 18474 8472 19890 8528
rect 19946 8472 19951 8528
rect 9692 8470 19951 8472
rect 9692 8468 9698 8470
rect 18413 8467 18479 8470
rect 19885 8467 19951 8470
rect 20161 8530 20227 8533
rect 20713 8530 20779 8533
rect 20161 8528 20779 8530
rect 20161 8472 20166 8528
rect 20222 8472 20718 8528
rect 20774 8472 20779 8528
rect 20161 8470 20779 8472
rect 20161 8467 20227 8470
rect 20713 8467 20779 8470
rect 2865 8392 3112 8394
rect 2865 8336 2870 8392
rect 2926 8336 3112 8392
rect 2865 8334 3112 8336
rect 4521 8394 4587 8397
rect 4981 8394 5047 8397
rect 5390 8394 5396 8396
rect 4521 8392 4768 8394
rect 4521 8336 4526 8392
rect 4582 8336 4768 8392
rect 4521 8334 4768 8336
rect 2865 8331 2931 8334
rect 4521 8331 4587 8334
rect 4708 8258 4768 8334
rect 4981 8392 5396 8394
rect 4981 8336 4986 8392
rect 5042 8336 5396 8392
rect 4981 8334 5396 8336
rect 4981 8331 5047 8334
rect 5390 8332 5396 8334
rect 5460 8332 5466 8396
rect 13813 8394 13879 8397
rect 14365 8394 14431 8397
rect 13813 8392 14431 8394
rect 13813 8336 13818 8392
rect 13874 8336 14370 8392
rect 14426 8336 14431 8392
rect 13813 8334 14431 8336
rect 13813 8331 13879 8334
rect 14365 8331 14431 8334
rect 15745 8394 15811 8397
rect 21265 8394 21331 8397
rect 15745 8392 21331 8394
rect 15745 8336 15750 8392
rect 15806 8336 21270 8392
rect 21326 8336 21331 8392
rect 15745 8334 21331 8336
rect 15745 8331 15811 8334
rect 21265 8331 21331 8334
rect 4981 8258 5047 8261
rect 4708 8256 5047 8258
rect 4708 8200 4986 8256
rect 5042 8200 5047 8256
rect 4708 8198 5047 8200
rect 4981 8195 5047 8198
rect 14457 8258 14523 8261
rect 18413 8258 18479 8261
rect 14457 8256 18479 8258
rect 14457 8200 14462 8256
rect 14518 8200 18418 8256
rect 18474 8200 18479 8256
rect 14457 8198 18479 8200
rect 14457 8195 14523 8198
rect 18413 8195 18479 8198
rect 20069 8258 20135 8261
rect 20253 8258 20319 8261
rect 20069 8256 20319 8258
rect 20069 8200 20074 8256
rect 20130 8200 20258 8256
rect 20314 8200 20319 8256
rect 20069 8198 20319 8200
rect 20069 8195 20135 8198
rect 20253 8195 20319 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19333 7986 19399 7989
rect 19290 7984 19399 7986
rect 19290 7928 19338 7984
rect 19394 7928 19399 7984
rect 19290 7923 19399 7928
rect 11278 7788 11284 7852
rect 11348 7850 11354 7852
rect 12157 7850 12223 7853
rect 11348 7848 12223 7850
rect 11348 7792 12162 7848
rect 12218 7792 12223 7848
rect 11348 7790 12223 7792
rect 11348 7788 11354 7790
rect 12157 7787 12223 7790
rect 200 7578 800 7608
rect 1393 7578 1459 7581
rect 200 7576 1459 7578
rect 200 7520 1398 7576
rect 1454 7520 1459 7576
rect 200 7518 1459 7520
rect 200 7488 800 7518
rect 1393 7515 1459 7518
rect 13997 7578 14063 7581
rect 15745 7578 15811 7581
rect 17769 7578 17835 7581
rect 13997 7576 17835 7578
rect 13997 7520 14002 7576
rect 14058 7520 15750 7576
rect 15806 7520 17774 7576
rect 17830 7520 17835 7576
rect 13997 7518 17835 7520
rect 13997 7515 14063 7518
rect 15745 7515 15811 7518
rect 17769 7515 17835 7518
rect 13997 7442 14063 7445
rect 15377 7442 15443 7445
rect 13997 7440 15443 7442
rect 13997 7384 14002 7440
rect 14058 7384 15382 7440
rect 15438 7384 15443 7440
rect 13997 7382 15443 7384
rect 13997 7379 14063 7382
rect 15377 7379 15443 7382
rect 9949 7170 10015 7173
rect 17493 7170 17559 7173
rect 9949 7168 17559 7170
rect 9949 7112 9954 7168
rect 10010 7112 17498 7168
rect 17554 7112 17559 7168
rect 9949 7110 17559 7112
rect 19290 7170 19350 7923
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 19425 7442 19491 7445
rect 22921 7442 22987 7445
rect 19425 7440 22987 7442
rect 19425 7384 19430 7440
rect 19486 7384 22926 7440
rect 22982 7384 22987 7440
rect 19425 7382 22987 7384
rect 19425 7379 19491 7382
rect 22921 7379 22987 7382
rect 19425 7306 19491 7309
rect 20161 7306 20227 7309
rect 19425 7304 20227 7306
rect 19425 7248 19430 7304
rect 19486 7248 20166 7304
rect 20222 7248 20227 7304
rect 19425 7246 20227 7248
rect 19425 7243 19491 7246
rect 20161 7243 20227 7246
rect 19425 7170 19491 7173
rect 19290 7168 19491 7170
rect 19290 7112 19430 7168
rect 19486 7112 19491 7168
rect 19290 7110 19491 7112
rect 9949 7107 10015 7110
rect 17493 7107 17559 7110
rect 19425 7107 19491 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 8150 6972 8156 7036
rect 8220 7034 8226 7036
rect 12341 7034 12407 7037
rect 8220 7032 12407 7034
rect 8220 6976 12346 7032
rect 12402 6976 12407 7032
rect 8220 6974 12407 6976
rect 8220 6972 8226 6974
rect 12341 6971 12407 6974
rect 15837 7034 15903 7037
rect 17401 7034 17467 7037
rect 15837 7032 17467 7034
rect 15837 6976 15842 7032
rect 15898 6976 17406 7032
rect 17462 6976 17467 7032
rect 15837 6974 17467 6976
rect 15837 6971 15903 6974
rect 17401 6971 17467 6974
rect 10685 6900 10751 6901
rect 10685 6896 10732 6900
rect 10796 6898 10802 6900
rect 12249 6898 12315 6901
rect 12433 6898 12499 6901
rect 10685 6840 10690 6896
rect 10685 6836 10732 6840
rect 10796 6838 10842 6898
rect 12249 6896 12499 6898
rect 12249 6840 12254 6896
rect 12310 6840 12438 6896
rect 12494 6840 12499 6896
rect 12249 6838 12499 6840
rect 10796 6836 10802 6838
rect 10685 6835 10751 6836
rect 12249 6835 12315 6838
rect 12433 6835 12499 6838
rect 19885 6898 19951 6901
rect 21357 6898 21423 6901
rect 19885 6896 21423 6898
rect 19885 6840 19890 6896
rect 19946 6840 21362 6896
rect 21418 6840 21423 6896
rect 19885 6838 21423 6840
rect 19885 6835 19951 6838
rect 21357 6835 21423 6838
rect 2957 6762 3023 6765
rect 6269 6762 6335 6765
rect 10133 6762 10199 6765
rect 2957 6760 10199 6762
rect 2957 6704 2962 6760
rect 3018 6704 6274 6760
rect 6330 6704 10138 6760
rect 10194 6704 10199 6760
rect 2957 6702 10199 6704
rect 2957 6699 3023 6702
rect 6269 6699 6335 6702
rect 10133 6699 10199 6702
rect 11697 6762 11763 6765
rect 13077 6762 13143 6765
rect 11697 6760 13143 6762
rect 11697 6704 11702 6760
rect 11758 6704 13082 6760
rect 13138 6704 13143 6760
rect 11697 6702 13143 6704
rect 11697 6699 11763 6702
rect 13077 6699 13143 6702
rect 16573 6762 16639 6765
rect 18137 6762 18203 6765
rect 16573 6760 18203 6762
rect 16573 6704 16578 6760
rect 16634 6704 18142 6760
rect 18198 6704 18203 6760
rect 16573 6702 18203 6704
rect 16573 6699 16639 6702
rect 18137 6699 18203 6702
rect 20161 6762 20227 6765
rect 23289 6762 23355 6765
rect 20161 6760 23355 6762
rect 20161 6704 20166 6760
rect 20222 6704 23294 6760
rect 23350 6704 23355 6760
rect 20161 6702 23355 6704
rect 20161 6699 20227 6702
rect 23289 6699 23355 6702
rect 12249 6626 12315 6629
rect 12433 6626 12499 6629
rect 12249 6624 12499 6626
rect 12249 6568 12254 6624
rect 12310 6568 12438 6624
rect 12494 6568 12499 6624
rect 12249 6566 12499 6568
rect 12249 6563 12315 6566
rect 12433 6563 12499 6566
rect 20253 6626 20319 6629
rect 20897 6626 20963 6629
rect 20253 6624 20963 6626
rect 20253 6568 20258 6624
rect 20314 6568 20902 6624
rect 20958 6568 20963 6624
rect 20253 6566 20963 6568
rect 20253 6563 20319 6566
rect 20897 6563 20963 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 6637 6492 6703 6493
rect 6637 6490 6684 6492
rect 6592 6488 6684 6490
rect 6592 6432 6642 6488
rect 6592 6430 6684 6432
rect 6637 6428 6684 6430
rect 6748 6428 6754 6492
rect 13997 6490 14063 6493
rect 16665 6490 16731 6493
rect 9630 6488 14063 6490
rect 9630 6432 14002 6488
rect 14058 6432 14063 6488
rect 9630 6430 14063 6432
rect 6637 6427 6703 6428
rect 3785 6354 3851 6357
rect 5901 6354 5967 6357
rect 9630 6354 9690 6430
rect 13997 6427 14063 6430
rect 14598 6488 16731 6490
rect 14598 6432 16670 6488
rect 16726 6432 16731 6488
rect 14598 6430 16731 6432
rect 3785 6352 9690 6354
rect 3785 6296 3790 6352
rect 3846 6296 5906 6352
rect 5962 6296 9690 6352
rect 3785 6294 9690 6296
rect 3785 6291 3851 6294
rect 5901 6291 5967 6294
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 6361 6218 6427 6221
rect 6913 6218 6979 6221
rect 6361 6216 6979 6218
rect 6361 6160 6366 6216
rect 6422 6160 6918 6216
rect 6974 6160 6979 6216
rect 6361 6158 6979 6160
rect 6361 6155 6427 6158
rect 6913 6155 6979 6158
rect 10409 6218 10475 6221
rect 11053 6218 11119 6221
rect 10409 6216 11119 6218
rect 10409 6160 10414 6216
rect 10470 6160 11058 6216
rect 11114 6160 11119 6216
rect 10409 6158 11119 6160
rect 10409 6155 10475 6158
rect 11053 6155 11119 6158
rect 9949 6082 10015 6085
rect 14598 6082 14658 6430
rect 16665 6427 16731 6430
rect 14825 6354 14891 6357
rect 37733 6354 37799 6357
rect 14825 6352 37799 6354
rect 14825 6296 14830 6352
rect 14886 6296 37738 6352
rect 37794 6296 37799 6352
rect 14825 6294 37799 6296
rect 14825 6291 14891 6294
rect 37733 6291 37799 6294
rect 37457 6218 37523 6221
rect 39200 6218 39800 6248
rect 37457 6216 39800 6218
rect 37457 6160 37462 6216
rect 37518 6160 39800 6216
rect 37457 6158 39800 6160
rect 37457 6155 37523 6158
rect 39200 6128 39800 6158
rect 9949 6080 14658 6082
rect 9949 6024 9954 6080
rect 10010 6024 14658 6080
rect 9949 6022 14658 6024
rect 9949 6019 10015 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 8201 5946 8267 5949
rect 12617 5946 12683 5949
rect 8201 5944 12683 5946
rect 8201 5888 8206 5944
rect 8262 5888 12622 5944
rect 12678 5888 12683 5944
rect 8201 5886 12683 5888
rect 8201 5883 8267 5886
rect 12617 5883 12683 5886
rect 17953 5946 18019 5949
rect 21081 5946 21147 5949
rect 17953 5944 21147 5946
rect 17953 5888 17958 5944
rect 18014 5888 21086 5944
rect 21142 5888 21147 5944
rect 17953 5886 21147 5888
rect 17953 5883 18019 5886
rect 21081 5883 21147 5886
rect 6545 5810 6611 5813
rect 7189 5810 7255 5813
rect 6545 5808 7255 5810
rect 6545 5752 6550 5808
rect 6606 5752 7194 5808
rect 7250 5752 7255 5808
rect 6545 5750 7255 5752
rect 6545 5747 6611 5750
rect 7189 5747 7255 5750
rect 8293 5812 8359 5813
rect 8293 5808 8340 5812
rect 8404 5810 8410 5812
rect 8937 5810 9003 5813
rect 9397 5810 9463 5813
rect 10409 5810 10475 5813
rect 10869 5812 10935 5813
rect 10869 5810 10916 5812
rect 8293 5752 8298 5808
rect 8293 5748 8340 5752
rect 8404 5750 8450 5810
rect 8937 5808 10475 5810
rect 8937 5752 8942 5808
rect 8998 5752 9402 5808
rect 9458 5752 10414 5808
rect 10470 5752 10475 5808
rect 8937 5750 10475 5752
rect 10824 5808 10916 5810
rect 10824 5752 10874 5808
rect 10824 5750 10916 5752
rect 8404 5748 8410 5750
rect 8293 5747 8359 5748
rect 8937 5747 9003 5750
rect 9397 5747 9463 5750
rect 10409 5747 10475 5750
rect 10869 5748 10916 5750
rect 10980 5748 10986 5812
rect 11053 5810 11119 5813
rect 14549 5810 14615 5813
rect 11053 5808 14615 5810
rect 11053 5752 11058 5808
rect 11114 5752 14554 5808
rect 14610 5752 14615 5808
rect 11053 5750 14615 5752
rect 10869 5747 10935 5748
rect 11053 5747 11119 5750
rect 14549 5747 14615 5750
rect 8201 5674 8267 5677
rect 8201 5672 19442 5674
rect 8201 5616 8206 5672
rect 8262 5616 19442 5672
rect 8201 5614 19442 5616
rect 8201 5611 8267 5614
rect 6269 5538 6335 5541
rect 7833 5538 7899 5541
rect 6269 5536 7899 5538
rect 6269 5480 6274 5536
rect 6330 5480 7838 5536
rect 7894 5480 7899 5536
rect 6269 5478 7899 5480
rect 6269 5475 6335 5478
rect 7833 5475 7899 5478
rect 7189 5402 7255 5405
rect 9029 5404 9095 5405
rect 7598 5402 7604 5404
rect 7189 5400 7604 5402
rect 7189 5344 7194 5400
rect 7250 5344 7604 5400
rect 7189 5342 7604 5344
rect 7189 5339 7255 5342
rect 7598 5340 7604 5342
rect 7668 5340 7674 5404
rect 9029 5402 9076 5404
rect 8984 5400 9076 5402
rect 8984 5344 9034 5400
rect 8984 5342 9076 5344
rect 9029 5340 9076 5342
rect 9140 5340 9146 5404
rect 12157 5402 12223 5405
rect 15653 5402 15719 5405
rect 12157 5400 15719 5402
rect 12157 5344 12162 5400
rect 12218 5344 15658 5400
rect 15714 5344 15719 5400
rect 12157 5342 15719 5344
rect 9029 5339 9095 5340
rect 12157 5339 12223 5342
rect 15653 5339 15719 5342
rect 9489 5266 9555 5269
rect 9765 5266 9831 5269
rect 9489 5264 9831 5266
rect 9489 5208 9494 5264
rect 9550 5208 9770 5264
rect 9826 5208 9831 5264
rect 9489 5206 9831 5208
rect 9489 5203 9555 5206
rect 9765 5203 9831 5206
rect 10133 5266 10199 5269
rect 11973 5266 12039 5269
rect 10133 5264 12039 5266
rect 10133 5208 10138 5264
rect 10194 5208 11978 5264
rect 12034 5208 12039 5264
rect 10133 5206 12039 5208
rect 10133 5203 10199 5206
rect 11973 5203 12039 5206
rect 12433 5266 12499 5269
rect 12985 5266 13051 5269
rect 12433 5264 13051 5266
rect 12433 5208 12438 5264
rect 12494 5208 12990 5264
rect 13046 5208 13051 5264
rect 12433 5206 13051 5208
rect 19382 5266 19442 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 23289 5266 23355 5269
rect 19382 5264 23355 5266
rect 19382 5208 23294 5264
rect 23350 5208 23355 5264
rect 19382 5206 23355 5208
rect 12433 5203 12499 5206
rect 12985 5203 13051 5206
rect 23289 5203 23355 5206
rect 6821 5130 6887 5133
rect 10409 5130 10475 5133
rect 6821 5128 10475 5130
rect 6821 5072 6826 5128
rect 6882 5072 10414 5128
rect 10470 5072 10475 5128
rect 6821 5070 10475 5072
rect 6821 5067 6887 5070
rect 10409 5067 10475 5070
rect 11421 4994 11487 4997
rect 16062 4994 16068 4996
rect 11421 4992 16068 4994
rect 11421 4936 11426 4992
rect 11482 4936 16068 4992
rect 11421 4934 16068 4936
rect 11421 4931 11487 4934
rect 16062 4932 16068 4934
rect 16132 4932 16138 4996
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1301 4858 1367 4861
rect 200 4856 1367 4858
rect 200 4800 1306 4856
rect 1362 4800 1367 4856
rect 200 4798 1367 4800
rect 200 4768 800 4798
rect 1301 4795 1367 4798
rect 16021 4858 16087 4861
rect 16246 4858 16252 4860
rect 16021 4856 16252 4858
rect 16021 4800 16026 4856
rect 16082 4800 16252 4856
rect 16021 4798 16252 4800
rect 16021 4795 16087 4798
rect 16246 4796 16252 4798
rect 16316 4796 16322 4860
rect 3049 4722 3115 4725
rect 9857 4722 9923 4725
rect 3049 4720 9923 4722
rect 3049 4664 3054 4720
rect 3110 4664 9862 4720
rect 9918 4664 9923 4720
rect 3049 4662 9923 4664
rect 3049 4659 3115 4662
rect 9857 4659 9923 4662
rect 15193 4722 15259 4725
rect 23197 4722 23263 4725
rect 15193 4720 23263 4722
rect 15193 4664 15198 4720
rect 15254 4664 23202 4720
rect 23258 4664 23263 4720
rect 15193 4662 23263 4664
rect 15193 4659 15259 4662
rect 23197 4659 23263 4662
rect 5441 4586 5507 4589
rect 18965 4586 19031 4589
rect 5441 4584 19031 4586
rect 5441 4528 5446 4584
rect 5502 4528 18970 4584
rect 19026 4528 19031 4584
rect 5441 4526 19031 4528
rect 5441 4523 5507 4526
rect 18965 4523 19031 4526
rect 10869 4450 10935 4453
rect 19057 4450 19123 4453
rect 10869 4448 19123 4450
rect 10869 4392 10874 4448
rect 10930 4392 19062 4448
rect 19118 4392 19123 4448
rect 10869 4390 19123 4392
rect 10869 4387 10935 4390
rect 19057 4387 19123 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 7649 4314 7715 4317
rect 9581 4314 9647 4317
rect 7649 4312 9647 4314
rect 7649 4256 7654 4312
rect 7710 4256 9586 4312
rect 9642 4256 9647 4312
rect 7649 4254 9647 4256
rect 7649 4251 7715 4254
rect 9581 4251 9647 4254
rect 9765 4178 9831 4181
rect 12198 4178 12204 4180
rect 9765 4176 12204 4178
rect 9765 4120 9770 4176
rect 9826 4120 12204 4176
rect 9765 4118 12204 4120
rect 9765 4115 9831 4118
rect 12198 4116 12204 4118
rect 12268 4116 12274 4180
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 3918 3980 3924 4044
rect 3988 4042 3994 4044
rect 10317 4042 10383 4045
rect 3988 4040 10383 4042
rect 3988 3984 10322 4040
rect 10378 3984 10383 4040
rect 3988 3982 10383 3984
rect 3988 3980 3994 3982
rect 10317 3979 10383 3982
rect 14273 3906 14339 3909
rect 19333 3906 19399 3909
rect 14273 3904 19399 3906
rect 14273 3848 14278 3904
rect 14334 3848 19338 3904
rect 19394 3848 19399 3904
rect 14273 3846 19399 3848
rect 14273 3843 14339 3846
rect 19333 3843 19399 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 6126 3708 6132 3772
rect 6196 3770 6202 3772
rect 13537 3770 13603 3773
rect 6196 3768 13603 3770
rect 6196 3712 13542 3768
rect 13598 3712 13603 3768
rect 6196 3710 13603 3712
rect 6196 3708 6202 3710
rect 13537 3707 13603 3710
rect 15929 3770 15995 3773
rect 16062 3770 16068 3772
rect 15929 3768 16068 3770
rect 15929 3712 15934 3768
rect 15990 3712 16068 3768
rect 15929 3710 16068 3712
rect 15929 3707 15995 3710
rect 16062 3708 16068 3710
rect 16132 3708 16138 3772
rect 12893 3634 12959 3637
rect 19517 3634 19583 3637
rect 20069 3634 20135 3637
rect 20253 3634 20319 3637
rect 12893 3632 20319 3634
rect 12893 3576 12898 3632
rect 12954 3576 19522 3632
rect 19578 3576 20074 3632
rect 20130 3576 20258 3632
rect 20314 3576 20319 3632
rect 12893 3574 20319 3576
rect 12893 3571 12959 3574
rect 19517 3571 19583 3574
rect 20069 3571 20135 3574
rect 20253 3571 20319 3574
rect 4245 3498 4311 3501
rect 8334 3498 8340 3500
rect 4245 3496 8340 3498
rect 4245 3440 4250 3496
rect 4306 3440 8340 3496
rect 4245 3438 8340 3440
rect 4245 3435 4311 3438
rect 8334 3436 8340 3438
rect 8404 3436 8410 3500
rect 9765 3498 9831 3501
rect 16481 3498 16547 3501
rect 20621 3498 20687 3501
rect 9765 3496 16314 3498
rect 9765 3440 9770 3496
rect 9826 3440 16314 3496
rect 9765 3438 16314 3440
rect 9765 3435 9831 3438
rect 13813 3362 13879 3365
rect 15469 3362 15535 3365
rect 13813 3360 15535 3362
rect 13813 3304 13818 3360
rect 13874 3304 15474 3360
rect 15530 3304 15535 3360
rect 13813 3302 15535 3304
rect 16254 3362 16314 3438
rect 16481 3496 20687 3498
rect 16481 3440 16486 3496
rect 16542 3440 20626 3496
rect 20682 3440 20687 3496
rect 16481 3438 20687 3440
rect 16481 3435 16547 3438
rect 20621 3435 20687 3438
rect 18505 3362 18571 3365
rect 16254 3360 18571 3362
rect 16254 3304 18510 3360
rect 18566 3304 18571 3360
rect 16254 3302 18571 3304
rect 13813 3299 13879 3302
rect 15469 3299 15535 3302
rect 18505 3299 18571 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 10225 3226 10291 3229
rect 17125 3226 17191 3229
rect 10225 3224 17191 3226
rect 10225 3168 10230 3224
rect 10286 3168 17130 3224
rect 17186 3168 17191 3224
rect 10225 3166 17191 3168
rect 10225 3163 10291 3166
rect 17125 3163 17191 3166
rect 14457 3090 14523 3093
rect 25773 3090 25839 3093
rect 14457 3088 25839 3090
rect 14457 3032 14462 3088
rect 14518 3032 25778 3088
rect 25834 3032 25839 3088
rect 14457 3030 25839 3032
rect 14457 3027 14523 3030
rect 25773 3027 25839 3030
rect 13629 2954 13695 2957
rect 15193 2954 15259 2957
rect 19425 2956 19491 2957
rect 13629 2952 15259 2954
rect 13629 2896 13634 2952
rect 13690 2896 15198 2952
rect 15254 2896 15259 2952
rect 13629 2894 15259 2896
rect 13629 2891 13695 2894
rect 15193 2891 15259 2894
rect 19374 2892 19380 2956
rect 19444 2954 19491 2956
rect 19444 2952 19536 2954
rect 19486 2896 19536 2952
rect 19444 2894 19536 2896
rect 19444 2892 19491 2894
rect 19425 2891 19491 2892
rect 200 2818 800 2848
rect 1393 2818 1459 2821
rect 200 2816 1459 2818
rect 200 2760 1398 2816
rect 1454 2760 1459 2816
rect 200 2758 1459 2760
rect 200 2728 800 2758
rect 1393 2755 1459 2758
rect 12065 2818 12131 2821
rect 12433 2818 12499 2821
rect 12065 2816 12499 2818
rect 12065 2760 12070 2816
rect 12126 2760 12438 2816
rect 12494 2760 12499 2816
rect 12065 2758 12499 2760
rect 12065 2755 12131 2758
rect 12433 2755 12499 2758
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 16021 2682 16087 2685
rect 17166 2682 17172 2684
rect 16021 2680 17172 2682
rect 16021 2624 16026 2680
rect 16082 2624 17172 2680
rect 16021 2622 17172 2624
rect 16021 2619 16087 2622
rect 17166 2620 17172 2622
rect 17236 2620 17242 2684
rect 3182 2484 3188 2548
rect 3252 2546 3258 2548
rect 4705 2546 4771 2549
rect 3252 2544 4771 2546
rect 3252 2488 4710 2544
rect 4766 2488 4771 2544
rect 3252 2486 4771 2488
rect 3252 2484 3258 2486
rect 4705 2483 4771 2486
rect 16113 2546 16179 2549
rect 18873 2546 18939 2549
rect 16113 2544 18939 2546
rect 16113 2488 16118 2544
rect 16174 2488 18878 2544
rect 18934 2488 18939 2544
rect 16113 2486 18939 2488
rect 16113 2483 16179 2486
rect 18873 2483 18939 2486
rect 5390 2348 5396 2412
rect 5460 2410 5466 2412
rect 23473 2410 23539 2413
rect 5460 2408 23539 2410
rect 5460 2352 23478 2408
rect 23534 2352 23539 2408
rect 5460 2350 23539 2352
rect 5460 2348 5466 2350
rect 23473 2347 23539 2350
rect 13445 2274 13511 2277
rect 17953 2274 18019 2277
rect 13445 2272 18019 2274
rect 13445 2216 13450 2272
rect 13506 2216 17958 2272
rect 18014 2216 18019 2272
rect 13445 2214 18019 2216
rect 13445 2211 13511 2214
rect 17953 2211 18019 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1368 800 1398
rect 2773 1395 2839 1398
rect 37181 1458 37247 1461
rect 39200 1458 39800 1488
rect 37181 1456 39800 1458
rect 37181 1400 37186 1456
rect 37242 1400 39800 1456
rect 37181 1398 39800 1400
rect 37181 1395 37247 1398
rect 39200 1368 39800 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 9076 22612 9140 22676
rect 11284 22476 11348 22540
rect 16068 22340 16132 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 17172 21932 17236 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 10916 20708 10980 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 10732 19620 10796 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 12204 18728 12268 18732
rect 12204 18672 12254 18728
rect 12254 18672 12268 18728
rect 12204 18668 12268 18672
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 7604 18124 7668 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 6684 17852 6748 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 16252 16492 16316 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 9628 13908 9692 13972
rect 3188 13772 3252 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 3924 12548 3988 12612
rect 6132 12548 6196 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 10548 12412 10612 12476
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 8156 11052 8220 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 19380 10372 19444 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 10548 9828 10612 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 9628 8468 9692 8532
rect 5396 8332 5460 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 11284 7788 11348 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 8156 6972 8220 7036
rect 10732 6896 10796 6900
rect 10732 6840 10746 6896
rect 10746 6840 10796 6896
rect 10732 6836 10796 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 6684 6488 6748 6492
rect 6684 6432 6698 6488
rect 6698 6432 6748 6488
rect 6684 6428 6748 6432
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 8340 5808 8404 5812
rect 8340 5752 8354 5808
rect 8354 5752 8404 5808
rect 8340 5748 8404 5752
rect 10916 5808 10980 5812
rect 10916 5752 10930 5808
rect 10930 5752 10980 5808
rect 10916 5748 10980 5752
rect 7604 5340 7668 5404
rect 9076 5400 9140 5404
rect 9076 5344 9090 5400
rect 9090 5344 9140 5400
rect 9076 5340 9140 5344
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 16068 4932 16132 4996
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 16252 4796 16316 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 12204 4116 12268 4180
rect 3924 3980 3988 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 6132 3708 6196 3772
rect 16068 3708 16132 3772
rect 8340 3436 8404 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 19380 2952 19444 2956
rect 19380 2896 19430 2952
rect 19430 2896 19444 2952
rect 19380 2892 19444 2896
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 17172 2620 17236 2684
rect 3188 2484 3252 2548
rect 5396 2348 5460 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 9075 22676 9141 22677
rect 9075 22612 9076 22676
rect 9140 22612 9141 22676
rect 9075 22611 9141 22612
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 7603 18188 7669 18189
rect 7603 18124 7604 18188
rect 7668 18124 7669 18188
rect 7603 18123 7669 18124
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 6683 17916 6749 17917
rect 6683 17852 6684 17916
rect 6748 17852 6749 17916
rect 6683 17851 6749 17852
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3187 13836 3253 13837
rect 3187 13772 3188 13836
rect 3252 13772 3253 13836
rect 3187 13771 3253 13772
rect 3190 2549 3250 13771
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3923 12612 3989 12613
rect 3923 12548 3924 12612
rect 3988 12548 3989 12612
rect 3923 12547 3989 12548
rect 3926 4045 3986 12547
rect 4208 12544 4528 13568
rect 6131 12612 6197 12613
rect 6131 12548 6132 12612
rect 6196 12548 6197 12612
rect 6131 12547 6197 12548
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3187 2548 3253 2549
rect 3187 2484 3188 2548
rect 3252 2484 3253 2548
rect 3187 2483 3253 2484
rect 4208 2128 4528 2688
rect 5398 2413 5458 8331
rect 6134 3773 6194 12547
rect 6686 6493 6746 17851
rect 6683 6492 6749 6493
rect 6683 6428 6684 6492
rect 6748 6428 6749 6492
rect 6683 6427 6749 6428
rect 7606 5405 7666 18123
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 8158 7037 8218 11051
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 8339 5812 8405 5813
rect 8339 5748 8340 5812
rect 8404 5748 8405 5812
rect 8339 5747 8405 5748
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 6131 3772 6197 3773
rect 6131 3708 6132 3772
rect 6196 3708 6197 3772
rect 6131 3707 6197 3708
rect 8342 3501 8402 5747
rect 9078 5405 9138 22611
rect 11283 22540 11349 22541
rect 11283 22476 11284 22540
rect 11348 22476 11349 22540
rect 11283 22475 11349 22476
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 10731 19684 10797 19685
rect 10731 19620 10732 19684
rect 10796 19620 10797 19684
rect 10731 19619 10797 19620
rect 9627 13972 9693 13973
rect 9627 13908 9628 13972
rect 9692 13908 9693 13972
rect 9627 13907 9693 13908
rect 9630 8533 9690 13907
rect 10547 12476 10613 12477
rect 10547 12412 10548 12476
rect 10612 12412 10613 12476
rect 10547 12411 10613 12412
rect 10550 9893 10610 12411
rect 10547 9892 10613 9893
rect 10547 9828 10548 9892
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 9627 8532 9693 8533
rect 9627 8468 9628 8532
rect 9692 8468 9693 8532
rect 9627 8467 9693 8468
rect 10734 6901 10794 19619
rect 10731 6900 10797 6901
rect 10731 6836 10732 6900
rect 10796 6836 10797 6900
rect 10731 6835 10797 6836
rect 10918 5813 10978 20707
rect 11286 7853 11346 22475
rect 16067 22404 16133 22405
rect 16067 22340 16068 22404
rect 16132 22340 16133 22404
rect 16067 22339 16133 22340
rect 12203 18732 12269 18733
rect 12203 18668 12204 18732
rect 12268 18668 12269 18732
rect 12203 18667 12269 18668
rect 11283 7852 11349 7853
rect 11283 7788 11284 7852
rect 11348 7788 11349 7852
rect 11283 7787 11349 7788
rect 10915 5812 10981 5813
rect 10915 5748 10916 5812
rect 10980 5748 10981 5812
rect 10915 5747 10981 5748
rect 9075 5404 9141 5405
rect 9075 5340 9076 5404
rect 9140 5340 9141 5404
rect 9075 5339 9141 5340
rect 12206 4181 12266 18667
rect 16070 4997 16130 22339
rect 17171 21996 17237 21997
rect 17171 21932 17172 21996
rect 17236 21932 17237 21996
rect 17171 21931 17237 21932
rect 16251 16556 16317 16557
rect 16251 16492 16252 16556
rect 16316 16492 16317 16556
rect 16251 16491 16317 16492
rect 16067 4996 16133 4997
rect 16067 4932 16068 4996
rect 16132 4932 16133 4996
rect 16067 4931 16133 4932
rect 12203 4180 12269 4181
rect 12203 4116 12204 4180
rect 12268 4116 12269 4180
rect 12203 4115 12269 4116
rect 16070 3773 16130 4931
rect 16254 4861 16314 16491
rect 16251 4860 16317 4861
rect 16251 4796 16252 4860
rect 16316 4796 16317 4860
rect 16251 4795 16317 4796
rect 16067 3772 16133 3773
rect 16067 3708 16068 3772
rect 16132 3708 16133 3772
rect 16067 3707 16133 3708
rect 8339 3500 8405 3501
rect 8339 3436 8340 3500
rect 8404 3436 8405 3500
rect 8339 3435 8405 3436
rect 17174 2685 17234 21931
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 10436 19445 10437
rect 19379 10372 19380 10436
rect 19444 10372 19445 10436
rect 19379 10371 19445 10372
rect 19382 2957 19442 10371
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 2956 19445 2957
rect 19379 2892 19380 2956
rect 19444 2892 19445 2956
rect 19379 2891 19445 2892
rect 17171 2684 17237 2685
rect 17171 2620 17172 2684
rect 17236 2620 17237 2684
rect 17171 2619 17237 2620
rect 5395 2412 5461 2413
rect 5395 2348 5396 2412
rect 5460 2348 5461 2412
rect 5395 2347 5461 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform -1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform -1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform -1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1667941163
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1667941163
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1667941163
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1667941163
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1667941163
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1667941163
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_286 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1667941163
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1667941163
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1667941163
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_98
timestamp 1667941163
transform 1 0 10120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_191
timestamp 1667941163
transform 1 0 18676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_208
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1667941163
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1667941163
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1667941163
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1667941163
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_124
timestamp 1667941163
transform 1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1667941163
transform 1 0 13248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1667941163
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_210
timestamp 1667941163
transform 1 0 20424 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_218
timestamp 1667941163
transform 1 0 21160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1667941163
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_229
timestamp 1667941163
transform 1 0 22172 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1667941163
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1667941163
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_383
timestamp 1667941163
transform 1 0 36340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_395
timestamp 1667941163
transform 1 0 37444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1667941163
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1667941163
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1667941163
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1667941163
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1667941163
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1667941163
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1667941163
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1667941163
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1667941163
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1667941163
transform 1 0 18032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1667941163
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1667941163
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1667941163
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_211
timestamp 1667941163
transform 1 0 20516 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1667941163
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_236
timestamp 1667941163
transform 1 0 22816 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1667941163
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1667941163
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1667941163
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_264
timestamp 1667941163
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1667941163
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_401
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1667941163
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1667941163
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_50
timestamp 1667941163
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1667941163
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1667941163
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1667941163
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1667941163
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_208
timestamp 1667941163
transform 1 0 20240 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_216
timestamp 1667941163
transform 1 0 20976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_224
timestamp 1667941163
transform 1 0 21712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1667941163
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1667941163
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_242
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1667941163
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_293
timestamp 1667941163
transform 1 0 28060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1667941163
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1667941163
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1667941163
transform 1 0 33212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1667941163
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_17
timestamp 1667941163
transform 1 0 2668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1667941163
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1667941163
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_63
timestamp 1667941163
transform 1 0 6900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1667941163
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_92
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1667941163
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1667941163
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_120
timestamp 1667941163
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1667941163
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_154
timestamp 1667941163
transform 1 0 15272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_162
timestamp 1667941163
transform 1 0 16008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1667941163
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1667941163
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_209
timestamp 1667941163
transform 1 0 20332 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1667941163
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1667941163
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1667941163
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1667941163
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1667941163
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1667941163
transform 1 0 25944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1667941163
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1667941163
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1667941163
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1667941163
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1667941163
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_110
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1667941163
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1667941163
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1667941163
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1667941163
transform 1 0 18308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1667941163
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_214
timestamp 1667941163
transform 1 0 20792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1667941163
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1667941163
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_242
timestamp 1667941163
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1667941163
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_317
timestamp 1667941163
transform 1 0 30268 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_322
timestamp 1667941163
transform 1 0 30728 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_334
timestamp 1667941163
transform 1 0 31832 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_346
timestamp 1667941163
transform 1 0 32936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1667941163
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_17
timestamp 1667941163
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1667941163
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1667941163
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1667941163
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_118
timestamp 1667941163
transform 1 0 11960 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1667941163
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_204
timestamp 1667941163
transform 1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1667941163
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_242
timestamp 1667941163
transform 1 0 23368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_266
timestamp 1667941163
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1667941163
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1667941163
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_123
timestamp 1667941163
transform 1 0 12420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1667941163
transform 1 0 12788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1667941163
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 1667941163
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1667941163
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1667941163
transform 1 0 20424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1667941163
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_228
timestamp 1667941163
transform 1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_235
timestamp 1667941163
transform 1 0 22724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_242
timestamp 1667941163
transform 1 0 23368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1667941163
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_295
timestamp 1667941163
transform 1 0 28244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1667941163
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_351
timestamp 1667941163
transform 1 0 33396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1667941163
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_383
timestamp 1667941163
transform 1 0 36340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1667941163
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_399
timestamp 1667941163
transform 1 0 37812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1667941163
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1667941163
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1667941163
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1667941163
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1667941163
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1667941163
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1667941163
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1667941163
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1667941163
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_187
timestamp 1667941163
transform 1 0 18308 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1667941163
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1667941163
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1667941163
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 1667941163
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1667941163
transform 1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_244
timestamp 1667941163
transform 1 0 23552 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1667941163
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1667941163
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp 1667941163
transform 1 0 28612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_303
timestamp 1667941163
transform 1 0 28980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_315
timestamp 1667941163
transform 1 0 30084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1667941163
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1667941163
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1667941163
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1667941163
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1667941163
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1667941163
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1667941163
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp 1667941163
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1667941163
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_208
timestamp 1667941163
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1667941163
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_227
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_234
timestamp 1667941163
transform 1 0 22632 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_238
timestamp 1667941163
transform 1 0 23000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1667941163
transform 1 0 23368 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1667941163
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_282
timestamp 1667941163
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1667941163
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1667941163
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1667941163
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1667941163
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1667941163
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1667941163
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_121
timestamp 1667941163
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1667941163
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1667941163
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_162
timestamp 1667941163
transform 1 0 16008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1667941163
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1667941163
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_204
timestamp 1667941163
transform 1 0 19872 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_208
timestamp 1667941163
transform 1 0 20240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1667941163
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1667941163
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1667941163
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_255
timestamp 1667941163
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_262
timestamp 1667941163
transform 1 0 25208 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1667941163
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_356
timestamp 1667941163
transform 1 0 33856 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_368
timestamp 1667941163
transform 1 0 34960 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_380
timestamp 1667941163
transform 1 0 36064 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1667941163
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1667941163
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1667941163
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_129
timestamp 1667941163
transform 1 0 12972 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1667941163
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_176
timestamp 1667941163
transform 1 0 17296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1667941163
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1667941163
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_216
timestamp 1667941163
transform 1 0 20976 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_228
timestamp 1667941163
transform 1 0 22080 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1667941163
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_23
timestamp 1667941163
transform 1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1667941163
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1667941163
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1667941163
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_204
timestamp 1667941163
transform 1 0 19872 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1667941163
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1667941163
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_234
timestamp 1667941163
transform 1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_240
timestamp 1667941163
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_268
timestamp 1667941163
transform 1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1667941163
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1667941163
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_289
timestamp 1667941163
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_301
timestamp 1667941163
transform 1 0 28796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_313
timestamp 1667941163
transform 1 0 29900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_325
timestamp 1667941163
transform 1 0 31004 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 1667941163
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1667941163
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1667941163
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1667941163
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1667941163
transform 1 0 16100 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_171
timestamp 1667941163
transform 1 0 16836 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1667941163
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1667941163
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1667941163
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_222
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1667941163
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1667941163
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_370
timestamp 1667941163
transform 1 0 35144 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_382
timestamp 1667941163
transform 1 0 36248 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_394
timestamp 1667941163
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1667941163
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1667941163
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1667941163
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1667941163
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1667941163
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1667941163
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_100
timestamp 1667941163
transform 1 0 10304 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1667941163
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1667941163
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1667941163
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1667941163
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_183
timestamp 1667941163
transform 1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1667941163
transform 1 0 19412 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1667941163
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_242
timestamp 1667941163
transform 1 0 23368 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_268
timestamp 1667941163
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_19
timestamp 1667941163
transform 1 0 2852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1667941163
transform 1 0 5796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1667941163
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1667941163
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_128
timestamp 1667941163
transform 1 0 12880 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1667941163
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1667941163
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_176
timestamp 1667941163
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1667941163
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1667941163
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_217
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1667941163
transform 1 0 21988 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1667941163
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1667941163
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_280
timestamp 1667941163
transform 1 0 26864 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_284
timestamp 1667941163
transform 1 0 27232 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_296
timestamp 1667941163
transform 1 0 28336 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_8
timestamp 1667941163
transform 1 0 1840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1667941163
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_75
timestamp 1667941163
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1667941163
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_119
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_132
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1667941163
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1667941163
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_177
timestamp 1667941163
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_195
timestamp 1667941163
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1667941163
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1667941163
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1667941163
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1667941163
transform 1 0 24840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_265
timestamp 1667941163
transform 1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1667941163
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1667941163
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1667941163
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_34
timestamp 1667941163
transform 1 0 4232 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_42
timestamp 1667941163
transform 1 0 4968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1667941163
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1667941163
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1667941163
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1667941163
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_95
timestamp 1667941163
transform 1 0 9844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1667941163
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1667941163
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1667941163
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_152
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_175
timestamp 1667941163
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1667941163
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1667941163
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_236
timestamp 1667941163
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1667941163
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_270
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_282
timestamp 1667941163
transform 1 0 27048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_294
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_392
timestamp 1667941163
transform 1 0 37168 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_398
timestamp 1667941163
transform 1 0 37720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1667941163
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_26
timestamp 1667941163
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_43
timestamp 1667941163
transform 1 0 5060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1667941163
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1667941163
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1667941163
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 1667941163
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_92
timestamp 1667941163
transform 1 0 9568 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1667941163
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1667941163
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1667941163
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1667941163
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1667941163
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1667941163
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1667941163
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1667941163
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1667941163
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_179
timestamp 1667941163
transform 1 0 17572 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1667941163
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_195
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_203
timestamp 1667941163
transform 1 0 19780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_210
timestamp 1667941163
transform 1 0 20424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_268
timestamp 1667941163
transform 1 0 25760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1667941163
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_345
timestamp 1667941163
transform 1 0 32844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_357
timestamp 1667941163
transform 1 0 33948 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_369
timestamp 1667941163
transform 1 0 35052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_381
timestamp 1667941163
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1667941163
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_8
timestamp 1667941163
transform 1 0 1840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_19
timestamp 1667941163
transform 1 0 2852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_36
timestamp 1667941163
transform 1 0 4416 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_48
timestamp 1667941163
transform 1 0 5520 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1667941163
transform 1 0 6624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1667941163
transform 1 0 6992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1667941163
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_75
timestamp 1667941163
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1667941163
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1667941163
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1667941163
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_115
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_124
timestamp 1667941163
transform 1 0 12512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1667941163
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1667941163
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1667941163
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_166
timestamp 1667941163
transform 1 0 16376 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1667941163
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1667941163
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_203
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_224
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1667941163
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1667941163
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1667941163
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1667941163
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1667941163
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_8
timestamp 1667941163
transform 1 0 1840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1667941163
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_30
timestamp 1667941163
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1667941163
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1667941163
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1667941163
transform 1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_124
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_132
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_150
timestamp 1667941163
transform 1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1667941163
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_187
timestamp 1667941163
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_191
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_209
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_235
timestamp 1667941163
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_242
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_248
timestamp 1667941163
transform 1 0 23920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1667941163
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1667941163
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_8
timestamp 1667941163
transform 1 0 1840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_12
timestamp 1667941163
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1667941163
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_37
timestamp 1667941163
transform 1 0 4508 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_43
timestamp 1667941163
transform 1 0 5060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_55
timestamp 1667941163
transform 1 0 6164 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_67
timestamp 1667941163
transform 1 0 7268 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1667941163
transform 1 0 7636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1667941163
transform 1 0 8004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1667941163
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_100
timestamp 1667941163
transform 1 0 10304 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1667941163
transform 1 0 10856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1667941163
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1667941163
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_204
timestamp 1667941163
transform 1 0 19872 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_208
timestamp 1667941163
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1667941163
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_219
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_228
timestamp 1667941163
transform 1 0 22080 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1667941163
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_263
timestamp 1667941163
transform 1 0 25300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1667941163
transform 1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_284
timestamp 1667941163
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_296
timestamp 1667941163
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_63
timestamp 1667941163
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_67
timestamp 1667941163
transform 1 0 7268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_74
timestamp 1667941163
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1667941163
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1667941163
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_130
timestamp 1667941163
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1667941163
transform 1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1667941163
transform 1 0 15364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_186
timestamp 1667941163
transform 1 0 18216 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1667941163
transform 1 0 18768 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1667941163
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_236
timestamp 1667941163
transform 1 0 22816 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1667941163
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1667941163
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1667941163
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_345
timestamp 1667941163
transform 1 0 32844 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_350
timestamp 1667941163
transform 1 0 33304 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_362
timestamp 1667941163
transform 1 0 34408 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_374
timestamp 1667941163
transform 1 0 35512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1667941163
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_70
timestamp 1667941163
transform 1 0 7544 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_78
timestamp 1667941163
transform 1 0 8280 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_95
timestamp 1667941163
transform 1 0 9844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_111
timestamp 1667941163
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1667941163
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1667941163
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_152
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_160
timestamp 1667941163
transform 1 0 15824 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_184
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1667941163
transform 1 0 18584 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1667941163
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1667941163
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_75
timestamp 1667941163
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1667941163
transform 1 0 8648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1667941163
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1667941163
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1667941163
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1667941163
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191
timestamp 1667941163
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1667941163
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1667941163
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_258
timestamp 1667941163
transform 1 0 24840 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1667941163
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_57
timestamp 1667941163
transform 1 0 6348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1667941163
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1667941163
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_95
timestamp 1667941163
transform 1 0 9844 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1667941163
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1667941163
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1667941163
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_134
timestamp 1667941163
transform 1 0 13432 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1667941163
transform 1 0 16652 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1667941163
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_223
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1667941163
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_237
timestamp 1667941163
transform 1 0 22908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1667941163
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_281
timestamp 1667941163
transform 1 0 26956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_285
timestamp 1667941163
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 1667941163
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1667941163
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1667941163
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1667941163
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1667941163
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1667941163
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_101
timestamp 1667941163
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1667941163
transform 1 0 13064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_142
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp 1667941163
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_175
timestamp 1667941163
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_191
timestamp 1667941163
transform 1 0 18676 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1667941163
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1667941163
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_247
timestamp 1667941163
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_259
timestamp 1667941163
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1667941163
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_47
timestamp 1667941163
transform 1 0 5428 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_59
timestamp 1667941163
transform 1 0 6532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1667941163
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_116
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_124
timestamp 1667941163
transform 1 0 12512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1667941163
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_151
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1667941163
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_179
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1667941163
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1667941163
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1667941163
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1667941163
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1667941163
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1667941163
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_83
timestamp 1667941163
transform 1 0 8740 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_90
timestamp 1667941163
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1667941163
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1667941163
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1667941163
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1667941163
transform 1 0 15180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1667941163
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_244
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_256
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1667941163
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_353
timestamp 1667941163
transform 1 0 33580 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_365
timestamp 1667941163
transform 1 0 34684 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_377
timestamp 1667941163
transform 1 0 35788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1667941163
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1667941163
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1667941163
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_104
timestamp 1667941163
transform 1 0 10672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1667941163
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 1667941163
transform 1 0 12512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1667941163
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1667941163
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1667941163
transform 1 0 16560 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_203
timestamp 1667941163
transform 1 0 19780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1667941163
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_240
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1667941163
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_8
timestamp 1667941163
transform 1 0 1840 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_20
timestamp 1667941163
transform 1 0 2944 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_32
timestamp 1667941163
transform 1 0 4048 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_44
timestamp 1667941163
transform 1 0 5152 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_50
timestamp 1667941163
transform 1 0 5704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1667941163
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1667941163
transform 1 0 7636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_78
timestamp 1667941163
transform 1 0 8280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1667941163
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_92
timestamp 1667941163
transform 1 0 9568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1667941163
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_123
timestamp 1667941163
transform 1 0 12420 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1667941163
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1667941163
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1667941163
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_206
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1667941163
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1667941163
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_242
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1667941163
transform 1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1667941163
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_101
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_127
timestamp 1667941163
transform 1 0 12788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1667941163
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1667941163
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1667941163
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1667941163
transform 1 0 18124 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1667941163
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1667941163
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_314
timestamp 1667941163
transform 1 0 29992 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_326
timestamp 1667941163
transform 1 0 31096 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_338
timestamp 1667941163
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_350
timestamp 1667941163
transform 1 0 33304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1667941163
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_66
timestamp 1667941163
transform 1 0 7176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1667941163
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_80
timestamp 1667941163
transform 1 0 8464 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_87
timestamp 1667941163
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1667941163
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_127
timestamp 1667941163
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1667941163
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1667941163
transform 1 0 14352 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_148
timestamp 1667941163
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1667941163
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_187
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 1667941163
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1667941163
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_244
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_256
timestamp 1667941163
transform 1 0 24656 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_268
timestamp 1667941163
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_61
timestamp 1667941163
transform 1 0 6716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_66
timestamp 1667941163
transform 1 0 7176 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_108
timestamp 1667941163
transform 1 0 11040 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp 1667941163
transform 1 0 11776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1667941163
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_152
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1667941163
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_182
timestamp 1667941163
transform 1 0 17848 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1667941163
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_212
timestamp 1667941163
transform 1 0 20608 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 1667941163
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_272
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_284
timestamp 1667941163
transform 1 0 27232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_296
timestamp 1667941163
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1667941163
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_90
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1667941163
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_126
timestamp 1667941163
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_133
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_146
timestamp 1667941163
transform 1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_154
timestamp 1667941163
transform 1 0 15272 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_159
timestamp 1667941163
transform 1 0 15732 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_180
timestamp 1667941163
transform 1 0 17664 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_188
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1667941163
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_242
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_254
timestamp 1667941163
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_90
timestamp 1667941163
transform 1 0 9384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_104
timestamp 1667941163
transform 1 0 10672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_111
timestamp 1667941163
transform 1 0 11316 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1667941163
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1667941163
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1667941163
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1667941163
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_228
timestamp 1667941163
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_285
timestamp 1667941163
transform 1 0 27324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1667941163
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1667941163
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_103
timestamp 1667941163
transform 1 0 10580 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1667941163
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_159
timestamp 1667941163
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_178
timestamp 1667941163
transform 1 0 17480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_191
timestamp 1667941163
transform 1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1667941163
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1667941163
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_242
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_254
timestamp 1667941163
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_266
timestamp 1667941163
transform 1 0 25576 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_345
timestamp 1667941163
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_128
timestamp 1667941163
transform 1 0 12880 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_134
timestamp 1667941163
transform 1 0 13432 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1667941163
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_149
timestamp 1667941163
transform 1 0 14812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_175
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1667941163
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1667941163
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_237
timestamp 1667941163
transform 1 0 22908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1667941163
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_34
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1667941163
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_132
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1667941163
transform 1 0 13892 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_143
timestamp 1667941163
transform 1 0 14260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_147
timestamp 1667941163
transform 1 0 14628 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1667941163
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1667941163
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_183
timestamp 1667941163
transform 1 0 17940 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_192
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_170
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_182
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_208
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_219
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1667941163
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_238
timestamp 1667941163
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_351
timestamp 1667941163
transform 1 0 33396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1667941163
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_155
timestamp 1667941163
transform 1 0 15364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_159
timestamp 1667941163
transform 1 0 15732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_174
timestamp 1667941163
transform 1 0 17112 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1667941163
transform 1 0 18400 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_200
timestamp 1667941163
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_208
timestamp 1667941163
transform 1 0 20240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_212
timestamp 1667941163
transform 1 0 20608 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1667941163
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1667941163
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_100
timestamp 1667941163
transform 1 0 10304 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_112
timestamp 1667941163
transform 1 0 11408 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_124
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1667941163
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_163
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_182
timestamp 1667941163
transform 1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1667941163
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_214
timestamp 1667941163
transform 1 0 20792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_226
timestamp 1667941163
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1667941163
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_329
timestamp 1667941163
transform 1 0 31372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_335
timestamp 1667941163
transform 1 0 31924 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_342
timestamp 1667941163
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1667941163
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_74
timestamp 1667941163
transform 1 0 7912 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_86
timestamp 1667941163
transform 1 0 9016 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_98
timestamp 1667941163
transform 1 0 10120 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1667941163
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_186
timestamp 1667941163
transform 1 0 18216 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_190
timestamp 1667941163
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1667941163
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_78
timestamp 1667941163
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_90
timestamp 1667941163
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_102
timestamp 1667941163
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_289
timestamp 1667941163
transform 1 0 27692 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_295
timestamp 1667941163
transform 1 0 28244 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_307
timestamp 1667941163
transform 1 0 29348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_319
timestamp 1667941163
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1667941163
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_226
timestamp 1667941163
transform 1 0 21896 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_238
timestamp 1667941163
transform 1 0 23000 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_352
timestamp 1667941163
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_85
timestamp 1667941163
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_97
timestamp 1667941163
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_118
timestamp 1667941163
transform 1 0 11960 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_130
timestamp 1667941163
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_134
timestamp 1667941163
transform 1 0 13432 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_138
timestamp 1667941163
transform 1 0 13800 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_150
timestamp 1667941163
transform 1 0 14904 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1667941163
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_301
timestamp 1667941163
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_159
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_173
timestamp 1667941163
transform 1 0 17020 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_185
timestamp 1667941163
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1667941163
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_44
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1667941163
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_118
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_130
timestamp 1667941163
transform 1 0 13064 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_142
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_154
timestamp 1667941163
transform 1 0 15272 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1667941163
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_248
timestamp 1667941163
transform 1 0 23920 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_260
timestamp 1667941163
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1667941163
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_75
timestamp 1667941163
transform 1 0 8004 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_79
timestamp 1667941163
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_91
timestamp 1667941163
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1667941163
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_321
timestamp 1667941163
transform 1 0 30636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_56
timestamp 1667941163
transform 1 0 6256 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_68
timestamp 1667941163
transform 1 0 7360 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1667941163
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1667941163
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_99
timestamp 1667941163
transform 1 0 10212 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_111
timestamp 1667941163
transform 1 0 11316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_123
timestamp 1667941163
transform 1 0 12420 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_241
timestamp 1667941163
transform 1 0 23276 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1667941163
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_262
timestamp 1667941163
transform 1 0 25208 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_268
timestamp 1667941163
transform 1 0 25760 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_272
timestamp 1667941163
transform 1 0 26128 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1667941163
transform 1 0 27232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_288
timestamp 1667941163
transform 1 0 27600 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_292
timestamp 1667941163
transform 1 0 27968 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1667941163
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_353
timestamp 1667941163
transform 1 0 33580 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_359
timestamp 1667941163
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_340
timestamp 1667941163
transform 1 0 32384 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_352
timestamp 1667941163
transform 1 0 33488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1667941163
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1667941163
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1667941163
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1667941163
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_65
timestamp 1667941163
transform 1 0 7084 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_71
timestamp 1667941163
transform 1 0 7636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_83
timestamp 1667941163
transform 1 0 8740 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_95
timestamp 1667941163
transform 1 0 9844 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_107
timestamp 1667941163
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_174
timestamp 1667941163
transform 1 0 17112 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_186
timestamp 1667941163
transform 1 0 18216 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_198
timestamp 1667941163
transform 1 0 19320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_204
timestamp 1667941163
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_208
timestamp 1667941163
transform 1 0 20240 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_212
timestamp 1667941163
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_401
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_93
timestamp 1667941163
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_174
timestamp 1667941163
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1667941163
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1667941163
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 1667941163
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1667941163
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_328
timestamp 1667941163
transform 1 0 31280 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_335
timestamp 1667941163
transform 1 0 31924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_347
timestamp 1667941163
transform 1 0 33028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1667941163
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1667941163
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1667941163
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_141
timestamp 1667941163
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_145
timestamp 1667941163
transform 1 0 14444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_202
timestamp 1667941163
transform 1 0 19688 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_214
timestamp 1667941163
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1667941163
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 1667941163
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_245
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_257
timestamp 1667941163
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_70
timestamp 1667941163
transform 1 0 7544 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_129
timestamp 1667941163
transform 1 0 12972 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_135
timestamp 1667941163
transform 1 0 13524 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_146
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_158
timestamp 1667941163
transform 1 0 15640 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_170
timestamp 1667941163
transform 1 0 16744 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_182
timestamp 1667941163
transform 1 0 17848 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1667941163
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_174
timestamp 1667941163
transform 1 0 17112 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_186
timestamp 1667941163
transform 1 0 18216 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_198
timestamp 1667941163
transform 1 0 19320 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_210
timestamp 1667941163
transform 1 0 20424 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_233
timestamp 1667941163
transform 1 0 22540 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_239
timestamp 1667941163
transform 1 0 23092 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_251
timestamp 1667941163
transform 1 0 24196 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_263
timestamp 1667941163
transform 1 0 25300 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1667941163
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_106
timestamp 1667941163
transform 1 0 10856 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_118
timestamp 1667941163
transform 1 0 11960 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_130
timestamp 1667941163
transform 1 0 13064 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_162
timestamp 1667941163
transform 1 0 16008 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_174
timestamp 1667941163
transform 1 0 17112 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 1667941163
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_8
timestamp 1667941163
transform 1 0 1840 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_20
timestamp 1667941163
transform 1 0 2944 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_32
timestamp 1667941163
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1667941163
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1667941163
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_398
timestamp 1667941163
transform 1 0 37720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_8
timestamp 1667941163
transform 1 0 1840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1667941163
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1667941163
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1667941163
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1667941163
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1667941163
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_386
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0416_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 10396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 20976 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 20332 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 21620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 20240 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 22724 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 10120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 7728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 7636 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 13524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 11316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 8648 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 8464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 7360 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 25208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 25208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 25668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 26312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 25760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 25484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 25208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform 1 0 21804 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 21804 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 13064 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 23276 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 14352 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 14996 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 23368 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 20976 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 22080 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 23736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 19504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 20424 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 14536 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 15364 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1667941163
transform 1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1667941163
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 17204 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 18124 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 17480 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1667941163
transform 1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1667941163
transform 1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 8372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0607_
timestamp 1667941163
transform 1 0 26404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 9108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 9752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 9752 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 8648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 11040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1667941163
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1667941163
transform 1 0 10396 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 14996 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 8280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1667941163
transform 1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 21804 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 6716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1667941163
transform 1 0 7544 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 7728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 11684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 23000 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1667941163
transform 1 0 22632 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 23092 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1667941163
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 7820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform 1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1667941163
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1667941163
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1667941163
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1667941163
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 23276 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1667941163
transform 1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0708_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 27416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 7636 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 10580 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 9936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 24932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 31648 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 9292 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 28336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 32108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 7360 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 5428 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 32292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 8096 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 6992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 5152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 27968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 19596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 31004 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 33212 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 33488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 16744 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 14168 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 23460 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 15456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 33028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 29256 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 33580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 26128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 27048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 7820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 16836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 31648 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 36432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 8648 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 36064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 16928 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 33304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 22540 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 23368 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 13524 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0818_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 4140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 2576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 4784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0829_
timestamp 1667941163
transform 1 0 20976 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 2852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0840_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0851_
timestamp 1667941163
transform 1 0 23184 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 21804 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 20516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0862_
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0873_
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11040 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0891_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0893_
timestamp 1667941163
transform 1 0 11592 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0894_
timestamp 1667941163
transform 1 0 6716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0895_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0898_
timestamp 1667941163
transform 1 0 6072 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0900_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 9108 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0907_
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0908_
timestamp 1667941163
transform 1 0 7912 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 8188 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0912_
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 8924 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 3496 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0916_
timestamp 1667941163
transform 1 0 7268 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 3772 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0918_
timestamp 1667941163
transform 1 0 13340 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0919_
timestamp 1667941163
transform 1 0 7268 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 10304 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 6900 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform 1 0 6532 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0924_
timestamp 1667941163
transform 1 0 12512 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0925_
timestamp 1667941163
transform 1 0 9108 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform 1 0 11500 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 7084 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0929_
timestamp 1667941163
transform 1 0 10948 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0931_
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0932_
timestamp 1667941163
transform 1 0 11960 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0933_
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 6716 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 6164 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 13800 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0942_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0943_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 2944 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1667941163
transform 1 0 2852 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 14352 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 2852 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 11776 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 9292 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0960_
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0961_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1667941163
transform 1 0 16560 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0964_
timestamp 1667941163
transform 1 0 13984 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1667941163
transform 1 0 11776 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform -1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 33856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 22816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 33580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 23092 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 13248 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 16836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 37812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 34132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 15732 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 33856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 4784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 32936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 7268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 30452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 19412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 9752 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 2208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform -1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 33488 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1043__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15548 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1043_
timestamp 1667941163
transform 1 0 17572 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 15272 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1045_
timestamp 1667941163
transform 1 0 15364 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 16560 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1049__101
timestamp 1667941163
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1050_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 16836 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 16928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1055__102
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1057_
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1061__103
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 13432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 12604 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 19504 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1067__104
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 19320 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1073__105
timestamp 1667941163
transform 1 0 21620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 16192 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 9844 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1079__106
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1081_
timestamp 1667941163
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 11040 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1084_
timestamp 1667941163
transform 1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1085__107
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 20608 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1091__108
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 13892 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1093_
timestamp 1667941163
transform 1 0 12788 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 9568 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 14260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 18676 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1097__109
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 16928 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 20700 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 14996 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1103__110
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 14352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform 1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 15088 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 11960 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1109__111
timestamp 1667941163
transform 1 0 12972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 12972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 11684 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 21804 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1114_
timestamp 1667941163
transform 1 0 10212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1115__112
timestamp 1667941163
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 12328 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1117_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 11684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1120_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1121__113
timestamp 1667941163
transform 1 0 18584 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 14444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1123_
timestamp 1667941163
transform 1 0 19136 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1127__114
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform 1 0 17112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1132_
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1133__115
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 19964 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1135_
timestamp 1667941163
transform 1 0 22356 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 23184 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1139__116
timestamp 1667941163
transform 1 0 22632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1140_
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 22540 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 21344 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1144_
timestamp 1667941163
transform 1 0 16468 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 18032 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1145__117
timestamp 1667941163
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1147_
timestamp 1667941163
transform 1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 16928 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 17020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 19504 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1151__118
timestamp 1667941163
transform 1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 19504 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1154_
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1156_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1157__119
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 23092 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1159_
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1163__120
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1164_
timestamp 1667941163
transform 1 0 24380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 16560 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1166_
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 23644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1169__121
timestamp 1667941163
transform 1 0 24564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1172_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1174__122
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 11776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1178__123
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 19044 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1182_
timestamp 1667941163
transform 1 0 23276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1182__124
timestamp 1667941163
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1184_
timestamp 1667941163
transform 1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1186__125
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 15272 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1190__126
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 20424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1194__127
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 17572 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 10580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 11868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1198__128
timestamp 1667941163
transform 1 0 10672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 9292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 10120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1202__129
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform -1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 17664 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1206__130
timestamp 1667941163
transform 1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 9936 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 16468 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 8832 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1210__131
timestamp 1667941163
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1210_
timestamp 1667941163
transform 1 0 16744 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1212_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1214__132
timestamp 1667941163
transform 1 0 25668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 22816 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1215_
timestamp 1667941163
transform 1 0 17848 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1218__133
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 19044 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 17572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1222__134
timestamp 1667941163
transform 1 0 21988 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1222_
timestamp 1667941163
transform 1 0 20148 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1223_
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1224_
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1225_
timestamp 1667941163
transform 1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1226__135
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 20700 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 20608 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 22172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 13156 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1230__136
timestamp 1667941163
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 13340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform 1 0 12880 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1234__137
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1234_
timestamp 1667941163
transform 1 0 20424 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1236_
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1237_
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1667941163
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1667941163
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1667941163
transform 1 0 6808 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1667941163
transform 1 0 11776 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1667941163
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 38088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 3864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 2208 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 1564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 1564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1667941163
transform 1 0 6532 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 25760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 13432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 3 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 4 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 5 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 6 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 7 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 8 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 9 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 10 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 11 nsew signal input
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 12 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 13 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 14 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 15 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 16 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 17 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 18 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 19 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 20 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 21 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 22 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 23 nsew signal tristate
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 24 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 26 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 27 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 28 nsew signal tristate
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 29 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 30 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 32 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 33 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 34 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 35 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 36 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 37 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 38 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 78 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 79 nsew signal input
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 80 nsew signal input
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 81 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 82 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 83 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 84 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 85 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 86 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 87 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 pReset
port 88 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 prog_clk
port 89 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 90 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 91 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 96 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 97 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 98 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 99 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 vssd1
port 101 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 3910 9486 3910 9486 0 _0000_
rlabel metal1 3319 4522 3319 4522 0 _0001_
rlabel metal2 9798 5848 9798 5848 0 _0002_
rlabel metal2 3726 10948 3726 10948 0 _0003_
rlabel metal1 4094 12682 4094 12682 0 _0004_
rlabel metal1 7951 5270 7951 5270 0 _0005_
rlabel metal1 2576 8806 2576 8806 0 _0006_
rlabel metal2 14122 5542 14122 5542 0 _0007_
rlabel metal1 11040 6154 11040 6154 0 _0008_
rlabel metal1 5428 4794 5428 4794 0 _0009_
rlabel metal1 3680 9350 3680 9350 0 _0010_
rlabel metal1 2530 7514 2530 7514 0 _0011_
rlabel metal1 7038 5338 7038 5338 0 _0012_
rlabel via1 13754 8245 13754 8245 0 _0013_
rlabel metal1 11178 4114 11178 4114 0 _0014_
rlabel metal2 4094 5746 4094 5746 0 _0015_
rlabel metal2 2070 6936 2070 6936 0 _0016_
rlabel metal1 11040 5338 11040 5338 0 _0017_
rlabel metal1 3910 2822 3910 2822 0 _0018_
rlabel via2 20286 6613 20286 6613 0 _0019_
rlabel metal1 20378 10710 20378 10710 0 _0020_
rlabel metal1 21344 6426 21344 6426 0 _0021_
rlabel metal1 20516 5338 20516 5338 0 _0022_
rlabel metal2 12466 6341 12466 6341 0 _0023_
rlabel metal3 19412 5440 19412 5440 0 _0024_
rlabel metal1 19419 5610 19419 5610 0 _0025_
rlabel metal1 21160 5882 21160 5882 0 _0026_
rlabel metal1 20700 5542 20700 5542 0 _0027_
rlabel metal1 21206 5542 21206 5542 0 _0028_
rlabel metal2 20286 5066 20286 5066 0 _0029_
rlabel metal2 20102 6341 20102 6341 0 _0030_
rlabel metal1 16153 3434 16153 3434 0 _0031_
rlabel metal1 19642 2822 19642 2822 0 _0032_
rlabel metal2 23506 2329 23506 2329 0 _0033_
rlabel metal1 17342 2040 17342 2040 0 _0034_
rlabel metal1 3365 3434 3365 3434 0 _0035_
rlabel metal1 9522 5066 9522 5066 0 _0036_
rlabel metal1 16107 8942 16107 8942 0 _0037_
rlabel metal2 10442 3672 10442 3672 0 _0038_
rlabel metal2 5382 11033 5382 11033 0 _0039_
rlabel via2 19458 2907 19458 2907 0 _0040_
rlabel metal1 11592 5882 11592 5882 0 _0041_
rlabel metal1 13294 9996 13294 9996 0 _0042_
rlabel metal2 20378 4828 20378 4828 0 _0043_
rlabel metal2 12834 7990 12834 7990 0 _0044_
rlabel via1 22034 5525 22034 5525 0 _0045_
rlabel metal1 13715 2346 13715 2346 0 _0046_
rlabel metal1 10863 4522 10863 4522 0 _0047_
rlabel metal1 18170 3706 18170 3706 0 _0048_
rlabel metal2 20470 3298 20470 3298 0 _0049_
rlabel metal2 15594 2006 15594 2006 0 _0050_
rlabel metal1 21298 3910 21298 3910 0 _0051_
rlabel metal2 17986 4012 17986 4012 0 _0052_
rlabel metal2 22586 4318 22586 4318 0 _0053_
rlabel metal1 14674 4216 14674 4216 0 _0054_
rlabel metal1 9844 6630 9844 6630 0 _0055_
rlabel metal1 19366 9656 19366 9656 0 _0056_
rlabel metal1 8924 4794 8924 4794 0 _0057_
rlabel metal2 8510 12121 8510 12121 0 _0058_
rlabel metal1 8287 2346 8287 2346 0 _0059_
rlabel metal1 6118 12274 6118 12274 0 _0060_
rlabel metal1 4876 2278 4876 2278 0 _0061_
rlabel metal1 6854 8806 6854 8806 0 _0062_
rlabel metal1 5842 6222 5842 6222 0 _0063_
rlabel metal3 3979 2516 3979 2516 0 _0064_
rlabel metal1 5474 13158 5474 13158 0 _0065_
rlabel metal1 6900 6086 6900 6086 0 _0066_
rlabel metal2 2346 9724 2346 9724 0 _0067_
rlabel metal1 2530 14246 2530 14246 0 _0068_
rlabel metal2 4094 9112 4094 9112 0 _0069_
rlabel metal1 4830 12138 4830 12138 0 _0070_
rlabel metal1 3864 13362 3864 13362 0 _0071_
rlabel metal1 4692 13838 4692 13838 0 _0072_
rlabel metal1 6302 12750 6302 12750 0 _0073_
rlabel metal1 4232 13226 4232 13226 0 _0074_
rlabel metal1 5106 7514 5106 7514 0 _0075_
rlabel metal1 14858 13260 14858 13260 0 _0076_
rlabel metal1 21758 18258 21758 18258 0 _0077_
rlabel metal1 12926 13396 12926 13396 0 _0078_
rlabel metal1 8142 19686 8142 19686 0 _0079_
rlabel metal1 20976 21862 20976 21862 0 _0080_
rlabel metal1 21850 24208 21850 24208 0 _0081_
rlabel metal1 7728 11866 7728 11866 0 _0082_
rlabel metal2 22862 14756 22862 14756 0 _0083_
rlabel metal1 23920 4250 23920 4250 0 _0084_
rlabel metal2 20102 9350 20102 9350 0 _0085_
rlabel metal1 15594 22406 15594 22406 0 _0086_
rlabel metal1 23230 10030 23230 10030 0 _0087_
rlabel metal1 8602 13260 8602 13260 0 _0088_
rlabel metal2 9338 11526 9338 11526 0 _0089_
rlabel metal1 13340 11118 13340 11118 0 _0090_
rlabel metal3 8418 10132 8418 10132 0 _0091_
rlabel metal1 13248 6970 13248 6970 0 _0092_
rlabel metal1 18906 8976 18906 8976 0 _0093_
rlabel via2 19458 7259 19458 7259 0 _0094_
rlabel metal1 6946 18394 6946 18394 0 _0095_
rlabel metal2 9154 21692 9154 21692 0 _0096_
rlabel metal2 9246 14382 9246 14382 0 _0097_
rlabel metal1 14260 5882 14260 5882 0 _0098_
rlabel metal1 20562 21454 20562 21454 0 _0099_
rlabel metal1 12627 23086 12627 23086 0 _0100_
rlabel metal2 11546 20026 11546 20026 0 _0101_
rlabel viali 9246 11732 9246 11732 0 _0102_
rlabel metal1 20148 3978 20148 3978 0 _0103_
rlabel metal1 23920 7990 23920 7990 0 _0104_
rlabel metal1 8556 17850 8556 17850 0 _0105_
rlabel metal1 20194 13498 20194 13498 0 _0106_
rlabel metal1 8372 15674 8372 15674 0 _0107_
rlabel metal1 18308 3978 18308 3978 0 _0108_
rlabel metal1 25668 11730 25668 11730 0 _0109_
rlabel metal1 26542 14348 26542 14348 0 _0110_
rlabel metal1 25622 15130 25622 15130 0 _0111_
rlabel metal1 24518 8500 24518 8500 0 _0112_
rlabel via1 21942 6613 21942 6613 0 _0113_
rlabel metal2 22034 12920 22034 12920 0 _0114_
rlabel metal2 21298 14212 21298 14212 0 _0115_
rlabel metal1 23046 9146 23046 9146 0 _0116_
rlabel metal1 24380 15674 24380 15674 0 _0117_
rlabel metal1 20562 21114 20562 21114 0 _0118_
rlabel metal1 13754 21658 13754 21658 0 _0119_
rlabel metal1 18906 19414 18906 19414 0 _0120_
rlabel metal1 17434 24650 17434 24650 0 _0121_
rlabel metal1 15226 23732 15226 23732 0 _0122_
rlabel metal1 15594 21862 15594 21862 0 _0123_
rlabel metal2 20378 11084 20378 11084 0 _0124_
rlabel metal1 23690 12614 23690 12614 0 _0125_
rlabel metal2 23506 17034 23506 17034 0 _0126_
rlabel metal1 20792 14382 20792 14382 0 _0127_
rlabel metal1 23046 9894 23046 9894 0 _0128_
rlabel metal2 20194 13124 20194 13124 0 _0129_
rlabel metal1 15870 24378 15870 24378 0 _0130_
rlabel metal1 12535 21522 12535 21522 0 _0131_
rlabel metal1 16330 17646 16330 17646 0 _0132_
rlabel metal1 9982 18292 9982 18292 0 _0133_
rlabel metal1 17802 22746 17802 22746 0 _0134_
rlabel metal1 15916 23290 15916 23290 0 _0135_
rlabel metal2 6946 17340 6946 17340 0 _0136_
rlabel metal1 7544 13498 7544 13498 0 _0137_
rlabel metal2 11454 14858 11454 14858 0 _0138_
rlabel metal2 26634 13668 26634 13668 0 _0139_
rlabel metal1 9982 21488 9982 21488 0 _0140_
rlabel metal2 8418 20230 8418 20230 0 _0141_
rlabel metal1 14122 13906 14122 13906 0 _0142_
rlabel metal1 9062 17850 9062 17850 0 _0143_
rlabel metal2 13110 22406 13110 22406 0 _0144_
rlabel metal1 13478 14586 13478 14586 0 _0145_
rlabel metal1 14858 18938 14858 18938 0 _0146_
rlabel metal1 21850 20808 21850 20808 0 _0147_
rlabel metal1 13202 12070 13202 12070 0 _0148_
rlabel metal1 10534 13872 10534 13872 0 _0149_
rlabel metal2 9706 14518 9706 14518 0 _0150_
rlabel metal2 18170 12036 18170 12036 0 _0151_
rlabel metal1 18906 5712 18906 5712 0 _0152_
rlabel metal2 21022 10948 21022 10948 0 _0153_
rlabel metal1 7590 19380 7590 19380 0 _0154_
rlabel metal1 7544 16218 7544 16218 0 _0155_
rlabel metal1 7774 20570 7774 20570 0 _0156_
rlabel via2 9890 19363 9890 19363 0 _0157_
rlabel metal2 18446 14212 18446 14212 0 _0158_
rlabel metal1 23276 19346 23276 19346 0 _0159_
rlabel metal1 20700 17306 20700 17306 0 _0160_
rlabel metal2 17158 13294 17158 13294 0 _0161_
rlabel metal1 20516 14042 20516 14042 0 _0162_
rlabel metal1 15042 14246 15042 14246 0 _0163_
rlabel metal2 8418 17510 8418 17510 0 _0164_
rlabel metal1 9154 16218 9154 16218 0 _0165_
rlabel metal2 18906 15300 18906 15300 0 _0166_
rlabel metal1 16928 17306 16928 17306 0 _0167_
rlabel metal2 15870 19210 15870 19210 0 _0168_
rlabel metal1 24012 6766 24012 6766 0 _0169_
rlabel metal1 13524 5542 13524 5542 0 _0170_
rlabel metal2 17158 12036 17158 12036 0 _0171_
rlabel metal2 13846 13668 13846 13668 0 _0172_
rlabel metal2 17434 14586 17434 14586 0 _0173_
rlabel metal2 22034 3094 22034 3094 0 _0174_
rlabel metal2 21574 5100 21574 5100 0 _0175_
rlabel metal2 14030 6613 14030 6613 0 _0176_
rlabel metal2 14122 3774 14122 3774 0 _0177_
rlabel metal1 1978 8976 1978 8976 0 _0178_
rlabel metal2 23230 3876 23230 3876 0 _0179_
rlabel metal1 19458 4590 19458 4590 0 _0180_
rlabel metal1 20240 2414 20240 2414 0 _0181_
rlabel metal1 10396 11594 10396 11594 0 _0182_
rlabel metal1 17526 14586 17526 14586 0 _0183_
rlabel metal1 14536 12682 14536 12682 0 _0184_
rlabel metal1 8418 10438 8418 10438 0 _0185_
rlabel metal1 14306 12954 14306 12954 0 _0186_
rlabel metal1 20194 17816 20194 17816 0 _0187_
rlabel metal1 17434 12410 17434 12410 0 _0188_
rlabel metal1 15594 8024 15594 8024 0 _0189_
rlabel via2 20194 6715 20194 6715 0 _0190_
rlabel metal1 16652 5338 16652 5338 0 _0191_
rlabel metal2 21850 8296 21850 8296 0 _0192_
rlabel metal1 16882 13226 16882 13226 0 _0193_
rlabel metal1 16836 18938 16836 18938 0 _0194_
rlabel metal1 15916 18938 15916 18938 0 _0195_
rlabel metal1 18860 15674 18860 15674 0 _0196_
rlabel metal1 20562 17544 20562 17544 0 _0197_
rlabel metal1 13524 20978 13524 20978 0 _0198_
rlabel metal1 21620 16762 21620 16762 0 _0199_
rlabel metal2 10994 17544 10994 17544 0 _0200_
rlabel metal1 13662 17238 13662 17238 0 _0201_
rlabel metal1 13708 16422 13708 16422 0 _0202_
rlabel metal2 12926 16082 12926 16082 0 _0203_
rlabel metal1 9476 12818 9476 12818 0 _0204_
rlabel metal1 16100 15130 16100 15130 0 _0205_
rlabel metal2 16974 14144 16974 14144 0 _0206_
rlabel metal1 19734 14892 19734 14892 0 _0207_
rlabel metal1 19596 17850 19596 17850 0 _0208_
rlabel metal1 16606 14518 16606 14518 0 _0209_
rlabel metal1 20470 12274 20470 12274 0 _0210_
rlabel metal1 19504 16490 19504 16490 0 _0211_
rlabel metal1 19412 14586 19412 14586 0 _0212_
rlabel metal1 22218 19244 22218 19244 0 _0213_
rlabel metal1 16422 19924 16422 19924 0 _0214_
rlabel metal1 18262 14586 18262 14586 0 _0215_
rlabel metal1 20930 19244 20930 19244 0 _0216_
rlabel metal2 18446 19108 18446 19108 0 _0217_
rlabel metal1 8234 16694 8234 16694 0 _0218_
rlabel metal1 9154 20978 9154 20978 0 _0219_
rlabel metal1 10442 18802 10442 18802 0 _0220_
rlabel metal1 8441 16422 8441 16422 0 _0221_
rlabel metal1 9890 19924 9890 19924 0 _0222_
rlabel metal1 11270 17748 11270 17748 0 _0223_
rlabel metal1 18952 5882 18952 5882 0 _0224_
rlabel metal2 21022 10268 21022 10268 0 _0225_
rlabel metal1 18078 12750 18078 12750 0 _0226_
rlabel metal1 19228 7514 19228 7514 0 _0227_
rlabel metal2 20838 8092 20838 8092 0 _0228_
rlabel metal1 16698 13396 16698 13396 0 _0229_
rlabel metal2 12466 16354 12466 16354 0 _0230_
rlabel metal2 13202 15844 13202 15844 0 _0231_
rlabel metal1 14122 14858 14122 14858 0 _0232_
rlabel metal1 13018 15368 13018 15368 0 _0233_
rlabel metal1 8832 14450 8832 14450 0 _0234_
rlabel metal1 14352 12818 14352 12818 0 _0235_
rlabel via1 18906 20485 18906 20485 0 _0236_
rlabel metal1 21505 20978 21505 20978 0 _0237_
rlabel metal1 11454 16116 11454 16116 0 _0238_
rlabel metal1 14904 18326 14904 18326 0 _0239_
rlabel metal2 20930 20060 20930 20060 0 _0240_
rlabel metal1 15502 14042 15502 14042 0 _0241_
rlabel metal1 8694 19312 8694 19312 0 _0242_
rlabel metal1 13754 22474 13754 22474 0 _0243_
rlabel metal1 14260 14042 14260 14042 0 _0244_
rlabel metal1 15042 14586 15042 14586 0 _0245_
rlabel metal1 11684 20978 11684 20978 0 _0246_
rlabel metal1 14720 16014 14720 16014 0 _0247_
rlabel metal2 12190 20910 12190 20910 0 _0248_
rlabel metal1 13202 19244 13202 19244 0 _0249_
rlabel metal1 24794 13192 24794 13192 0 _0250_
rlabel metal1 10810 19754 10810 19754 0 _0251_
rlabel metal1 11868 19278 11868 19278 0 _0252_
rlabel via1 22034 19771 22034 19771 0 _0253_
rlabel metal2 7774 14484 7774 14484 0 _0254_
rlabel metal2 8418 15334 8418 15334 0 _0255_
rlabel metal1 9522 17068 9522 17068 0 _0256_
rlabel metal2 7222 14722 7222 14722 0 _0257_
rlabel metal1 11914 15572 11914 15572 0 _0258_
rlabel metal1 8188 16626 8188 16626 0 _0259_
rlabel metal2 19642 24378 19642 24378 0 _0260_
rlabel metal1 17986 24174 17986 24174 0 _0261_
rlabel via2 14674 18173 14674 18173 0 _0262_
rlabel metal2 19366 24446 19366 24446 0 _0263_
rlabel metal2 18262 24140 18262 24140 0 _0264_
rlabel metal1 16560 23222 16560 23222 0 _0265_
rlabel metal1 16790 20502 16790 20502 0 _0266_
rlabel metal1 16744 17850 16744 17850 0 _0267_
rlabel metal1 16606 23698 16606 23698 0 _0268_
rlabel metal1 15732 21930 15732 21930 0 _0269_
rlabel metal1 16882 14586 16882 14586 0 _0270_
rlabel metal1 17526 24242 17526 24242 0 _0271_
rlabel metal2 23782 11424 23782 11424 0 _0272_
rlabel metal1 21022 12852 21022 12852 0 _0273_
rlabel metal1 20286 14586 20286 14586 0 _0274_
rlabel metal2 22494 10370 22494 10370 0 _0275_
rlabel metal1 20148 12614 20148 12614 0 _0276_
rlabel metal2 22126 15300 22126 15300 0 _0277_
rlabel metal1 23414 12920 23414 12920 0 _0278_
rlabel metal2 23322 16932 23322 16932 0 _0279_
rlabel metal1 20378 10778 20378 10778 0 _0280_
rlabel metal1 24196 10710 24196 10710 0 _0281_
rlabel metal1 22494 17170 22494 17170 0 _0282_
rlabel metal1 22770 8942 22770 8942 0 _0283_
rlabel metal2 16698 23358 16698 23358 0 _0284_
rlabel metal1 17204 22474 17204 22474 0 _0285_
rlabel metal2 18998 25228 18998 25228 0 _0286_
rlabel metal1 16100 24242 16100 24242 0 _0287_
rlabel metal1 17388 20026 17388 20026 0 _0288_
rlabel metal2 15870 24140 15870 24140 0 _0289_
rlabel via2 17250 20859 17250 20859 0 _0290_
rlabel metal2 18722 19618 18722 19618 0 _0291_
rlabel metal2 21850 22406 21850 22406 0 _0292_
rlabel metal1 16560 22406 16560 22406 0 _0293_
rlabel metal1 19182 18156 19182 18156 0 _0294_
rlabel metal1 20608 23154 20608 23154 0 _0295_
rlabel metal1 24702 11322 24702 11322 0 _0296_
rlabel metal2 23322 15708 23322 15708 0 _0297_
rlabel metal2 22218 14076 22218 14076 0 _0298_
rlabel metal1 24472 10234 24472 10234 0 _0299_
rlabel metal1 24196 14926 24196 14926 0 _0300_
rlabel metal1 23414 13362 23414 13362 0 _0301_
rlabel metal2 19090 6562 19090 6562 0 _0302_
rlabel metal2 23046 13532 23046 13532 0 _0303_
rlabel metal1 24472 8602 24472 8602 0 _0304_
rlabel metal2 16790 5304 16790 5304 0 _0305_
rlabel metal1 25070 12886 25070 12886 0 _0306_
rlabel metal1 24288 7310 24288 7310 0 _0307_
rlabel metal2 24242 14246 24242 14246 0 _0308_
rlabel metal1 24564 14994 24564 14994 0 _0309_
rlabel metal1 24932 12750 24932 12750 0 _0310_
rlabel metal2 25346 11560 25346 11560 0 _0311_
rlabel metal1 25944 14450 25944 14450 0 _0312_
rlabel metal2 25346 10404 25346 10404 0 _0313_
rlabel metal2 19274 9112 19274 9112 0 _0314_
rlabel metal1 10718 17204 10718 17204 0 _0315_
rlabel metal1 14858 7718 14858 7718 0 _0316_
rlabel metal1 12006 13940 12006 13940 0 _0317_
rlabel metal1 20792 15130 20792 15130 0 _0318_
rlabel metal1 14490 17578 14490 17578 0 _0319_
rlabel metal1 19504 14042 19504 14042 0 _0320_
rlabel metal1 14306 16660 14306 16660 0 _0321_
rlabel metal1 24380 9146 24380 9146 0 _0322_
rlabel metal1 21298 4794 21298 4794 0 _0323_
rlabel metal2 23874 8228 23874 8228 0 _0324_
rlabel metal1 19872 4114 19872 4114 0 _0325_
rlabel metal2 9430 11492 9430 11492 0 _0326_
rlabel metal2 15318 20196 15318 20196 0 _0327_
rlabel metal1 13294 14008 13294 14008 0 _0328_
rlabel metal2 13938 19074 13938 19074 0 _0329_
rlabel metal1 12926 22950 12926 22950 0 _0330_
rlabel metal1 20654 21420 20654 21420 0 _0331_
rlabel metal1 13800 22406 13800 22406 0 _0332_
rlabel metal1 19136 21114 19136 21114 0 _0333_
rlabel metal1 16606 8602 16606 8602 0 _0334_
rlabel metal1 9292 14042 9292 14042 0 _0335_
rlabel metal2 13018 7650 13018 7650 0 _0336_
rlabel metal2 11086 15504 11086 15504 0 _0337_
rlabel metal1 10626 21624 10626 21624 0 _0338_
rlabel metal1 9522 18700 9522 18700 0 _0339_
rlabel metal1 10212 22406 10212 22406 0 _0340_
rlabel metal1 8004 18938 8004 18938 0 _0341_
rlabel metal2 19458 9520 19458 9520 0 _0342_
rlabel metal1 18676 9146 18676 9146 0 _0343_
rlabel metal1 17066 7480 17066 7480 0 _0344_
rlabel metal2 19918 6817 19918 6817 0 _0345_
rlabel metal2 12558 7344 12558 7344 0 _0346_
rlabel metal1 9568 9146 9568 9146 0 _0347_
rlabel metal2 15870 10914 15870 10914 0 _0348_
rlabel metal1 9062 12716 9062 12716 0 _0349_
rlabel metal1 16928 10710 16928 10710 0 _0350_
rlabel metal1 9890 13498 9890 13498 0 _0351_
rlabel metal1 12834 13294 12834 13294 0 _0352_
rlabel via2 9338 12291 9338 12291 0 _0353_
rlabel metal1 22908 10234 22908 10234 0 _0354_
rlabel metal1 15502 21624 15502 21624 0 _0355_
rlabel metal1 22034 11322 22034 11322 0 _0356_
rlabel metal1 19136 20230 19136 20230 0 _0357_
rlabel metal2 18262 8942 18262 8942 0 _0358_
rlabel metal1 20079 4658 20079 4658 0 _0359_
rlabel metal1 19642 5338 19642 5338 0 _0360_
rlabel metal1 18676 2074 18676 2074 0 _0361_
rlabel metal2 20378 16354 20378 16354 0 _0362_
rlabel metal1 8878 11832 8878 11832 0 _0363_
rlabel metal1 18860 12954 18860 12954 0 _0364_
rlabel metal1 9890 14586 9890 14586 0 _0365_
rlabel metal2 20930 23902 20930 23902 0 _0366_
rlabel metal1 20838 22508 20838 22508 0 _0367_
rlabel metal2 22126 23256 22126 23256 0 _0368_
rlabel metal2 22402 23630 22402 23630 0 _0369_
rlabel metal1 13386 20536 13386 20536 0 _0370_
rlabel metal1 13432 13158 13432 13158 0 _0371_
rlabel metal1 12742 18632 12742 18632 0 _0372_
rlabel metal1 10028 8058 10028 8058 0 _0373_
rlabel metal1 20976 18394 20976 18394 0 _0374_
rlabel metal1 15732 13158 15732 13158 0 _0375_
rlabel metal2 20286 18632 20286 18632 0 _0376_
rlabel metal1 12098 15130 12098 15130 0 _0377_
rlabel via2 37490 6205 37490 6205 0 ccff_head
rlabel via2 38226 33371 38226 33371 0 ccff_tail
rlabel metal1 22724 37230 22724 37230 0 chanx_left_in[0]
rlabel metal1 37766 36142 37766 36142 0 chanx_left_in[10]
rlabel metal3 1234 12308 1234 12308 0 chanx_left_in[11]
rlabel metal2 34822 1588 34822 1588 0 chanx_left_in[12]
rlabel metal3 1234 36788 1234 36788 0 chanx_left_in[13]
rlabel metal1 38180 36754 38180 36754 0 chanx_left_in[14]
rlabel metal2 29026 1588 29026 1588 0 chanx_left_in[15]
rlabel metal3 1050 7548 1050 7548 0 chanx_left_in[16]
rlabel metal3 1234 30668 1234 30668 0 chanx_left_in[17]
rlabel metal3 4025 12580 4025 12580 0 chanx_left_in[18]
rlabel metal3 1740 38148 1740 38148 0 chanx_left_in[1]
rlabel metal2 4554 823 4554 823 0 chanx_left_in[2]
rlabel metal3 1234 20468 1234 20468 0 chanx_left_in[3]
rlabel metal3 1234 17748 1234 17748 0 chanx_left_in[4]
rlabel metal2 38318 28883 38318 28883 0 chanx_left_in[5]
rlabel metal1 18216 37230 18216 37230 0 chanx_left_in[6]
rlabel metal2 33534 1588 33534 1588 0 chanx_left_in[7]
rlabel metal3 1234 25228 1234 25228 0 chanx_left_in[8]
rlabel metal3 1234 32028 1234 32028 0 chanx_left_in[9]
rlabel metal3 1234 27268 1234 27268 0 chanx_left_out[0]
rlabel metal2 22586 1520 22586 1520 0 chanx_left_out[10]
rlabel metal1 14260 3366 14260 3366 0 chanx_left_out[11]
rlabel metal2 39330 1520 39330 1520 0 chanx_left_out[12]
rlabel metal3 1740 1428 1740 1428 0 chanx_left_out[13]
rlabel metal2 38226 20621 38226 20621 0 chanx_left_out[14]
rlabel metal1 24656 37094 24656 37094 0 chanx_left_out[15]
rlabel metal1 14030 37094 14030 37094 0 chanx_left_out[16]
rlabel metal2 38226 36941 38226 36941 0 chanx_left_out[17]
rlabel metal2 16790 1520 16790 1520 0 chanx_left_out[18]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[1]
rlabel metal2 38226 34833 38226 34833 0 chanx_left_out[2]
rlabel metal1 15640 37094 15640 37094 0 chanx_left_out[3]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[4]
rlabel metal2 38226 12461 38226 12461 0 chanx_left_out[5]
rlabel metal1 16928 37094 16928 37094 0 chanx_left_out[6]
rlabel metal1 10488 37094 10488 37094 0 chanx_left_out[7]
rlabel metal2 25806 1520 25806 1520 0 chanx_left_out[8]
rlabel metal1 9522 2822 9522 2822 0 chanx_left_out[9]
rlabel metal2 38318 30107 38318 30107 0 chany_top_in[0]
rlabel metal2 38042 1367 38042 1367 0 chany_top_in[10]
rlabel metal2 38318 15895 38318 15895 0 chany_top_in[11]
rlabel metal1 29486 37230 29486 37230 0 chany_top_in[12]
rlabel metal1 12512 37230 12512 37230 0 chany_top_in[13]
rlabel metal1 37766 4114 37766 4114 0 chany_top_in[14]
rlabel metal2 38318 32215 38318 32215 0 chany_top_in[15]
rlabel metal1 36846 37230 36846 37230 0 chany_top_in[16]
rlabel metal1 21758 37230 21758 37230 0 chany_top_in[17]
rlabel metal3 1234 19108 1234 19108 0 chany_top_in[18]
rlabel metal2 38318 7701 38318 7701 0 chany_top_in[1]
rlabel metal3 1234 22508 1234 22508 0 chany_top_in[2]
rlabel metal3 1050 2788 1050 2788 0 chany_top_in[3]
rlabel metal1 25944 37230 25944 37230 0 chany_top_in[4]
rlabel metal3 1234 28628 1234 28628 0 chany_top_in[5]
rlabel metal2 30314 1588 30314 1588 0 chany_top_in[6]
rlabel metal1 33672 37230 33672 37230 0 chany_top_in[7]
rlabel metal3 1234 9588 1234 9588 0 chany_top_in[8]
rlabel metal2 2622 1350 2622 1350 0 chany_top_in[9]
rlabel metal1 11362 2822 11362 2822 0 chany_top_out[0]
rlabel metal2 36110 1520 36110 1520 0 chany_top_out[10]
rlabel via2 38226 17051 38226 17051 0 chany_top_out[11]
rlabel metal2 38226 11101 38226 11101 0 chany_top_out[12]
rlabel metal3 1234 6188 1234 6188 0 chany_top_out[13]
rlabel metal3 1234 33388 1234 33388 0 chany_top_out[14]
rlabel via2 38226 2805 38226 2805 0 chany_top_out[15]
rlabel metal1 4738 37094 4738 37094 0 chany_top_out[16]
rlabel metal2 38226 14297 38226 14297 0 chany_top_out[17]
rlabel metal2 38226 25177 38226 25177 0 chany_top_out[18]
rlabel metal2 31602 1520 31602 1520 0 chany_top_out[1]
rlabel via2 38226 27285 38226 27285 0 chany_top_out[2]
rlabel metal1 6302 37094 6302 37094 0 chany_top_out[3]
rlabel metal3 1234 23868 1234 23868 0 chany_top_out[4]
rlabel metal2 19366 1520 19366 1520 0 chany_top_out[5]
rlabel metal2 46 2880 46 2880 0 chany_top_out[6]
rlabel metal2 23874 1520 23874 1520 0 chany_top_out[7]
rlabel metal1 7912 37094 7912 37094 0 chany_top_out[8]
rlabel metal1 20148 37094 20148 37094 0 chany_top_out[9]
rlabel metal1 1656 6698 1656 6698 0 clknet_0_prog_clk
rlabel metal2 1610 2992 1610 2992 0 clknet_3_0__leaf_prog_clk
rlabel metal1 6578 6358 6578 6358 0 clknet_3_1__leaf_prog_clk
rlabel metal1 3542 7786 3542 7786 0 clknet_3_2__leaf_prog_clk
rlabel metal2 6762 7650 6762 7650 0 clknet_3_3__leaf_prog_clk
rlabel metal1 13294 4012 13294 4012 0 clknet_3_4__leaf_prog_clk
rlabel metal1 12972 5134 12972 5134 0 clknet_3_5__leaf_prog_clk
rlabel metal1 8694 10098 8694 10098 0 clknet_3_6__leaf_prog_clk
rlabel metal2 14306 7412 14306 7412 0 clknet_3_7__leaf_prog_clk
rlabel metal1 1794 12172 1794 12172 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 2990 37230 2990 37230 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5842 1761 5842 1761 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 1334 1860 1334 1860 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 34960 37230 34960 37230 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 27876 37230 27876 37230 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 18078 1761 18078 1761 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 37674 36788 37674 36788 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 38318 4369 38318 4369 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 1564 37230 1564 37230 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 14674 14365 14674 14365 0 mem_left_track_1.DFFR_0_.D
rlabel metal1 8924 19822 8924 19822 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 8234 20400 8234 20400 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 9522 10982 9522 10982 0 mem_left_track_11.DFFR_0_.D
rlabel metal1 21758 9112 21758 9112 0 mem_left_track_11.DFFR_0_.Q
rlabel metal2 16882 9928 16882 9928 0 mem_left_track_11.DFFR_1_.Q
rlabel metal1 15640 18870 15640 18870 0 mem_left_track_13.DFFR_0_.Q
rlabel metal1 14260 6426 14260 6426 0 mem_left_track_13.DFFR_1_.Q
rlabel metal1 20332 20978 20332 20978 0 mem_left_track_15.DFFR_0_.Q
rlabel metal2 13294 6256 13294 6256 0 mem_left_track_15.DFFR_1_.Q
rlabel metal1 18630 13362 18630 13362 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 14490 10234 14490 10234 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 16054 10778 16054 10778 0 mem_left_track_19.DFFR_0_.Q
rlabel metal2 8234 11271 8234 11271 0 mem_left_track_19.DFFR_1_.Q
rlabel metal1 7038 12818 7038 12818 0 mem_left_track_21.DFFR_0_.Q
rlabel metal2 13754 6596 13754 6596 0 mem_left_track_21.DFFR_1_.Q
rlabel metal1 7866 13294 7866 13294 0 mem_left_track_23.DFFR_0_.Q
rlabel metal2 7498 10897 7498 10897 0 mem_left_track_23.DFFR_1_.Q
rlabel metal1 18078 20332 18078 20332 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 15962 2315 15962 2315 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 13800 2618 13800 2618 0 mem_left_track_27.DFFR_0_.Q
rlabel metal1 20286 8976 20286 8976 0 mem_left_track_27.DFFR_1_.Q
rlabel metal1 8602 8840 8602 8840 0 mem_left_track_29.DFFR_0_.Q
rlabel metal1 14398 2346 14398 2346 0 mem_left_track_29.DFFR_1_.Q
rlabel metal2 10718 13209 10718 13209 0 mem_left_track_3.DFFR_0_.Q
rlabel metal1 7360 13294 7360 13294 0 mem_left_track_3.DFFR_1_.Q
rlabel metal3 16629 2652 16629 2652 0 mem_left_track_31.DFFR_0_.Q
rlabel metal2 16928 17204 16928 17204 0 mem_left_track_31.DFFR_1_.Q
rlabel metal2 17158 3145 17158 3145 0 mem_left_track_33.DFFR_0_.Q
rlabel via2 12466 2805 12466 2805 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 13616 4046 13616 4046 0 mem_left_track_35.DFFR_0_.Q
rlabel metal1 18354 16422 18354 16422 0 mem_left_track_35.DFFR_1_.Q
rlabel metal1 18124 9690 18124 9690 0 mem_left_track_37.DFFR_0_.Q
rlabel metal1 15870 23052 15870 23052 0 mem_left_track_5.DFFR_0_.Q
rlabel via2 17434 22627 17434 22627 0 mem_left_track_5.DFFR_1_.Q
rlabel metal1 14858 18734 14858 18734 0 mem_left_track_7.DFFR_0_.Q
rlabel via1 13202 21675 13202 21675 0 mem_left_track_7.DFFR_1_.Q
rlabel metal1 19550 12852 19550 12852 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 16146 9486 16146 9486 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 8970 11118 8970 11118 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 15962 14093 15962 14093 0 mem_top_track_10.DFFR_0_.D
rlabel metal2 18354 19686 18354 19686 0 mem_top_track_10.DFFR_0_.Q
rlabel metal2 8418 6086 8418 6086 0 mem_top_track_10.DFFR_1_.Q
rlabel metal1 1886 5576 1886 5576 0 mem_top_track_12.DFFR_0_.Q
rlabel metal1 6118 16082 6118 16082 0 mem_top_track_12.DFFR_1_.Q
rlabel metal1 19964 11118 19964 11118 0 mem_top_track_14.DFFR_0_.Q
rlabel metal1 20102 7344 20102 7344 0 mem_top_track_14.DFFR_1_.Q
rlabel via2 13386 12189 13386 12189 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 8326 14994 8326 14994 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 21114 20672 21114 20672 0 mem_top_track_18.DFFR_0_.Q
rlabel metal2 12650 18751 12650 18751 0 mem_top_track_18.DFFR_1_.Q
rlabel metal2 17342 11934 17342 11934 0 mem_top_track_2.DFFR_0_.Q
rlabel metal1 10159 10234 10159 10234 0 mem_top_track_2.DFFR_1_.Q
rlabel metal1 8326 13906 8326 13906 0 mem_top_track_20.DFFR_0_.Q
rlabel metal1 14628 7786 14628 7786 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 16192 8058 16192 8058 0 mem_top_track_22.DFFR_0_.Q
rlabel metal1 19412 13294 19412 13294 0 mem_top_track_22.DFFR_1_.Q
rlabel metal1 15548 8262 15548 8262 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 16146 9894 16146 9894 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 13294 18870 13294 18870 0 mem_top_track_26.DFFR_0_.Q
rlabel metal2 14582 5542 14582 5542 0 mem_top_track_26.DFFR_1_.Q
rlabel metal1 18630 20910 18630 20910 0 mem_top_track_28.DFFR_0_.Q
rlabel metal1 16008 3638 16008 3638 0 mem_top_track_28.DFFR_1_.Q
rlabel metal1 7498 14994 7498 14994 0 mem_top_track_30.DFFR_0_.Q
rlabel metal2 12926 6681 12926 6681 0 mem_top_track_30.DFFR_1_.Q
rlabel metal2 1886 3740 1886 3740 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 7222 21318 7222 21318 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 9338 9112 9338 9112 0 mem_top_track_34.DFFR_0_.Q
rlabel metal1 13110 7446 13110 7446 0 mem_top_track_34.DFFR_1_.Q
rlabel metal1 12742 14280 12742 14280 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 19090 14960 19090 14960 0 mem_top_track_4.DFFR_0_.Q
rlabel metal1 13294 1972 13294 1972 0 mem_top_track_4.DFFR_1_.Q
rlabel metal2 1886 2176 1886 2176 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 4968 2482 4968 2482 0 mem_top_track_6.DFFR_1_.Q
rlabel metal1 19550 16626 19550 16626 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 32430 22508 32430 22508 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 24564 12818 24564 12818 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 9384 17102 9384 17102 0 mux_left_track_1.INVTX1_2_.out
rlabel metal2 12466 20060 12466 20060 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12374 19924 12374 19924 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12558 20094 12558 20094 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 5566 23222 5566 23222 0 mux_left_track_1.out
rlabel metal1 25162 6766 25162 6766 0 mux_left_track_11.INVTX1_0_.out
rlabel metal2 20470 11424 20470 11424 0 mux_left_track_11.INVTX1_1_.out
rlabel metal1 21850 17170 21850 17170 0 mux_left_track_11.INVTX1_2_.out
rlabel metal2 22126 10098 22126 10098 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23460 16966 23460 16966 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23552 12750 23552 12750 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 37536 12206 37536 12206 0 mux_left_track_11.out
rlabel metal1 14996 33286 14996 33286 0 mux_left_track_13.INVTX1_0_.out
rlabel metal1 15042 18666 15042 18666 0 mux_left_track_13.INVTX1_2_.out
rlabel metal1 16560 24174 16560 24174 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17342 22644 17342 22644 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16744 24378 16744 24378 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16974 28730 16974 28730 0 mux_left_track_13.out
rlabel metal1 19918 23222 19918 23222 0 mux_left_track_15.INVTX1_0_.out
rlabel metal1 20010 13838 20010 13838 0 mux_left_track_15.INVTX1_2_.out
rlabel metal1 17710 21454 17710 21454 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19688 20026 19688 20026 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17618 21284 17618 21284 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14030 33898 14030 33898 0 mux_left_track_15.out
rlabel metal2 33166 14280 33166 14280 0 mux_left_track_17.INVTX1_0_.out
rlabel metal2 24610 14620 24610 14620 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 23138 13498 23138 13498 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23690 15334 23690 15334 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24426 12342 24426 12342 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 23414 6290 23414 6290 0 mux_left_track_17.out
rlabel metal2 31970 6052 31970 6052 0 mux_left_track_19.INVTX1_0_.out
rlabel metal1 18538 5032 18538 5032 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22494 14008 22494 14008 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20654 5508 20654 5508 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 21298 5644 21298 5644 0 mux_left_track_19.out
rlabel metal1 8832 12750 8832 12750 0 mux_left_track_21.INVTX1_0_.out
rlabel metal2 10626 11305 10626 11305 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19918 6052 19918 6052 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25070 3502 25070 3502 0 mux_left_track_21.out
rlabel metal1 5382 8398 5382 8398 0 mux_left_track_23.INVTX1_0_.out
rlabel metal2 12466 17952 12466 17952 0 mux_left_track_23.INVTX1_1_.out
rlabel metal1 10672 12342 10672 12342 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17158 7344 17158 7344 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16606 3978 16606 3978 0 mux_left_track_23.out
rlabel metal1 24518 22066 24518 22066 0 mux_left_track_25.INVTX1_0_.out
rlabel metal2 16882 26316 16882 26316 0 mux_left_track_25.INVTX1_1_.out
rlabel metal2 21390 17340 21390 17340 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23368 12682 23368 12682 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 36938 3196 36938 3196 0 mux_left_track_25.out
rlabel metal2 19320 2652 19320 2652 0 mux_left_track_27.INVTX1_0_.out
rlabel metal1 16882 15980 16882 15980 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 18446 2618 18446 2618 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel via2 1610 13923 1610 13923 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2346 12818 2346 12818 0 mux_left_track_27.out
rlabel metal1 11040 16626 11040 16626 0 mux_left_track_29.INVTX1_0_.out
rlabel metal1 12788 11662 12788 11662 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20792 16694 20792 16694 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 33442 18564 33442 18564 0 mux_left_track_29.out
rlabel metal2 9154 17068 9154 17068 0 mux_left_track_3.INVTX1_0_.out
rlabel metal2 9706 16864 9706 16864 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12052 15606 12052 15606 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 9798 15232 9798 15232 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 5014 14586 5014 14586 0 mux_left_track_3.out
rlabel metal1 22862 33286 22862 33286 0 mux_left_track_31.INVTX1_0_.out
rlabel metal1 21114 22984 21114 22984 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22586 26452 22586 26452 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 22862 29274 22862 29274 0 mux_left_track_31.out
rlabel metal1 9936 8942 9936 8942 0 mux_left_track_33.INVTX1_0_.out
rlabel metal1 12558 18768 12558 18768 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13846 19584 13846 19584 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14076 33966 14076 33966 0 mux_left_track_33.out
rlabel metal2 9062 18972 9062 18972 0 mux_left_track_35.INVTX1_0_.out
rlabel metal1 19757 18190 19757 18190 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20838 18564 20838 18564 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30544 31790 30544 31790 0 mux_left_track_35.out
rlabel metal2 33718 9554 33718 9554 0 mux_left_track_37.INVTX1_0_.out
rlabel metal1 24610 11662 24610 11662 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 24426 14314 24426 14314 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24518 11594 24518 11594 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 20378 8398 20378 8398 0 mux_left_track_37.out
rlabel metal1 18906 32198 18906 32198 0 mux_left_track_5.INVTX1_0_.out
rlabel metal1 15594 18394 15594 18394 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19228 24106 19228 24106 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19918 23800 19918 23800 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31786 28900 31786 28900 0 mux_left_track_5.out
rlabel metal1 17158 24276 17158 24276 0 mux_left_track_7.INVTX1_0_.out
rlabel metal1 16422 23494 16422 23494 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17710 17782 17710 17782 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16928 32402 16928 32402 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 15962 34340 15962 34340 0 mux_left_track_7.out
rlabel metal2 33350 21454 33350 21454 0 mux_left_track_9.INVTX1_0_.out
rlabel metal1 21620 15334 21620 15334 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21160 11866 21160 11866 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25024 11050 25024 11050 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 28934 10540 28934 10540 0 mux_left_track_9.out
rlabel via2 15318 13277 15318 13277 0 mux_top_track_0.INVTX1_0_.out
rlabel metal2 17618 13634 17618 13634 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 20102 18190 20102 18190 0 mux_top_track_0.INVTX1_2_.out
rlabel metal2 15870 13634 15870 13634 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17066 16966 17066 16966 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16560 12614 16560 12614 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17664 11050 17664 11050 0 mux_top_track_0.out
rlabel metal1 19320 19278 19320 19278 0 mux_top_track_10.INVTX1_0_.out
rlabel via2 16238 19907 16238 19907 0 mux_top_track_10.INVTX1_1_.out
rlabel metal1 31832 32742 31832 32742 0 mux_top_track_10.INVTX1_2_.out
rlabel metal1 17894 19686 17894 19686 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21114 19346 21114 19346 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19596 17034 19596 17034 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 18998 5032 18998 5032 0 mux_top_track_10.out
rlabel metal1 14260 19278 14260 19278 0 mux_top_track_12.INVTX1_1_.out
rlabel metal1 9752 19890 9752 19890 0 mux_top_track_12.INVTX1_2_.out
rlabel metal2 11730 18224 11730 18224 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10534 20026 10534 20026 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 10166 17714 10166 17714 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 2438 11900 2438 11900 0 mux_top_track_12.out
rlabel metal2 21022 7072 21022 7072 0 mux_top_track_14.INVTX1_1_.out
rlabel metal1 26496 6970 26496 6970 0 mux_top_track_14.INVTX1_2_.out
rlabel metal2 18078 12920 18078 12920 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21390 8058 21390 8058 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 18722 7582 18722 7582 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel via2 13662 2907 13662 2907 0 mux_top_track_14.out
rlabel metal1 13800 14926 13800 14926 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 9062 14382 9062 14382 0 mux_top_track_16.INVTX1_2_.out
rlabel metal2 14306 15232 14306 15232 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12006 16626 12006 16626 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 13156 15538 13156 15538 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 10902 32878 10902 32878 0 mux_top_track_16.out
rlabel metal2 32246 25874 32246 25874 0 mux_top_track_18.INVTX1_2_.out
rlabel via1 16698 16218 16698 16218 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21068 20026 21068 20026 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 19366 19567 19366 19567 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 19550 33490 19550 33490 0 mux_top_track_18.out
rlabel metal1 16100 16558 16100 16558 0 mux_top_track_2.INVTX1_1_.out
rlabel metal2 17342 8636 17342 8636 0 mux_top_track_2.INVTX1_2_.out
rlabel metal1 17710 13430 17710 13430 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17342 7582 17342 7582 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18308 7786 18308 7786 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 26542 6222 26542 6222 0 mux_top_track_2.out
rlabel metal1 9292 17714 9292 17714 0 mux_top_track_20.INVTX1_1_.out
rlabel metal2 12466 14178 12466 14178 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19458 9452 19458 9452 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30452 5678 30452 5678 0 mux_top_track_20.out
rlabel metal2 13110 19652 13110 19652 0 mux_top_track_22.INVTX1_1_.out
rlabel metal2 16606 17068 16606 17068 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21482 15912 21482 15912 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33810 16524 33810 16524 0 mux_top_track_22.out
rlabel metal1 18998 16014 18998 16014 0 mux_top_track_24.INVTX1_0_.out
rlabel metal1 26542 4794 26542 4794 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 21091 5814 21091 5814 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25714 9622 25714 9622 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 35098 9826 35098 9826 0 mux_top_track_24.out
rlabel metal1 18262 18700 18262 18700 0 mux_top_track_26.INVTX1_0_.out
rlabel metal1 16054 32742 16054 32742 0 mux_top_track_26.INVTX1_1_.out
rlabel metal2 15962 17374 15962 17374 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14306 15538 14306 15538 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 2898 8636 2898 8636 0 mux_top_track_26.out
rlabel metal2 31786 23358 31786 23358 0 mux_top_track_28.INVTX1_1_.out
rlabel metal1 18262 21318 18262 21318 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13754 21896 13754 21896 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 10166 27302 10166 27302 0 mux_top_track_28.out
rlabel metal1 9016 15538 9016 15538 0 mux_top_track_30.INVTX1_1_.out
rlabel metal1 12650 8534 12650 8534 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17986 9724 17986 9724 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 38042 5916 38042 5916 0 mux_top_track_30.out
rlabel metal1 8924 18802 8924 18802 0 mux_top_track_32.INVTX1_1_.out
rlabel metal2 10350 19788 10350 19788 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 11086 20944 11086 20944 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8142 33966 8142 33966 0 mux_top_track_32.out
rlabel metal1 8418 11016 8418 11016 0 mux_top_track_34.INVTX1_1_.out
rlabel metal2 18354 8636 18354 8636 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19734 10098 19734 10098 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30958 12818 30958 12818 0 mux_top_track_34.out
rlabel metal1 9752 20774 9752 20774 0 mux_top_track_36.INVTX1_2_.out
rlabel metal2 15226 16456 15226 16456 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13708 21046 13708 21046 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16169 19822 16169 19822 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 33166 21692 33166 21692 0 mux_top_track_36.out
rlabel metal1 8694 25670 8694 25670 0 mux_top_track_4.INVTX1_2_.out
rlabel metal1 20792 17714 20792 17714 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15042 21114 15042 21114 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 21114 20502 21114 20502 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 28980 21998 28980 21998 0 mux_top_track_4.out
rlabel metal1 8648 12614 8648 12614 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 15042 17782 15042 17782 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12144 17102 12144 17102 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12558 31790 12558 31790 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 10028 36754 10028 36754 0 mux_top_track_6.out
rlabel metal1 20654 12172 20654 12172 0 mux_top_track_8.INVTX1_2_.out
rlabel metal1 18952 18938 18952 18938 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19780 15130 19780 15130 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17618 19040 17618 19040 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 8510 18513 8510 18513 0 mux_top_track_8.out
rlabel via2 37766 6307 37766 6307 0 net1
rlabel metal2 5566 28356 5566 28356 0 net10
rlabel metal1 17618 17204 17618 17204 0 net100
rlabel metal1 13846 7310 13846 7310 0 net101
rlabel metal1 15318 19482 15318 19482 0 net102
rlabel via2 11086 17493 11086 17493 0 net103
rlabel metal2 19642 14688 19642 14688 0 net104
rlabel metal1 21850 18802 21850 18802 0 net105
rlabel metal1 9384 20910 9384 20910 0 net106
rlabel metal1 20884 9690 20884 9690 0 net107
rlabel via1 12926 14467 12926 14467 0 net108
rlabel metal1 21390 20570 21390 20570 0 net109
rlabel metal2 20746 10285 20746 10285 0 net11
rlabel metal2 14398 21529 14398 21529 0 net110
rlabel metal2 13018 21488 13018 21488 0 net111
rlabel metal2 9798 15742 9798 15742 0 net112
rlabel metal1 18446 24242 18446 24242 0 net113
rlabel metal1 16974 19346 16974 19346 0 net114
rlabel metal2 20838 12988 20838 12988 0 net115
rlabel metal1 22908 16626 22908 16626 0 net116
rlabel metal1 17112 21658 17112 21658 0 net117
rlabel metal1 19504 18802 19504 18802 0 net118
rlabel metal2 23138 15776 23138 15776 0 net119
rlabel metal1 3818 37162 3818 37162 0 net12
rlabel metal2 23138 13566 23138 13566 0 net120
rlabel metal2 24058 15504 24058 15504 0 net121
rlabel metal1 18814 9486 18814 9486 0 net122
rlabel metal1 21436 16014 21436 16014 0 net123
rlabel metal1 23506 8602 23506 8602 0 net124
rlabel metal1 10856 11866 10856 11866 0 net125
rlabel metal1 13018 22066 13018 22066 0 net126
rlabel metal1 17802 10098 17802 10098 0 net127
rlabel metal1 10396 21590 10396 21590 0 net128
rlabel metal2 19550 10336 19550 10336 0 net129
rlabel metal1 2622 11220 2622 11220 0 net13
rlabel metal1 12052 5338 12052 5338 0 net130
rlabel metal2 15502 11050 15502 11050 0 net131
rlabel metal2 22954 11900 22954 11900 0 net132
rlabel metal2 19458 6987 19458 6987 0 net133
rlabel metal1 22034 16592 22034 16592 0 net134
rlabel metal1 21758 23630 21758 23630 0 net135
rlabel metal2 12282 20366 12282 20366 0 net136
rlabel metal1 20562 18632 20562 18632 0 net137
rlabel metal2 5842 20060 5842 20060 0 net14
rlabel metal2 5566 16762 5566 16762 0 net15
rlabel metal2 38134 27200 38134 27200 0 net16
rlabel metal1 17664 37094 17664 37094 0 net17
rlabel metal2 33626 3570 33626 3570 0 net18
rlabel metal1 5980 21522 5980 21522 0 net19
rlabel metal1 21528 37162 21528 37162 0 net2
rlabel metal1 4186 32198 4186 32198 0 net20
rlabel metal1 37352 30022 37352 30022 0 net21
rlabel metal2 33902 4148 33902 4148 0 net22
rlabel metal2 37030 15436 37030 15436 0 net23
rlabel metal2 24886 35156 24886 35156 0 net24
rlabel metal1 13294 33490 13294 33490 0 net25
rlabel metal1 37260 3978 37260 3978 0 net26
rlabel metal2 33258 29818 33258 29818 0 net27
rlabel metal1 36064 37094 36064 37094 0 net28
rlabel metal1 21252 37094 21252 37094 0 net29
rlabel metal1 37030 36006 37030 36006 0 net3
rlabel metal2 5198 18564 5198 18564 0 net30
rlabel metal2 34730 8262 34730 8262 0 net31
rlabel metal1 6348 19822 6348 19822 0 net32
rlabel metal1 2185 11594 2185 11594 0 net33
rlabel metal1 24656 37162 24656 37162 0 net34
rlabel metal1 2185 29274 2185 29274 0 net35
rlabel metal1 30130 2618 30130 2618 0 net36
rlabel metal1 33028 37094 33028 37094 0 net37
rlabel metal2 3726 9588 3726 9588 0 net38
rlabel metal2 1702 9996 1702 9996 0 net39
rlabel metal1 1610 12716 1610 12716 0 net4
rlabel metal2 1610 11968 1610 11968 0 net40
rlabel metal1 7314 29070 7314 29070 0 net41
rlabel metal3 14628 6256 14628 6256 0 net42
rlabel metal2 3358 3060 3358 3060 0 net43
rlabel metal1 33764 37162 33764 37162 0 net44
rlabel metal1 27738 37094 27738 37094 0 net45
rlabel metal1 13754 8364 13754 8364 0 net46
rlabel metal1 33396 36550 33396 36550 0 net47
rlabel metal1 36984 4794 36984 4794 0 net48
rlabel metal1 4048 36890 4048 36890 0 net49
rlabel metal1 32614 2550 32614 2550 0 net5
rlabel metal1 38088 21862 38088 21862 0 net50
rlabel metal1 7406 12954 7406 12954 0 net51
rlabel metal2 6578 13702 6578 13702 0 net52
rlabel metal2 37030 21930 37030 21930 0 net53
rlabel metal2 20102 3145 20102 3145 0 net54
rlabel metal1 31004 37162 31004 37162 0 net55
rlabel metal1 30130 37094 30130 37094 0 net56
rlabel metal2 4002 36958 4002 36958 0 net57
rlabel metal1 9246 37094 9246 37094 0 net58
rlabel metal1 22034 7344 22034 7344 0 net59
rlabel metal1 2162 36550 2162 36550 0 net6
rlabel metal2 4094 11271 4094 11271 0 net60
rlabel metal1 37950 33490 37950 33490 0 net61
rlabel metal2 4002 25636 4002 25636 0 net62
rlabel metal1 23276 2414 23276 2414 0 net63
rlabel metal2 12742 4522 12742 4522 0 net64
rlabel metal2 38042 2618 38042 2618 0 net65
rlabel metal1 2300 5202 2300 5202 0 net66
rlabel metal2 33626 19924 33626 19924 0 net67
rlabel metal1 23736 34714 23736 34714 0 net68
rlabel metal2 14306 35700 14306 35700 0 net69
rlabel metal2 38134 34714 38134 34714 0 net7
rlabel metal1 38042 37196 38042 37196 0 net70
rlabel metal1 16744 2414 16744 2414 0 net71
rlabel metal2 4830 15334 4830 15334 0 net72
rlabel metal2 33902 32980 33902 32980 0 net73
rlabel metal2 15778 36788 15778 36788 0 net74
rlabel metal2 34822 9418 34822 9418 0 net75
rlabel metal1 37950 12410 37950 12410 0 net76
rlabel metal2 16882 35972 16882 35972 0 net77
rlabel metal1 11868 34170 11868 34170 0 net78
rlabel metal1 25300 2414 25300 2414 0 net79
rlabel metal1 27370 8466 27370 8466 0 net8
rlabel metal2 13846 3145 13846 3145 0 net80
rlabel metal2 13202 5916 13202 5916 0 net81
rlabel metal1 36041 2414 36041 2414 0 net82
rlabel metal1 36294 17170 36294 17170 0 net83
rlabel metal2 36110 10676 36110 10676 0 net84
rlabel metal1 1702 6834 1702 6834 0 net85
rlabel metal1 2530 33490 2530 33490 0 net86
rlabel metal2 38042 4012 38042 4012 0 net87
rlabel metal1 5060 37230 5060 37230 0 net88
rlabel metal2 36478 13668 36478 13668 0 net89
rlabel metal1 3726 13430 3726 13430 0 net9
rlabel metal2 36938 24004 36938 24004 0 net90
rlabel metal2 32338 3706 32338 3706 0 net91
rlabel metal2 33534 25908 33534 25908 0 net92
rlabel metal2 6578 37060 6578 37060 0 net93
rlabel metal1 6578 21114 6578 21114 0 net94
rlabel metal1 19458 2380 19458 2380 0 net95
rlabel metal1 1564 6426 1564 6426 0 net96
rlabel metal1 13294 2516 13294 2516 0 net97
rlabel metal1 8832 33082 8832 33082 0 net98
rlabel metal1 19780 33626 19780 33626 0 net99
rlabel metal2 38134 21879 38134 21879 0 pReset
rlabel metal1 8142 8602 8142 8602 0 prog_clk
rlabel metal2 13570 2251 13570 2251 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal3 1234 14348 1234 14348 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 38318 24021 38318 24021 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21298 1860 21298 1860 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 32384 37230 32384 37230 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 30498 37230 30498 37230 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 3726 37230 3726 37230 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 9200 37230 9200 37230 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 27094 1588 27094 1588 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 10948 1234 10948 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
