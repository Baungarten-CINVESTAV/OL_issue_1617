// This is the unpowered netlist.
module cbx_1__0_ (bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_,
    bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_,
    vccd1,
    vssd1,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out);
 output bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
 output bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
 inout vccd1;
 inout vssd1;
 input [0:18] chanx_left_in;
 output [0:18] chanx_left_out;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire \mem_bottom_ipin_0.DFFR_0_.Q ;
 wire \mem_bottom_ipin_0.DFFR_1_.Q ;
 wire \mem_bottom_ipin_0.DFFR_2_.Q ;
 wire \mem_bottom_ipin_0.DFFR_3_.Q ;
 wire \mem_bottom_ipin_0.DFFR_4_.Q ;
 wire \mem_bottom_ipin_0.DFFR_5_.Q ;
 wire \mem_bottom_ipin_1.DFFR_0_.Q ;
 wire \mem_bottom_ipin_1.DFFR_1_.Q ;
 wire \mem_bottom_ipin_1.DFFR_2_.Q ;
 wire \mem_bottom_ipin_1.DFFR_3_.Q ;
 wire \mem_bottom_ipin_1.DFFR_4_.Q ;
 wire \mem_bottom_ipin_1.DFFR_5_.Q ;
 wire \mem_bottom_ipin_2.DFFR_0_.Q ;
 wire \mem_bottom_ipin_2.DFFR_1_.Q ;
 wire \mem_bottom_ipin_2.DFFR_2_.Q ;
 wire \mem_bottom_ipin_2.DFFR_3_.Q ;
 wire \mem_bottom_ipin_2.DFFR_4_.Q ;
 wire \mem_bottom_ipin_2.DFFR_5_.Q ;
 wire \mem_top_ipin_0.DFFR_0_.Q ;
 wire \mem_top_ipin_0.DFFR_1_.Q ;
 wire \mem_top_ipin_0.DFFR_2_.Q ;
 wire \mem_top_ipin_0.DFFR_3_.Q ;
 wire \mem_top_ipin_0.DFFR_4_.Q ;
 wire \mem_top_ipin_0.DFFR_5_.Q ;
 wire \mem_top_ipin_1.DFFR_0_.Q ;
 wire \mem_top_ipin_1.DFFR_1_.Q ;
 wire \mem_top_ipin_1.DFFR_2_.Q ;
 wire \mem_top_ipin_1.DFFR_3_.Q ;
 wire \mem_top_ipin_1.DFFR_4_.Q ;
 wire \mem_top_ipin_1.DFFR_5_.Q ;
 wire \mem_top_ipin_2.DFFR_0_.Q ;
 wire \mem_top_ipin_2.DFFR_1_.Q ;
 wire \mem_top_ipin_2.DFFR_2_.Q ;
 wire \mem_top_ipin_2.DFFR_3_.Q ;
 wire \mem_top_ipin_2.DFFR_4_.Q ;
 wire \mem_top_ipin_2.DFFR_5_.Q ;
 wire \mem_top_ipin_3.DFFR_0_.Q ;
 wire \mem_top_ipin_3.DFFR_1_.Q ;
 wire \mem_top_ipin_3.DFFR_2_.Q ;
 wire \mem_top_ipin_3.DFFR_3_.Q ;
 wire \mem_top_ipin_3.DFFR_4_.Q ;
 wire \mem_top_ipin_3.DFFR_5_.Q ;
 wire \mem_top_ipin_4.DFFR_0_.Q ;
 wire \mem_top_ipin_4.DFFR_1_.Q ;
 wire \mem_top_ipin_4.DFFR_2_.Q ;
 wire \mem_top_ipin_4.DFFR_3_.Q ;
 wire \mem_top_ipin_4.DFFR_4_.Q ;
 wire \mem_top_ipin_4.DFFR_5_.Q ;
 wire \mem_top_ipin_5.DFFR_0_.Q ;
 wire \mem_top_ipin_5.DFFR_1_.Q ;
 wire \mem_top_ipin_5.DFFR_2_.Q ;
 wire \mem_top_ipin_5.DFFR_3_.Q ;
 wire \mem_top_ipin_5.DFFR_4_.Q ;
 wire \mem_top_ipin_5.DFFR_5_.Q ;
 wire \mem_top_ipin_6.DFFR_0_.Q ;
 wire \mem_top_ipin_6.DFFR_1_.Q ;
 wire \mem_top_ipin_6.DFFR_2_.Q ;
 wire \mem_top_ipin_6.DFFR_3_.Q ;
 wire \mem_top_ipin_6.DFFR_4_.Q ;
 wire \mem_top_ipin_6.DFFR_5_.Q ;
 wire \mem_top_ipin_7.DFFR_0_.Q ;
 wire \mem_top_ipin_7.DFFR_1_.Q ;
 wire \mem_top_ipin_7.DFFR_2_.Q ;
 wire \mem_top_ipin_7.DFFR_3_.Q ;
 wire \mem_top_ipin_7.DFFR_4_.Q ;
 wire \mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \mux_bottom_ipin_0.INVTX1_2_.out ;
 wire \mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \mux_bottom_ipin_0.INVTX1_4_.out ;
 wire \mux_bottom_ipin_0.INVTX1_5_.out ;
 wire \mux_bottom_ipin_0.INVTX1_6_.out ;
 wire \mux_bottom_ipin_0.INVTX1_7_.out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_1.INVTX1_2_.out ;
 wire \mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \mux_bottom_ipin_1.INVTX1_4_.out ;
 wire \mux_bottom_ipin_1.INVTX1_5_.out ;
 wire \mux_bottom_ipin_1.INVTX1_6_.out ;
 wire \mux_bottom_ipin_1.INVTX1_7_.out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_0.INVTX1_2_.out ;
 wire \mux_top_ipin_0.INVTX1_3_.out ;
 wire \mux_top_ipin_0.INVTX1_4_.out ;
 wire \mux_top_ipin_0.INVTX1_5_.out ;
 wire \mux_top_ipin_0.INVTX1_6_.out ;
 wire \mux_top_ipin_0.INVTX1_7_.out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_1.INVTX1_2_.out ;
 wire \mux_top_ipin_1.INVTX1_3_.out ;
 wire \mux_top_ipin_1.INVTX1_4_.out ;
 wire \mux_top_ipin_1.INVTX1_5_.out ;
 wire \mux_top_ipin_1.INVTX1_6_.out ;
 wire \mux_top_ipin_1.INVTX1_7_.out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_2.INVTX1_2_.out ;
 wire \mux_top_ipin_2.INVTX1_3_.out ;
 wire \mux_top_ipin_2.INVTX1_6_.out ;
 wire \mux_top_ipin_2.INVTX1_7_.out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_5.INVTX1_4_.out ;
 wire \mux_top_ipin_5.INVTX1_5_.out ;
 wire \mux_top_ipin_5.INVTX1_6_.out ;
 wire \mux_top_ipin_5.INVTX1_7_.out ;
 wire \mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;

 sky130_fd_sc_hd__inv_2 _213_ (.A(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .Y(_199_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_201_));
 sky130_fd_sc_hd__inv_2 _215_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_198_));
 sky130_fd_sc_hd__inv_2 _216_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_197_));
 sky130_fd_sc_hd__inv_2 _217_ (.A(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .Y(_194_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .Y(_193_));
 sky130_fd_sc_hd__inv_2 _219_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_200_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_196_));
 sky130_fd_sc_hd__inv_2 _221_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_195_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(\mem_top_ipin_7.DFFR_3_.Q ),
    .Y(_189_));
 sky130_fd_sc_hd__inv_2 _223_ (.A(\mem_top_ipin_7.DFFR_0_.Q ),
    .Y(_192_));
 sky130_fd_sc_hd__inv_2 _224_ (.A(\mem_top_ipin_7.DFFR_2_.Q ),
    .Y(_188_));
 sky130_fd_sc_hd__inv_2 _225_ (.A(\mem_top_ipin_7.DFFR_1_.Q ),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(net49),
    .Y(_182_));
 sky130_fd_sc_hd__inv_2 _227_ (.A(\mem_top_ipin_7.DFFR_0_.Q ),
    .Y(_190_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(\mem_top_ipin_7.DFFR_2_.Q ),
    .Y(_184_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(\mem_top_ipin_7.DFFR_1_.Q ),
    .Y(_183_));
 sky130_fd_sc_hd__inv_2 _230_ (.A(\mem_top_ipin_7.DFFR_4_.Q ),
    .Y(_181_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(\mem_top_ipin_7.DFFR_0_.Q ),
    .Y(_191_));
 sky130_fd_sc_hd__inv_2 _232_ (.A(\mem_top_ipin_7.DFFR_2_.Q ),
    .Y(_186_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(\mem_top_ipin_7.DFFR_1_.Q ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_2 _234_ (.A(\mem_top_ipin_6.DFFR_3_.Q ),
    .Y(_177_));
 sky130_fd_sc_hd__inv_2 _235_ (.A(\mem_top_ipin_6.DFFR_0_.Q ),
    .Y(_180_));
 sky130_fd_sc_hd__inv_2 _236_ (.A(\mem_top_ipin_6.DFFR_2_.Q ),
    .Y(_176_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(\mem_top_ipin_6.DFFR_1_.Q ),
    .Y(_175_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(\mem_top_ipin_6.DFFR_5_.Q ),
    .Y(_170_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\mem_top_ipin_6.DFFR_0_.Q ),
    .Y(_178_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(\mem_top_ipin_6.DFFR_2_.Q ),
    .Y(_172_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(\mem_top_ipin_6.DFFR_1_.Q ),
    .Y(_171_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(\mem_top_ipin_6.DFFR_4_.Q ),
    .Y(_169_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(\mem_top_ipin_6.DFFR_0_.Q ),
    .Y(_179_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(\mem_top_ipin_6.DFFR_2_.Q ),
    .Y(_174_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(\mem_top_ipin_6.DFFR_1_.Q ),
    .Y(_173_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(\mem_top_ipin_5.DFFR_3_.Q ),
    .Y(_165_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(\mem_top_ipin_5.DFFR_0_.Q ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(\mem_top_ipin_5.DFFR_2_.Q ),
    .Y(_164_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(\mem_top_ipin_5.DFFR_1_.Q ),
    .Y(_163_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(\mem_top_ipin_5.DFFR_5_.Q ),
    .Y(_158_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(\mem_top_ipin_5.DFFR_0_.Q ),
    .Y(_166_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(\mem_top_ipin_5.DFFR_2_.Q ),
    .Y(_160_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(\mem_top_ipin_5.DFFR_1_.Q ),
    .Y(_159_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(\mem_top_ipin_5.DFFR_4_.Q ),
    .Y(_157_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(\mem_top_ipin_5.DFFR_0_.Q ),
    .Y(_167_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(\mem_top_ipin_5.DFFR_2_.Q ),
    .Y(_162_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(\mem_top_ipin_5.DFFR_1_.Q ),
    .Y(_161_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(\mem_top_ipin_4.DFFR_3_.Q ),
    .Y(_153_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(\mem_top_ipin_4.DFFR_0_.Q ),
    .Y(_156_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(\mem_top_ipin_4.DFFR_2_.Q ),
    .Y(_152_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(\mem_top_ipin_4.DFFR_1_.Q ),
    .Y(_151_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(\mem_top_ipin_4.DFFR_5_.Q ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(\mem_top_ipin_4.DFFR_0_.Q ),
    .Y(_154_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(\mem_top_ipin_4.DFFR_2_.Q ),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(\mem_top_ipin_4.DFFR_1_.Q ),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(\mem_top_ipin_4.DFFR_4_.Q ),
    .Y(_145_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(\mem_top_ipin_4.DFFR_0_.Q ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(\mem_top_ipin_4.DFFR_2_.Q ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(\mem_top_ipin_4.DFFR_1_.Q ),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _270_ (.A(\mem_top_ipin_3.DFFR_3_.Q ),
    .Y(_141_));
 sky130_fd_sc_hd__inv_2 _271_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_144_));
 sky130_fd_sc_hd__inv_2 _272_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_140_));
 sky130_fd_sc_hd__inv_2 _273_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _274_ (.A(\mem_top_ipin_3.DFFR_5_.Q ),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _275_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_142_));
 sky130_fd_sc_hd__inv_2 _276_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _277_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _278_ (.A(\mem_top_ipin_3.DFFR_4_.Q ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_143_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_138_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(\mem_top_ipin_2.DFFR_3_.Q ),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_128_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_127_));
 sky130_fd_sc_hd__inv_2 _286_ (.A(\mem_top_ipin_2.DFFR_5_.Q ),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _289_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _290_ (.A(\mem_top_ipin_2.DFFR_4_.Q ),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _292_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(\mem_top_ipin_1.DFFR_3_.Q ),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _297_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(\mem_top_ipin_1.DFFR_5_.Q ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _302_ (.A(\mem_top_ipin_1.DFFR_4_.Q ),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _303_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _305_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _306_ (.A(\mem_top_ipin_0.DFFR_3_.Q ),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _307_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _308_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _309_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(\mem_top_ipin_0.DFFR_5_.Q ),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _311_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _312_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _313_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _314_ (.A(\mem_top_ipin_0.DFFR_4_.Q ),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _316_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _318_ (.A(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _319_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _320_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _321_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _322_ (.A(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _323_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _324_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _325_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _327_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _329_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _331_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _332_ (.A(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _334_ (.A(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _335_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _341_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _342_ (.A(net24),
    .Y(\mux_bottom_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _343_ (.A(net11),
    .Y(\mux_bottom_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _344_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _345_ (.A(net30),
    .Y(\mux_bottom_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _346_ (.A(net2),
    .Y(\mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _347_ (.A(net21),
    .Y(\mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _348_ (.A(net17),
    .Y(\mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _349_ (.A(net36),
    .Y(\mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _350_ (.A(net5),
    .Y(\mux_bottom_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _351_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _352_ (.A(net6),
    .Y(\mux_bottom_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _353_ (.A(net37),
    .Y(\mux_bottom_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _354_ (.A(net18),
    .Y(\mux_bottom_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _355_ (.A(net31),
    .Y(\mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _356_ (.A(net12),
    .Y(\mux_bottom_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _357_ (.A(net25),
    .Y(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _359_ (.A(net8),
    .Y(\mux_top_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _360_ (.A(net39),
    .Y(\mux_top_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _361_ (.A(net20),
    .Y(\mux_top_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _362_ (.A(net33),
    .Y(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _363_ (.A(net14),
    .Y(\mux_top_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _364_ (.A(net27),
    .Y(\mux_top_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _366_ (.A(net9),
    .Y(\mux_top_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _367_ (.A(net22),
    .Y(\mux_top_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _368_ (.A(net3),
    .Y(\mux_top_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _369_ (.A(net34),
    .Y(\mux_top_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _370_ (.A(net15),
    .Y(\mux_top_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net28),
    .Y(\mux_top_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _372_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net43));
 sky130_fd_sc_hd__clkinv_2 _373_ (.A(net10),
    .Y(\mux_top_ipin_2.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _374_ (.A(net35),
    .Y(\mux_top_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _375_ (.A(net16),
    .Y(\mux_top_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _376_ (.A(net29),
    .Y(\mux_top_ipin_2.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _377_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _378_ (.A(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net45));
 sky130_fd_sc_hd__inv_2 _379_ (.A(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net46));
 sky130_fd_sc_hd__clkinv_2 _380_ (.A(net7),
    .Y(\mux_top_ipin_5.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _381_ (.A(net38),
    .Y(\mux_top_ipin_5.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _382_ (.A(net19),
    .Y(\mux_top_ipin_5.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _383_ (.A(net26),
    .Y(\mux_top_ipin_5.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _384_ (.A(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net47));
 sky130_fd_sc_hd__inv_2 _385_ (.A(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net48));
 sky130_fd_sc_hd__inv_2 _386_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _387_ (.A(net4),
    .Y(\mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net32),
    .Y(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net13),
    .Y(\mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net23),
    .Y(\mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_4 _391_ (.A(net40),
    .X(_066_));
 sky130_fd_sc_hd__buf_4 _392_ (.A(_066_),
    .X(_067_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(_067_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(_067_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(_067_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(_067_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(_067_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(_067_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(_067_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(_067_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(_067_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(_067_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_4 _403_ (.A(_066_),
    .X(_068_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(_068_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(_068_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _406_ (.A(_068_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(_068_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(_068_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(_068_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _410_ (.A(_068_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(_068_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _412_ (.A(_068_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _413_ (.A(_068_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _414_ (.A(_066_),
    .X(_069_));
 sky130_fd_sc_hd__inv_2 _415_ (.A(_069_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _416_ (.A(_069_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _417_ (.A(_069_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _418_ (.A(_069_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _419_ (.A(_069_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(_069_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _421_ (.A(_069_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _422_ (.A(_069_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _423_ (.A(_069_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _424_ (.A(_069_),
    .Y(_029_));
 sky130_fd_sc_hd__buf_4 _425_ (.A(_066_),
    .X(_070_));
 sky130_fd_sc_hd__inv_2 _426_ (.A(_070_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _427_ (.A(_070_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _428_ (.A(_070_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(_070_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_070_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(_070_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(_070_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(_070_),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _434_ (.A(_070_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(_070_),
    .Y(_039_));
 sky130_fd_sc_hd__buf_4 _436_ (.A(net40),
    .X(_071_));
 sky130_fd_sc_hd__inv_2 _437_ (.A(_071_),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _438_ (.A(_071_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _439_ (.A(_071_),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _440_ (.A(_071_),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _441_ (.A(_071_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _442_ (.A(_071_),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _443_ (.A(_071_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _444_ (.A(_071_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(_071_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _446_ (.A(_071_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_4 _447_ (.A(net40),
    .X(_072_));
 sky130_fd_sc_hd__inv_2 _448_ (.A(_072_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(_072_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(_072_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(_072_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(_072_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(_072_),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _454_ (.A(_072_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(_072_),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(_072_),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(_072_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _458_ (.A(_066_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _459_ (.A(_066_),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(_066_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _461_ (.A(_066_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _462_ (.A(_066_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _463_ (.A(_066_),
    .Y(_065_));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .RESET_B(_000_),
    .Q(\mem_bottom_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .RESET_B(_001_),
    .Q(\mem_bottom_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .RESET_B(_002_),
    .Q(\mem_bottom_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _467_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .RESET_B(_003_),
    .Q(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _468_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .RESET_B(_004_),
    .Q(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _469_ (.CLK(prog_clk),
    .D(net1),
    .RESET_B(_005_),
    .Q(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _470_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .RESET_B(_006_),
    .Q(\mem_bottom_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _471_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .RESET_B(_007_),
    .Q(\mem_bottom_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _472_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .RESET_B(_008_),
    .Q(\mem_bottom_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _473_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .RESET_B(_009_),
    .Q(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _474_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .RESET_B(_010_),
    .Q(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _475_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .RESET_B(_011_),
    .Q(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_4_.Q ),
    .RESET_B(_012_),
    .Q(\mem_top_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_3_.Q ),
    .RESET_B(_013_),
    .Q(\mem_top_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_2_.Q ),
    .RESET_B(_014_),
    .Q(\mem_top_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _479_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_1_.Q ),
    .RESET_B(_015_),
    .Q(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _480_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_0_.Q ),
    .RESET_B(_016_),
    .Q(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _481_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .RESET_B(_017_),
    .Q(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _482_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_4_.Q ),
    .RESET_B(_018_),
    .Q(\mem_top_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _483_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_3_.Q ),
    .RESET_B(_019_),
    .Q(\mem_top_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _484_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_2_.Q ),
    .RESET_B(_020_),
    .Q(\mem_top_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _485_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_1_.Q ),
    .RESET_B(_021_),
    .Q(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _486_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_0_.Q ),
    .RESET_B(_022_),
    .Q(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _487_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_5_.Q ),
    .RESET_B(_023_),
    .Q(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _488_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_4_.Q ),
    .RESET_B(_024_),
    .Q(\mem_top_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _489_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_3_.Q ),
    .RESET_B(_025_),
    .Q(\mem_top_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _490_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_2_.Q ),
    .RESET_B(_026_),
    .Q(\mem_top_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _491_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_1_.Q ),
    .RESET_B(_027_),
    .Q(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _492_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_0_.Q ),
    .RESET_B(_028_),
    .Q(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _493_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_5_.Q ),
    .RESET_B(_029_),
    .Q(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_4_.Q ),
    .RESET_B(_030_),
    .Q(\mem_top_ipin_3.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_3_.Q ),
    .RESET_B(_031_),
    .Q(\mem_top_ipin_3.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_2_.Q ),
    .RESET_B(_032_),
    .Q(\mem_top_ipin_3.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _497_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_1_.Q ),
    .RESET_B(_033_),
    .Q(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _498_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_0_.Q ),
    .RESET_B(_034_),
    .Q(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _499_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_5_.Q ),
    .RESET_B(_035_),
    .Q(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_4_.Q ),
    .RESET_B(_036_),
    .Q(\mem_top_ipin_4.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_3_.Q ),
    .RESET_B(_037_),
    .Q(\mem_top_ipin_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_2_.Q ),
    .RESET_B(_038_),
    .Q(\mem_top_ipin_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _503_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_1_.Q ),
    .RESET_B(_039_),
    .Q(\mem_top_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _504_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_0_.Q ),
    .RESET_B(_040_),
    .Q(\mem_top_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _505_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_5_.Q ),
    .RESET_B(_041_),
    .Q(\mem_top_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_4_.Q ),
    .RESET_B(_042_),
    .Q(\mem_top_ipin_5.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _507_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_3_.Q ),
    .RESET_B(_043_),
    .Q(\mem_top_ipin_5.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_2_.Q ),
    .RESET_B(_044_),
    .Q(\mem_top_ipin_5.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _509_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_1_.Q ),
    .RESET_B(_045_),
    .Q(\mem_top_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _510_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_0_.Q ),
    .RESET_B(_046_),
    .Q(\mem_top_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _511_ (.CLK(prog_clk),
    .D(\mem_top_ipin_4.DFFR_5_.Q ),
    .RESET_B(_047_),
    .Q(\mem_top_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_4_.Q ),
    .RESET_B(_048_),
    .Q(\mem_top_ipin_6.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _513_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_3_.Q ),
    .RESET_B(_049_),
    .Q(\mem_top_ipin_6.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_2_.Q ),
    .RESET_B(_050_),
    .Q(\mem_top_ipin_6.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _515_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_1_.Q ),
    .RESET_B(_051_),
    .Q(\mem_top_ipin_6.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _516_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_0_.Q ),
    .RESET_B(_052_),
    .Q(\mem_top_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _517_ (.CLK(prog_clk),
    .D(\mem_top_ipin_5.DFFR_5_.Q ),
    .RESET_B(_053_),
    .Q(\mem_top_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _518_ (.CLK(prog_clk),
    .D(\mem_top_ipin_7.DFFR_4_.Q ),
    .RESET_B(_054_),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _519_ (.CLK(prog_clk),
    .D(\mem_top_ipin_7.DFFR_3_.Q ),
    .RESET_B(_055_),
    .Q(\mem_top_ipin_7.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(prog_clk),
    .D(\mem_top_ipin_7.DFFR_2_.Q ),
    .RESET_B(_056_),
    .Q(\mem_top_ipin_7.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _521_ (.CLK(prog_clk),
    .D(\mem_top_ipin_7.DFFR_1_.Q ),
    .RESET_B(_057_),
    .Q(\mem_top_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _522_ (.CLK(prog_clk),
    .D(\mem_top_ipin_7.DFFR_0_.Q ),
    .RESET_B(_058_),
    .Q(\mem_top_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _523_ (.CLK(prog_clk),
    .D(\mem_top_ipin_6.DFFR_5_.Q ),
    .RESET_B(_059_),
    .Q(\mem_top_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .RESET_B(_060_),
    .Q(\mem_bottom_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _525_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .RESET_B(_061_),
    .Q(\mem_bottom_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .RESET_B(_062_),
    .Q(\mem_bottom_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _527_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .RESET_B(_063_),
    .Q(\mem_bottom_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _528_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .RESET_B(_064_),
    .Q(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _529_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .RESET_B(_065_),
    .Q(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _592__92 (.HI(net92));
 sky130_fd_sc_hd__conb_1 _606__93 (.HI(net93));
 sky130_fd_sc_hd__conb_1 _618__94 (.HI(net94));
 sky130_fd_sc_hd__conb_1 _630__95 (.HI(net95));
 sky130_fd_sc_hd__conb_1 _642__96 (.HI(net96));
 sky130_fd_sc_hd__conb_1 _654__97 (.HI(net97));
 sky130_fd_sc_hd__conb_1 _666__98 (.HI(net98));
 sky130_fd_sc_hd__conb_1 _678__99 (.HI(net99));
 sky130_fd_sc_hd__conb_1 _690__100 (.HI(net100));
 sky130_fd_sc_hd__conb_1 _700__101 (.HI(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__520__RESET_B (.DIODE(_056_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(net4),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _542_ (.A(net3),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 _543_ (.A(net20),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 _544_ (.A(net19),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _545_ (.A(net18),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _546_ (.A(net17),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _547_ (.A(net16),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _548_ (.A(net15),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _549_ (.A(net14),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 _550_ (.A(net13),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 _551_ (.A(net12),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(net2),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 _553_ (.A(net30),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(net29),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 _555_ (.A(net28),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 _556_ (.A(net27),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _557_ (.A(net26),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _558_ (.A(net25),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _559_ (.A(net24),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _560_ (.A(net23),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _561_ (.A(net22),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _562_ (.A(net39),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _563_ (.A(net38),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _564_ (.A(net37),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _565_ (.A(net36),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 _566_ (.A(net35),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(net34),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _568_ (.A(net33),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(net32),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _570_ (.A(net31),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(net21),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _572_ (.A(net11),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(net10),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _574_ (.A(net9),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _575_ (.A(net8),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 _576_ (.A(net7),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _577_ (.A(net6),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _578_ (.A(net5),
    .X(net72));
 sky130_fd_sc_hd__ebufn_2 _579_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_073_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _580_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_074_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _581_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_075_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _582_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_076_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _583_ (.A(net91),
    .TE_B(_077_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _584_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_078_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _585_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_079_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _586_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_080_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _587_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_081_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _588_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_082_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _589_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_083_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _590_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_084_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _591_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_085_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _592_ (.A(net92),
    .TE_B(_086_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _593_ (.A(\mux_bottom_ipin_1.INVTX1_7_.out ),
    .TE_B(_087_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _594_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_088_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _595_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_089_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _596_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_090_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _597_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_091_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _598_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_092_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _599_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_093_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _600_ (.A(\mux_bottom_ipin_1.INVTX1_6_.out ),
    .TE_B(_094_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _601_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_095_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _602_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_096_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _603_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_097_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _604_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_098_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _605_ (.A(\mux_top_ipin_0.INVTX1_7_.out ),
    .TE_B(_099_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _606_ (.A(net93),
    .TE_B(_100_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _607_ (.A(\mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_101_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _608_ (.A(\mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_102_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _609_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_103_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _610_ (.A(\mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_104_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _611_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_105_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _612_ (.A(\mux_top_ipin_0.INVTX1_6_.out ),
    .TE_B(_106_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _613_ (.A(\mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_107_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _614_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_108_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _615_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_109_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _616_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_110_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _617_ (.A(\mux_top_ipin_1.INVTX1_7_.out ),
    .TE_B(_111_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _618_ (.A(net94),
    .TE_B(_112_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _619_ (.A(\mux_top_ipin_1.INVTX1_4_.out ),
    .TE_B(_113_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _620_ (.A(\mux_top_ipin_1.INVTX1_5_.out ),
    .TE_B(_114_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _621_ (.A(\mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_115_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _622_ (.A(\mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_116_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _623_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_117_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _624_ (.A(\mux_top_ipin_1.INVTX1_6_.out ),
    .TE_B(_118_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _625_ (.A(\mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_119_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _626_ (.A(\mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_120_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _627_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_121_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _628_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_122_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _629_ (.A(\mux_top_ipin_2.INVTX1_7_.out ),
    .TE_B(_123_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _630_ (.A(net95),
    .TE_B(_124_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _631_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_125_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _632_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_126_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _633_ (.A(\mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_127_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _634_ (.A(\mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_128_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _635_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_129_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _636_ (.A(\mux_top_ipin_2.INVTX1_6_.out ),
    .TE_B(_130_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _637_ (.A(\mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_131_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _638_ (.A(\mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_132_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _639_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_133_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _640_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_134_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _641_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_135_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _642_ (.A(net96),
    .TE_B(_136_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _643_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_137_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _644_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_138_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _645_ (.A(\mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_139_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _646_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_140_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _647_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_141_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _648_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_142_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _649_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_143_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _650_ (.A(\mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_144_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _651_ (.A(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_145_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _652_ (.A(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_146_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _653_ (.A(\mux_bottom_ipin_1.INVTX1_7_.out ),
    .TE_B(_147_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _654_ (.A(net97),
    .TE_B(_148_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _655_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_149_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _656_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_150_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _657_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_151_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _658_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_152_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _659_ (.A(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_153_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _660_ (.A(\mux_bottom_ipin_1.INVTX1_6_.out ),
    .TE_B(_154_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _661_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_155_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _662_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_156_),
    .Z(\mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _663_ (.A(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_157_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _664_ (.A(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_158_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _665_ (.A(\mux_top_ipin_5.INVTX1_7_.out ),
    .TE_B(_159_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _666_ (.A(net98),
    .TE_B(_160_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _667_ (.A(\mux_top_ipin_5.INVTX1_4_.out ),
    .TE_B(_161_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _668_ (.A(\mux_top_ipin_5.INVTX1_5_.out ),
    .TE_B(_162_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _669_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_163_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _670_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_164_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _671_ (.A(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_165_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _672_ (.A(\mux_top_ipin_5.INVTX1_6_.out ),
    .TE_B(_166_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _673_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_167_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _674_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_168_),
    .Z(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _675_ (.A(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_169_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _676_ (.A(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_170_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _677_ (.A(\mux_top_ipin_0.INVTX1_7_.out ),
    .TE_B(_171_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _678_ (.A(net99),
    .TE_B(_172_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _679_ (.A(\mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_173_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _680_ (.A(\mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_174_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _681_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_175_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _682_ (.A(\mux_top_ipin_5.INVTX1_4_.out ),
    .TE_B(_176_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _683_ (.A(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_177_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _684_ (.A(\mux_top_ipin_0.INVTX1_6_.out ),
    .TE_B(_178_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _685_ (.A(\mux_top_ipin_5.INVTX1_5_.out ),
    .TE_B(_179_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _686_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_180_),
    .Z(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _687_ (.A(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_181_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _688_ (.A(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_182_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _689_ (.A(\mux_top_ipin_1.INVTX1_7_.out ),
    .TE_B(_183_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _690_ (.A(net100),
    .TE_B(_184_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _691_ (.A(\mux_top_ipin_1.INVTX1_4_.out ),
    .TE_B(_185_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _692_ (.A(\mux_top_ipin_1.INVTX1_5_.out ),
    .TE_B(_186_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _693_ (.A(\mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_187_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _694_ (.A(\mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_188_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _695_ (.A(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_189_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _696_ (.A(\mux_top_ipin_1.INVTX1_6_.out ),
    .TE_B(_190_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _697_ (.A(\mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_191_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _698_ (.A(\mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_192_),
    .Z(\mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _699_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_193_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _700_ (.A(net101),
    .TE_B(_194_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _701_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_195_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _702_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_196_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _703_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_197_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _704_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_198_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _705_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_199_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _706_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_200_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _707_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_201_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ccff_head),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(chanx_left_in[0]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(chanx_left_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(chanx_left_in[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(chanx_left_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(chanx_left_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(chanx_left_in[14]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(chanx_left_in[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(chanx_left_in[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(chanx_left_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(chanx_left_in[18]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(chanx_left_in[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(chanx_left_in[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(chanx_left_in[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(chanx_left_in[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(chanx_left_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chanx_left_in[6]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(chanx_left_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(chanx_left_in[8]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(chanx_left_in[9]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(chanx_right_in[0]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(chanx_right_in[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(chanx_right_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chanx_right_in[12]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(chanx_right_in[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(chanx_right_in[14]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(chanx_right_in[15]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(chanx_right_in[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(chanx_right_in[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(chanx_right_in[18]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(chanx_right_in[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chanx_right_in[2]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(chanx_right_in[3]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(chanx_right_in[4]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(chanx_right_in[5]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(chanx_right_in[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(chanx_right_in[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(chanx_right_in[8]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(chanx_right_in[9]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(pReset),
    .X(net40));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_));
 sky130_fd_sc_hd__conb_1 _583__91 (.HI(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__525__RESET_B (.DIODE(_061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__402__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__401__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__400__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__399__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__398__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__397__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__396__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__395__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__393__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__413__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__412__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__411__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__410__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__409__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__408__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__404__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__424__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__423__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__422__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__421__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__420__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__419__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__418__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__417__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__416__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__415__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__435__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__434__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__432__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__430__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__429__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__428__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__427__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__426__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__446__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__445__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__443__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__442__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__441__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__440__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__439__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__438__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__437__A (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__640__TE_B (.DIODE(_134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(chanx_left_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(chanx_left_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(chanx_left_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(chanx_left_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(chanx_left_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(chanx_left_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(chanx_left_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(chanx_left_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(chanx_left_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(chanx_left_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chanx_left_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chanx_left_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chanx_left_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chanx_left_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chanx_left_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chanx_left_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chanx_left_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chanx_left_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chanx_left_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chanx_right_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chanx_right_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chanx_right_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chanx_right_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chanx_right_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chanx_right_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chanx_right_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chanx_right_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chanx_right_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chanx_right_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chanx_right_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chanx_right_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chanx_right_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chanx_right_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chanx_right_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chanx_right_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chanx_right_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chanx_right_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chanx_right_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__468__D (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__335__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__333__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__331__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__D (.DIODE(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__340__A (.DIODE(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__A (.DIODE(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__336__A (.DIODE(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__D (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__341__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__339__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__337__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__D (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__327__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__323__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__319__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__473__D (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__328__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__324__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__320__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__472__D (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__329__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__325__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__321__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__525__D (.DIODE(\mem_bottom_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A (.DIODE(\mem_bottom_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__D (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__315__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__307__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__479__D (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__317__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__313__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__309__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__D (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__316__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__308__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__D (.DIODE(\mem_top_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__314__A (.DIODE(\mem_top_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__485__D (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__305__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__301__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__297__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__D (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__304__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__D (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__491__D (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__293__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__D (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__292__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__D (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__D (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__D (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__D (.DIODE(\mem_top_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A (.DIODE(\mem_top_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A (.DIODE(\mem_top_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__A (.DIODE(\mem_top_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__501__D (.DIODE(\mem_top_ipin_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A (.DIODE(\mem_top_ipin_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__500__D (.DIODE(\mem_top_ipin_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A (.DIODE(\mem_top_ipin_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__D (.DIODE(\mem_top_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A (.DIODE(\mem_top_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A (.DIODE(\mem_top_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A (.DIODE(\mem_top_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__509__D (.DIODE(\mem_top_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__257__A (.DIODE(\mem_top_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A (.DIODE(\mem_top_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__A (.DIODE(\mem_top_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__D (.DIODE(\mem_top_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A (.DIODE(\mem_top_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A (.DIODE(\mem_top_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(\mem_top_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__516__D (.DIODE(\mem_top_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A (.DIODE(\mem_top_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A (.DIODE(\mem_top_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A (.DIODE(\mem_top_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__D (.DIODE(\mem_top_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A (.DIODE(\mem_top_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__A (.DIODE(\mem_top_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__A (.DIODE(\mem_top_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__522__D (.DIODE(\mem_top_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__A (.DIODE(\mem_top_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__A (.DIODE(\mem_top_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__A (.DIODE(\mem_top_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__520__D (.DIODE(\mem_top_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__232__A (.DIODE(\mem_top_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__228__A (.DIODE(\mem_top_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__224__A (.DIODE(\mem_top_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__344__A (.DIODE(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__653__A (.DIODE(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__593__A (.DIODE(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__693__A (.DIODE(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__621__A (.DIODE(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__613__A (.DIODE(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__615__A (.DIODE(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__365__A (.DIODE(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__372__A (.DIODE(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__377__A (.DIODE(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__671__A (.DIODE(\mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(\mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(pReset));
 sky130_fd_sc_hd__diode_2 ANTENNA__529__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__528__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__527__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__526__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__525__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__524__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__523__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__522__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__521__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__520__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__519__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__518__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__517__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__516__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__514__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__513__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__512__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__511__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__509__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__507__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__506__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__505__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__504__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__503__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__501__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__500__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__495__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__491__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__489__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__488__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__487__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__486__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__485__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__483__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__482__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__481__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__479__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__477__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__475__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__473__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__472__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__471__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__470__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__469__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__468__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__465__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__469__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__542__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__368__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__541__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__387__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__578__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__350__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__577__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__352__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__576__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__380__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__574__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__366__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__573__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__373__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__572__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__343__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__550__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__549__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__363__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__548__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__370__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__547__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__375__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__546__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__348__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__543__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__361__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__571__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__347__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__560__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__559__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__342__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__557__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__383__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__556__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__364__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__555__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__371__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__554__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__376__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__553__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__345__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__570__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__355__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__568__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__362__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__565__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__349__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__564__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__353__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__563__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__381__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__562__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__360__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_399 ();
endmodule

