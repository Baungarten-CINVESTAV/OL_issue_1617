magic
tech sky130A
magscale 1 2
timestamp 1674174962
<< viali >>
rect 19698 37417 19732 37451
rect 8401 37349 8435 37383
rect 10425 37349 10459 37383
rect 18429 37349 18463 37383
rect 18797 37349 18831 37383
rect 23397 37349 23431 37383
rect 1593 37281 1627 37315
rect 5181 37281 5215 37315
rect 6561 37281 6595 37315
rect 11805 37281 11839 37315
rect 12357 37281 12391 37315
rect 15485 37281 15519 37315
rect 22937 37281 22971 37315
rect 25145 37281 25179 37315
rect 29745 37281 29779 37315
rect 32689 37281 32723 37315
rect 35173 37281 35207 37315
rect 37473 37281 37507 37315
rect 1869 37213 1903 37247
rect 2881 37213 2915 37247
rect 3985 37213 4019 37247
rect 5457 37213 5491 37247
rect 6837 37213 6871 37247
rect 8585 37213 8619 37247
rect 9873 37213 9907 37247
rect 10333 37213 10367 37247
rect 11161 37213 11195 37247
rect 11713 37213 11747 37247
rect 12633 37213 12667 37247
rect 14749 37213 14783 37247
rect 15761 37213 15795 37247
rect 18245 37213 18279 37247
rect 19441 37213 19475 37247
rect 22201 37213 22235 37247
rect 22753 37213 22787 37247
rect 23581 37213 23615 37247
rect 24869 37213 24903 37247
rect 27169 37213 27203 37247
rect 28089 37213 28123 37247
rect 28733 37213 28767 37247
rect 30021 37213 30055 37247
rect 31217 37213 31251 37247
rect 32413 37213 32447 37247
rect 34989 37213 35023 37247
rect 36185 37213 36219 37247
rect 37749 37213 37783 37247
rect 16957 37145 16991 37179
rect 17049 37145 17083 37179
rect 17969 37145 18003 37179
rect 3065 37077 3099 37111
rect 4169 37077 4203 37111
rect 9689 37077 9723 37111
rect 10977 37077 11011 37111
rect 14933 37077 14967 37111
rect 21189 37077 21223 37111
rect 22017 37077 22051 37111
rect 26617 37077 26651 37111
rect 27353 37077 27387 37111
rect 27905 37077 27939 37111
rect 28549 37077 28583 37111
rect 31033 37077 31067 37111
rect 34161 37077 34195 37111
rect 36369 37077 36403 37111
rect 3801 36873 3835 36907
rect 5181 36873 5215 36907
rect 12357 36873 12391 36907
rect 13829 36873 13863 36907
rect 25881 36873 25915 36907
rect 32505 36873 32539 36907
rect 33241 36873 33275 36907
rect 37657 36873 37691 36907
rect 1685 36805 1719 36839
rect 1777 36805 1811 36839
rect 9137 36805 9171 36839
rect 15393 36805 15427 36839
rect 23581 36805 23615 36839
rect 30205 36805 30239 36839
rect 3341 36737 3375 36771
rect 3985 36737 4019 36771
rect 4721 36737 4755 36771
rect 5365 36737 5399 36771
rect 6009 36737 6043 36771
rect 7021 36737 7055 36771
rect 7849 36737 7883 36771
rect 8401 36737 8435 36771
rect 9045 36737 9079 36771
rect 10517 36737 10551 36771
rect 10977 36737 11011 36771
rect 11897 36737 11931 36771
rect 13001 36737 13035 36771
rect 13645 36737 13679 36771
rect 14381 36737 14415 36771
rect 16865 36737 16899 36771
rect 25789 36737 25823 36771
rect 26617 36737 26651 36771
rect 30113 36737 30147 36771
rect 31125 36737 31159 36771
rect 31585 36737 31619 36771
rect 32321 36737 32355 36771
rect 33057 36737 33091 36771
rect 33977 36737 34011 36771
rect 36737 36737 36771 36771
rect 37473 36737 37507 36771
rect 2697 36669 2731 36703
rect 9689 36669 9723 36703
rect 11713 36669 11747 36703
rect 15301 36669 15335 36703
rect 16313 36669 16347 36703
rect 17141 36669 17175 36703
rect 18153 36669 18187 36703
rect 18429 36669 18463 36703
rect 20361 36669 20395 36703
rect 20637 36669 20671 36703
rect 23305 36669 23339 36703
rect 25329 36669 25363 36703
rect 27629 36669 27663 36703
rect 27905 36669 27939 36703
rect 29653 36669 29687 36703
rect 34437 36669 34471 36703
rect 34713 36669 34747 36703
rect 4537 36601 4571 36635
rect 7113 36601 7147 36635
rect 8585 36601 8619 36635
rect 30941 36601 30975 36635
rect 3157 36533 3191 36567
rect 5825 36533 5859 36567
rect 7665 36533 7699 36567
rect 10333 36533 10367 36567
rect 11069 36533 11103 36567
rect 12817 36533 12851 36567
rect 14381 36533 14415 36567
rect 19901 36533 19935 36567
rect 26433 36533 26467 36567
rect 31677 36533 31711 36567
rect 33793 36533 33827 36567
rect 36185 36533 36219 36567
rect 36829 36533 36863 36567
rect 7113 36329 7147 36363
rect 8493 36329 8527 36363
rect 29009 36329 29043 36363
rect 7849 36261 7883 36295
rect 10149 36261 10183 36295
rect 14933 36261 14967 36295
rect 26341 36261 26375 36295
rect 37565 36261 37599 36295
rect 2697 36193 2731 36227
rect 10793 36193 10827 36227
rect 12817 36193 12851 36227
rect 13461 36193 13495 36227
rect 15577 36193 15611 36227
rect 16773 36193 16807 36227
rect 21741 36193 21775 36227
rect 26801 36193 26835 36227
rect 29745 36193 29779 36227
rect 32229 36193 32263 36227
rect 34897 36193 34931 36227
rect 1777 36125 1811 36159
rect 4169 36125 4203 36159
rect 6009 36125 6043 36159
rect 6469 36125 6503 36159
rect 7297 36125 7331 36159
rect 7757 36125 7791 36159
rect 8401 36125 8435 36159
rect 9321 36125 9355 36159
rect 10057 36125 10091 36159
rect 13001 36125 13035 36159
rect 14841 36125 14875 36159
rect 18245 36125 18279 36159
rect 19441 36125 19475 36159
rect 24593 36125 24627 36159
rect 29193 36125 29227 36159
rect 37381 36125 37415 36159
rect 38025 36125 38059 36159
rect 2421 36057 2455 36091
rect 2513 36057 2547 36091
rect 9413 36057 9447 36091
rect 10885 36057 10919 36091
rect 11805 36057 11839 36091
rect 15669 36057 15703 36091
rect 16221 36057 16255 36091
rect 16865 36057 16899 36091
rect 17785 36057 17819 36091
rect 19717 36057 19751 36091
rect 22017 36057 22051 36091
rect 24869 36057 24903 36091
rect 27077 36057 27111 36091
rect 30021 36057 30055 36091
rect 31769 36057 31803 36091
rect 32505 36057 32539 36091
rect 35173 36057 35207 36091
rect 1593 35989 1627 36023
rect 3985 35989 4019 36023
rect 5825 35989 5859 36023
rect 6561 35989 6595 36023
rect 18337 35989 18371 36023
rect 21189 35989 21223 36023
rect 23489 35989 23523 36023
rect 28549 35989 28583 36023
rect 33977 35989 34011 36023
rect 36645 35989 36679 36023
rect 38209 35989 38243 36023
rect 3341 35785 3375 35819
rect 13093 35785 13127 35819
rect 35633 35785 35667 35819
rect 36829 35785 36863 35819
rect 1685 35717 1719 35751
rect 1777 35717 1811 35751
rect 2697 35717 2731 35751
rect 7849 35717 7883 35751
rect 10609 35717 10643 35751
rect 17049 35717 17083 35751
rect 17601 35717 17635 35751
rect 18429 35717 18463 35751
rect 28273 35717 28307 35751
rect 3249 35649 3283 35683
rect 9781 35649 9815 35683
rect 11805 35649 11839 35683
rect 12449 35649 12483 35683
rect 14105 35649 14139 35683
rect 14749 35649 14783 35683
rect 15393 35649 15427 35683
rect 16313 35649 16347 35683
rect 18153 35649 18187 35683
rect 27353 35649 27387 35683
rect 30297 35649 30331 35683
rect 30389 35649 30423 35683
rect 31217 35649 31251 35683
rect 32321 35649 32355 35683
rect 34897 35649 34931 35683
rect 35541 35649 35575 35683
rect 36737 35649 36771 35683
rect 38025 35649 38059 35683
rect 7021 35581 7055 35615
rect 7757 35581 7791 35615
rect 8769 35581 8803 35615
rect 10517 35581 10551 35615
rect 12633 35581 12667 35615
rect 14197 35581 14231 35615
rect 16957 35581 16991 35615
rect 24869 35581 24903 35615
rect 25145 35581 25179 35615
rect 27445 35581 27479 35615
rect 27997 35581 28031 35615
rect 9873 35513 9907 35547
rect 11069 35513 11103 35547
rect 31033 35513 31067 35547
rect 11897 35445 11931 35479
rect 14841 35445 14875 35479
rect 15485 35445 15519 35479
rect 16129 35445 16163 35479
rect 19901 35445 19935 35479
rect 26617 35445 26651 35479
rect 29745 35445 29779 35479
rect 32413 35445 32447 35479
rect 34989 35445 35023 35479
rect 38209 35445 38243 35479
rect 7665 35241 7699 35275
rect 10333 35241 10367 35275
rect 11069 35241 11103 35275
rect 13645 35241 13679 35275
rect 34989 35241 35023 35275
rect 36737 35241 36771 35275
rect 37381 35241 37415 35275
rect 38209 35241 38243 35275
rect 6561 35173 6595 35207
rect 11713 35173 11747 35207
rect 9137 35105 9171 35139
rect 9321 35105 9355 35139
rect 14565 35105 14599 35139
rect 24961 35105 24995 35139
rect 31493 35105 31527 35139
rect 31861 35105 31895 35139
rect 32597 35105 32631 35139
rect 1777 35037 1811 35071
rect 4353 35037 4387 35071
rect 6745 35037 6779 35071
rect 7573 35037 7607 35071
rect 8401 35037 8435 35071
rect 10241 35037 10275 35071
rect 10977 35037 11011 35071
rect 11621 35037 11655 35071
rect 12265 35037 12299 35071
rect 12909 35037 12943 35071
rect 13553 35037 13587 35071
rect 16405 35037 16439 35071
rect 27169 35037 27203 35071
rect 34897 35037 34931 35071
rect 36093 35037 36127 35071
rect 36921 35037 36955 35071
rect 37565 35037 37599 35071
rect 38025 35037 38059 35071
rect 12357 34969 12391 35003
rect 13001 34969 13035 35003
rect 14657 34969 14691 35003
rect 15577 34969 15611 35003
rect 16589 34969 16623 35003
rect 18245 34969 18279 35003
rect 21005 34969 21039 35003
rect 21833 34969 21867 35003
rect 25237 34969 25271 35003
rect 27905 34969 27939 35003
rect 29745 34969 29779 35003
rect 30573 34969 30607 35003
rect 31585 34969 31619 35003
rect 32873 34969 32907 35003
rect 1593 34901 1627 34935
rect 4169 34901 4203 34935
rect 8493 34901 8527 34935
rect 9781 34901 9815 34935
rect 26709 34901 26743 34935
rect 34345 34901 34379 34935
rect 36185 34901 36219 34935
rect 2421 34697 2455 34731
rect 21465 34697 21499 34731
rect 32965 34697 32999 34731
rect 35357 34697 35391 34731
rect 36829 34697 36863 34731
rect 11805 34629 11839 34663
rect 11897 34629 11931 34663
rect 13553 34629 13587 34663
rect 14105 34629 14139 34663
rect 15761 34629 15795 34663
rect 1593 34561 1627 34595
rect 2329 34561 2363 34595
rect 8309 34561 8343 34595
rect 8401 34561 8435 34595
rect 9597 34561 9631 34595
rect 10977 34561 11011 34595
rect 14565 34561 14599 34595
rect 14657 34561 14691 34595
rect 17233 34561 17267 34595
rect 24317 34561 24351 34595
rect 29285 34561 29319 34595
rect 32321 34561 32355 34595
rect 33609 34561 33643 34595
rect 34253 34561 34287 34595
rect 36277 34561 36311 34595
rect 36737 34561 36771 34595
rect 38025 34561 38059 34595
rect 9413 34493 9447 34527
rect 11069 34493 11103 34527
rect 13461 34493 13495 34527
rect 15669 34493 15703 34527
rect 19717 34493 19751 34527
rect 19993 34493 20027 34527
rect 22017 34493 22051 34527
rect 22293 34493 22327 34527
rect 23765 34493 23799 34527
rect 24593 34493 24627 34527
rect 26065 34493 26099 34527
rect 29561 34493 29595 34527
rect 31309 34493 31343 34527
rect 32505 34493 32539 34527
rect 34713 34493 34747 34527
rect 34897 34493 34931 34527
rect 9781 34425 9815 34459
rect 12357 34425 12391 34459
rect 16221 34425 16255 34459
rect 33425 34425 33459 34459
rect 34069 34425 34103 34459
rect 1777 34357 1811 34391
rect 17325 34357 17359 34391
rect 36093 34357 36127 34391
rect 38209 34357 38243 34391
rect 8493 34153 8527 34187
rect 11529 34153 11563 34187
rect 13553 34153 13587 34187
rect 16497 34153 16531 34187
rect 34253 34153 34287 34187
rect 10885 34085 10919 34119
rect 14657 34085 14691 34119
rect 24041 34085 24075 34119
rect 26617 34017 26651 34051
rect 26893 34017 26927 34051
rect 34989 34017 35023 34051
rect 35449 34017 35483 34051
rect 8401 33949 8435 33983
rect 9505 33949 9539 33983
rect 10149 33949 10183 33983
rect 10793 33949 10827 33983
rect 11437 33949 11471 33983
rect 13461 33949 13495 33983
rect 14565 33949 14599 33983
rect 16405 33949 16439 33983
rect 22293 33949 22327 33983
rect 32781 33949 32815 33983
rect 34161 33949 34195 33983
rect 36645 33949 36679 33983
rect 12173 33881 12207 33915
rect 12265 33881 12299 33915
rect 12817 33881 12851 33915
rect 15301 33881 15335 33915
rect 15393 33881 15427 33915
rect 15945 33881 15979 33915
rect 22569 33881 22603 33915
rect 31217 33881 31251 33915
rect 31309 33881 31343 33915
rect 31861 33881 31895 33915
rect 33517 33881 33551 33915
rect 35081 33881 35115 33915
rect 9597 33813 9631 33847
rect 10241 33813 10275 33847
rect 28365 33813 28399 33847
rect 36737 33813 36771 33847
rect 37565 33813 37599 33847
rect 6837 33609 6871 33643
rect 8585 33609 8619 33643
rect 15025 33609 15059 33643
rect 17141 33609 17175 33643
rect 31493 33609 31527 33643
rect 32413 33609 32447 33643
rect 35633 33609 35667 33643
rect 11897 33541 11931 33575
rect 13921 33541 13955 33575
rect 14473 33541 14507 33575
rect 15669 33541 15703 33575
rect 25145 33541 25179 33575
rect 6745 33473 6779 33507
rect 8493 33473 8527 33507
rect 9505 33473 9539 33507
rect 9597 33473 9631 33507
rect 10149 33473 10183 33507
rect 10977 33473 11011 33507
rect 13093 33473 13127 33507
rect 14933 33473 14967 33507
rect 15577 33473 15611 33507
rect 17049 33473 17083 33507
rect 31401 33473 31435 33507
rect 32321 33473 32355 33507
rect 32965 33473 32999 33507
rect 35541 33473 35575 33507
rect 36369 33473 36403 33507
rect 38117 33473 38151 33507
rect 11805 33405 11839 33439
rect 13829 33405 13863 33439
rect 18153 33405 18187 33439
rect 18429 33405 18463 33439
rect 24869 33405 24903 33439
rect 33241 33405 33275 33439
rect 12357 33337 12391 33371
rect 19901 33337 19935 33371
rect 38301 33337 38335 33371
rect 10241 33269 10275 33303
rect 11069 33269 11103 33303
rect 13185 33269 13219 33303
rect 26617 33269 26651 33303
rect 34713 33269 34747 33303
rect 36185 33269 36219 33303
rect 21189 33065 21223 33099
rect 34253 33065 34287 33099
rect 36645 33065 36679 33099
rect 37473 33065 37507 33099
rect 10609 32997 10643 33031
rect 12173 32929 12207 32963
rect 16037 32929 16071 32963
rect 17233 32929 17267 32963
rect 19441 32929 19475 32963
rect 24869 32929 24903 32963
rect 30757 32929 30791 32963
rect 34897 32929 34931 32963
rect 1593 32861 1627 32895
rect 7205 32861 7239 32895
rect 8585 32861 8619 32895
rect 9229 32861 9263 32895
rect 9873 32861 9907 32895
rect 10517 32861 10551 32895
rect 11161 32861 11195 32895
rect 13553 32861 13587 32895
rect 14381 32861 14415 32895
rect 15025 32861 15059 32895
rect 17141 32861 17175 32895
rect 24593 32861 24627 32895
rect 34161 32861 34195 32895
rect 37381 32861 37415 32895
rect 38025 32861 38059 32895
rect 9965 32793 9999 32827
rect 11897 32793 11931 32827
rect 11989 32793 12023 32827
rect 14473 32793 14507 32827
rect 16129 32793 16163 32827
rect 16681 32793 16715 32827
rect 19717 32793 19751 32827
rect 31033 32793 31067 32827
rect 35173 32793 35207 32827
rect 1777 32725 1811 32759
rect 7297 32725 7331 32759
rect 8401 32725 8435 32759
rect 9321 32725 9355 32759
rect 11253 32725 11287 32759
rect 13645 32725 13679 32759
rect 15117 32725 15151 32759
rect 26341 32725 26375 32759
rect 32505 32725 32539 32759
rect 38209 32725 38243 32759
rect 15025 32521 15059 32555
rect 22845 32521 22879 32555
rect 32781 32521 32815 32555
rect 9873 32453 9907 32487
rect 10793 32453 10827 32487
rect 11897 32453 11931 32487
rect 15761 32453 15795 32487
rect 24041 32453 24075 32487
rect 35173 32453 35207 32487
rect 1593 32385 1627 32419
rect 9229 32385 9263 32419
rect 12909 32385 12943 32419
rect 14013 32385 14047 32419
rect 14933 32385 14967 32419
rect 20361 32385 20395 32419
rect 22753 32385 22787 32419
rect 23765 32385 23799 32419
rect 27537 32385 27571 32419
rect 32689 32385 32723 32419
rect 34897 32385 34931 32419
rect 37657 32385 37691 32419
rect 9781 32317 9815 32351
rect 11805 32317 11839 32351
rect 14105 32317 14139 32351
rect 15669 32317 15703 32351
rect 15945 32317 15979 32351
rect 18337 32317 18371 32351
rect 18613 32317 18647 32351
rect 25789 32317 25823 32351
rect 36921 32317 36955 32351
rect 37473 32317 37507 32351
rect 9045 32249 9079 32283
rect 12357 32249 12391 32283
rect 1777 32181 1811 32215
rect 13001 32181 13035 32215
rect 27353 32181 27387 32215
rect 37841 32181 37875 32215
rect 9413 31977 9447 32011
rect 15117 31977 15151 32011
rect 17049 31977 17083 32011
rect 23581 31977 23615 32011
rect 6561 31909 6595 31943
rect 7757 31909 7791 31943
rect 13645 31909 13679 31943
rect 12081 31841 12115 31875
rect 12725 31841 12759 31875
rect 15761 31841 15795 31875
rect 21189 31841 21223 31875
rect 21833 31841 21867 31875
rect 24593 31841 24627 31875
rect 24869 31841 24903 31875
rect 26341 31841 26375 31875
rect 27629 31841 27663 31875
rect 36461 31841 36495 31875
rect 6745 31773 6779 31807
rect 7665 31773 7699 31807
rect 8493 31773 8527 31807
rect 9321 31773 9355 31807
rect 9965 31773 9999 31807
rect 10701 31773 10735 31807
rect 11345 31773 11379 31807
rect 13553 31773 13587 31807
rect 14289 31773 14323 31807
rect 14381 31773 14415 31807
rect 15025 31773 15059 31807
rect 16405 31773 16439 31807
rect 16957 31773 16991 31807
rect 19441 31773 19475 31807
rect 38301 31773 38335 31807
rect 11437 31705 11471 31739
rect 12173 31705 12207 31739
rect 15853 31705 15887 31739
rect 19717 31705 19751 31739
rect 22109 31705 22143 31739
rect 26893 31705 26927 31739
rect 36645 31705 36679 31739
rect 8309 31637 8343 31671
rect 10057 31637 10091 31671
rect 10793 31637 10827 31671
rect 9045 31433 9079 31467
rect 10425 31433 10459 31467
rect 15853 31433 15887 31467
rect 36829 31433 36863 31467
rect 9781 31365 9815 31399
rect 11805 31365 11839 31399
rect 14381 31365 14415 31399
rect 15301 31365 15335 31399
rect 20545 31365 20579 31399
rect 8401 31297 8435 31331
rect 9229 31297 9263 31331
rect 9689 31297 9723 31331
rect 10333 31297 10367 31331
rect 10977 31297 11011 31331
rect 11713 31297 11747 31331
rect 12909 31297 12943 31331
rect 13553 31297 13587 31331
rect 15761 31297 15795 31331
rect 18245 31297 18279 31331
rect 27261 31297 27295 31331
rect 36737 31297 36771 31331
rect 14289 31229 14323 31263
rect 18521 31229 18555 31263
rect 21373 31229 21407 31263
rect 23213 31229 23247 31263
rect 23489 31229 23523 31263
rect 25421 31229 25455 31263
rect 27537 31229 27571 31263
rect 29837 31229 29871 31263
rect 30113 31229 30147 31263
rect 32413 31229 32447 31263
rect 32689 31229 32723 31263
rect 37565 31229 37599 31263
rect 11069 31161 11103 31195
rect 13001 31161 13035 31195
rect 8493 31093 8527 31127
rect 13645 31093 13679 31127
rect 19993 31093 20027 31127
rect 24961 31093 24995 31127
rect 29009 31093 29043 31127
rect 31585 31093 31619 31127
rect 34161 31093 34195 31127
rect 16865 30889 16899 30923
rect 17404 30889 17438 30923
rect 18889 30889 18923 30923
rect 37841 30889 37875 30923
rect 7941 30753 7975 30787
rect 8125 30753 8159 30787
rect 9229 30753 9263 30787
rect 10793 30753 10827 30787
rect 11253 30753 11287 30787
rect 12633 30753 12667 30787
rect 17141 30753 17175 30787
rect 21005 30753 21039 30787
rect 24593 30753 24627 30787
rect 26433 30753 26467 30787
rect 29193 30753 29227 30787
rect 31033 30753 31067 30787
rect 35173 30753 35207 30787
rect 37473 30753 37507 30787
rect 1593 30685 1627 30719
rect 11897 30685 11931 30719
rect 27445 30685 27479 30719
rect 30757 30685 30791 30719
rect 34161 30685 34195 30719
rect 34897 30685 34931 30719
rect 37657 30685 37691 30719
rect 9321 30617 9355 30651
rect 10241 30617 10275 30651
rect 10885 30617 10919 30651
rect 12725 30617 12759 30651
rect 13277 30617 13311 30651
rect 15485 30617 15519 30651
rect 15577 30617 15611 30651
rect 16497 30617 16531 30651
rect 21281 30617 21315 30651
rect 23029 30617 23063 30651
rect 24777 30617 24811 30651
rect 27721 30617 27755 30651
rect 33425 30617 33459 30651
rect 1777 30549 1811 30583
rect 8585 30549 8619 30583
rect 11989 30549 12023 30583
rect 14289 30549 14323 30583
rect 32505 30549 32539 30583
rect 36645 30549 36679 30583
rect 38209 30345 38243 30379
rect 14197 30277 14231 30311
rect 14749 30277 14783 30311
rect 15301 30277 15335 30311
rect 15393 30277 15427 30311
rect 16957 30277 16991 30311
rect 30205 30277 30239 30311
rect 33425 30277 33459 30311
rect 36737 30277 36771 30311
rect 10333 30209 10367 30243
rect 10977 30209 11011 30243
rect 11805 30209 11839 30243
rect 12449 30209 12483 30243
rect 13185 30209 13219 30243
rect 16865 30209 16899 30243
rect 18245 30209 18279 30243
rect 24225 30209 24259 30243
rect 27169 30209 27203 30243
rect 33333 30209 33367 30243
rect 34713 30209 34747 30243
rect 38025 30209 38059 30243
rect 9689 30141 9723 30175
rect 14105 30141 14139 30175
rect 15577 30141 15611 30175
rect 18521 30141 18555 30175
rect 19993 30141 20027 30175
rect 26249 30141 26283 30175
rect 27445 30141 27479 30175
rect 29929 30141 29963 30175
rect 34989 30141 35023 30175
rect 10425 30073 10459 30107
rect 11897 30073 11931 30107
rect 11069 30005 11103 30039
rect 12541 30005 12575 30039
rect 13277 30005 13311 30039
rect 24482 30005 24516 30039
rect 28917 30005 28951 30039
rect 31677 30005 31711 30039
rect 8217 29801 8251 29835
rect 10609 29801 10643 29835
rect 14841 29801 14875 29835
rect 19698 29801 19732 29835
rect 1593 29733 1627 29767
rect 13645 29733 13679 29767
rect 16037 29733 16071 29767
rect 9965 29665 9999 29699
rect 11529 29665 11563 29699
rect 13093 29665 13127 29699
rect 21189 29665 21223 29699
rect 24593 29665 24627 29699
rect 30481 29665 30515 29699
rect 31401 29665 31435 29699
rect 34897 29665 34931 29699
rect 36645 29665 36679 29699
rect 1777 29597 1811 29631
rect 7573 29597 7607 29631
rect 7757 29597 7791 29631
rect 9505 29597 9539 29631
rect 10149 29597 10183 29631
rect 14749 29597 14783 29631
rect 19441 29597 19475 29631
rect 26985 29597 27019 29631
rect 29745 29597 29779 29631
rect 37289 29597 37323 29631
rect 38025 29597 38059 29631
rect 11161 29529 11195 29563
rect 11253 29529 11287 29563
rect 13185 29529 13219 29563
rect 15485 29529 15519 29563
rect 15577 29529 15611 29563
rect 24869 29529 24903 29563
rect 31677 29529 31711 29563
rect 35173 29529 35207 29563
rect 9321 29461 9355 29495
rect 26341 29461 26375 29495
rect 28273 29461 28307 29495
rect 33149 29461 33183 29495
rect 37105 29461 37139 29495
rect 38209 29461 38243 29495
rect 9781 29257 9815 29291
rect 13645 29257 13679 29291
rect 34253 29257 34287 29291
rect 11069 29189 11103 29223
rect 11897 29189 11931 29223
rect 14473 29189 14507 29223
rect 15662 29189 15696 29223
rect 20545 29189 20579 29223
rect 23305 29189 23339 29223
rect 25329 29189 25363 29223
rect 1593 29121 1627 29155
rect 9689 29121 9723 29155
rect 10333 29121 10367 29155
rect 10977 29121 11011 29155
rect 12909 29121 12943 29155
rect 13553 29121 13587 29155
rect 16865 29121 16899 29155
rect 32505 29121 32539 29155
rect 38025 29121 38059 29155
rect 10425 29053 10459 29087
rect 11805 29053 11839 29087
rect 12173 29053 12207 29087
rect 14381 29053 14415 29087
rect 14657 29053 14691 29087
rect 15577 29053 15611 29087
rect 16221 29053 16255 29087
rect 18245 29053 18279 29087
rect 21281 29053 21315 29087
rect 23029 29053 23063 29087
rect 24777 29053 24811 29087
rect 26065 29053 26099 29087
rect 1777 28985 1811 29019
rect 19993 28985 20027 29019
rect 38209 28985 38243 29019
rect 13001 28917 13035 28951
rect 16957 28917 16991 28951
rect 18508 28917 18542 28951
rect 32762 28917 32796 28951
rect 6653 28713 6687 28747
rect 10517 28713 10551 28747
rect 11713 28713 11747 28747
rect 13645 28713 13679 28747
rect 14381 28713 14415 28747
rect 15025 28713 15059 28747
rect 37473 28713 37507 28747
rect 7757 28577 7791 28611
rect 11253 28577 11287 28611
rect 16221 28577 16255 28611
rect 17417 28577 17451 28611
rect 20729 28577 20763 28611
rect 26341 28577 26375 28611
rect 31401 28577 31435 28611
rect 6837 28509 6871 28543
rect 7941 28509 7975 28543
rect 9137 28509 9171 28543
rect 10425 28509 10459 28543
rect 11069 28509 11103 28543
rect 12173 28509 12207 28543
rect 12817 28509 12851 28543
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 14933 28509 14967 28543
rect 16037 28509 16071 28543
rect 24593 28509 24627 28543
rect 28825 28509 28859 28543
rect 31125 28509 31159 28543
rect 34897 28509 34931 28543
rect 37657 28509 37691 28543
rect 38301 28509 38335 28543
rect 21005 28441 21039 28475
rect 22753 28441 22787 28475
rect 24869 28441 24903 28475
rect 28089 28441 28123 28475
rect 35173 28441 35207 28475
rect 8401 28373 8435 28407
rect 9229 28373 9263 28407
rect 12265 28373 12299 28407
rect 12909 28373 12943 28407
rect 32873 28373 32907 28407
rect 36645 28373 36679 28407
rect 38117 28373 38151 28407
rect 7573 28169 7607 28203
rect 8217 28169 8251 28203
rect 6929 28101 6963 28135
rect 10149 28101 10183 28135
rect 11069 28101 11103 28135
rect 11897 28101 11931 28135
rect 14197 28101 14231 28135
rect 15393 28101 15427 28135
rect 20269 28101 20303 28135
rect 33333 28101 33367 28135
rect 6837 28033 6871 28067
rect 7481 28033 7515 28067
rect 8125 28033 8159 28067
rect 10977 28033 11011 28067
rect 13369 28033 13403 28067
rect 22845 28033 22879 28067
rect 37749 28033 37783 28067
rect 11805 27965 11839 27999
rect 12449 27965 12483 27999
rect 14105 27965 14139 27999
rect 14565 27965 14599 27999
rect 15301 27965 15335 27999
rect 16221 27965 16255 27999
rect 18245 27965 18279 27999
rect 18521 27965 18555 27999
rect 23121 27965 23155 27999
rect 27629 27965 27663 27999
rect 27905 27965 27939 27999
rect 34069 27965 34103 27999
rect 10333 27897 10367 27931
rect 13461 27897 13495 27931
rect 24593 27829 24627 27863
rect 29377 27829 29411 27863
rect 37841 27829 37875 27863
rect 32210 27625 32244 27659
rect 35154 27625 35188 27659
rect 9689 27557 9723 27591
rect 13645 27557 13679 27591
rect 14289 27557 14323 27591
rect 26433 27557 26467 27591
rect 11897 27489 11931 27523
rect 27353 27489 27387 27523
rect 31493 27489 31527 27523
rect 31953 27489 31987 27523
rect 33701 27489 33735 27523
rect 34897 27489 34931 27523
rect 1777 27421 1811 27455
rect 9873 27421 9907 27455
rect 10333 27421 10367 27455
rect 13553 27421 13587 27455
rect 14473 27421 14507 27455
rect 15117 27421 15151 27455
rect 15209 27421 15243 27455
rect 24685 27421 24719 27455
rect 29745 27421 29779 27455
rect 38025 27421 38059 27455
rect 11989 27353 12023 27387
rect 12541 27353 12575 27387
rect 15853 27353 15887 27387
rect 15945 27353 15979 27387
rect 16865 27353 16899 27387
rect 24961 27353 24995 27387
rect 27629 27353 27663 27387
rect 30021 27353 30055 27387
rect 1593 27285 1627 27319
rect 10425 27285 10459 27319
rect 29101 27285 29135 27319
rect 36645 27285 36679 27319
rect 37657 27285 37691 27319
rect 38209 27285 38243 27319
rect 9229 27081 9263 27115
rect 13645 27081 13679 27115
rect 25145 27013 25179 27047
rect 9413 26945 9447 26979
rect 10977 26945 11011 26979
rect 11989 26945 12023 26979
rect 12633 26945 12667 26979
rect 13829 26945 13863 26979
rect 18153 26945 18187 26979
rect 22017 26945 22051 26979
rect 24869 26945 24903 26979
rect 27169 26945 27203 26979
rect 29469 26945 29503 26979
rect 32873 26945 32907 26979
rect 18429 26877 18463 26911
rect 20177 26877 20211 26911
rect 22293 26877 22327 26911
rect 24041 26877 24075 26911
rect 27445 26877 27479 26911
rect 29745 26877 29779 26911
rect 33149 26877 33183 26911
rect 11069 26809 11103 26843
rect 12081 26741 12115 26775
rect 12725 26741 12759 26775
rect 26617 26741 26651 26775
rect 28917 26741 28951 26775
rect 31217 26741 31251 26775
rect 34621 26741 34655 26775
rect 9781 26537 9815 26571
rect 13553 26537 13587 26571
rect 15577 26537 15611 26571
rect 21465 26537 21499 26571
rect 36645 26537 36679 26571
rect 1593 26469 1627 26503
rect 14381 26401 14415 26435
rect 14657 26401 14691 26435
rect 24593 26401 24627 26435
rect 24869 26401 24903 26435
rect 30849 26401 30883 26435
rect 32321 26401 32355 26435
rect 34897 26401 34931 26435
rect 37197 26401 37231 26435
rect 1777 26333 1811 26367
rect 8401 26333 8435 26367
rect 9137 26333 9171 26367
rect 9321 26333 9355 26367
rect 13737 26333 13771 26367
rect 15485 26333 15519 26367
rect 19717 26333 19751 26367
rect 22017 26333 22051 26367
rect 30573 26333 30607 26367
rect 10333 26265 10367 26299
rect 10425 26265 10459 26299
rect 11345 26265 11379 26299
rect 14473 26265 14507 26299
rect 19993 26265 20027 26299
rect 26617 26265 26651 26299
rect 35173 26265 35207 26299
rect 37289 26265 37323 26299
rect 38209 26265 38243 26299
rect 22109 26197 22143 26231
rect 8309 25993 8343 26027
rect 10609 25925 10643 25959
rect 12725 25925 12759 25959
rect 17417 25925 17451 25959
rect 32597 25925 32631 25959
rect 34989 25925 35023 25959
rect 5181 25857 5215 25891
rect 8493 25857 8527 25891
rect 11897 25857 11931 25891
rect 14933 25857 14967 25891
rect 22017 25857 22051 25891
rect 32321 25857 32355 25891
rect 38301 25857 38335 25891
rect 10517 25789 10551 25823
rect 12633 25789 12667 25823
rect 13277 25789 13311 25823
rect 17141 25789 17175 25823
rect 18889 25789 18923 25823
rect 19349 25789 19383 25823
rect 19625 25789 19659 25823
rect 22753 25789 22787 25823
rect 28733 25789 28767 25823
rect 29009 25789 29043 25823
rect 30757 25789 30791 25823
rect 34713 25789 34747 25823
rect 11069 25721 11103 25755
rect 34069 25721 34103 25755
rect 4997 25653 5031 25687
rect 11989 25653 12023 25687
rect 15025 25653 15059 25687
rect 21097 25653 21131 25687
rect 36461 25653 36495 25687
rect 38117 25653 38151 25687
rect 7757 25449 7791 25483
rect 9781 25449 9815 25483
rect 14381 25449 14415 25483
rect 16221 25449 16255 25483
rect 24041 25449 24075 25483
rect 37013 25449 37047 25483
rect 6929 25381 6963 25415
rect 37657 25381 37691 25415
rect 8493 25313 8527 25347
rect 9321 25313 9355 25347
rect 19441 25313 19475 25347
rect 22293 25313 22327 25347
rect 24593 25313 24627 25347
rect 7113 25245 7147 25279
rect 7941 25245 7975 25279
rect 8401 25245 8435 25279
rect 9137 25245 9171 25279
rect 14289 25245 14323 25279
rect 16129 25245 16163 25279
rect 33609 25245 33643 25279
rect 36921 25245 36955 25279
rect 38025 25245 38059 25279
rect 11621 25177 11655 25211
rect 11713 25177 11747 25211
rect 12265 25177 12299 25211
rect 15025 25177 15059 25211
rect 15117 25177 15151 25211
rect 15669 25177 15703 25211
rect 19717 25177 19751 25211
rect 21465 25177 21499 25211
rect 22569 25177 22603 25211
rect 24869 25177 24903 25211
rect 32873 25177 32907 25211
rect 26341 25109 26375 25143
rect 38209 25109 38243 25143
rect 24593 24905 24627 24939
rect 10517 24837 10551 24871
rect 12357 24837 12391 24871
rect 14657 24837 14691 24871
rect 23121 24837 23155 24871
rect 25053 24837 25087 24871
rect 1593 24769 1627 24803
rect 7849 24769 7883 24803
rect 8677 24769 8711 24803
rect 13829 24769 13863 24803
rect 13921 24769 13955 24803
rect 15669 24769 15703 24803
rect 15761 24769 15795 24803
rect 19165 24769 19199 24803
rect 32321 24769 32355 24803
rect 10425 24701 10459 24735
rect 12265 24701 12299 24735
rect 12817 24701 12851 24735
rect 14565 24701 14599 24735
rect 19441 24701 19475 24735
rect 22845 24701 22879 24735
rect 25789 24701 25823 24735
rect 27169 24701 27203 24735
rect 27445 24701 27479 24735
rect 29469 24701 29503 24735
rect 29745 24701 29779 24735
rect 32597 24701 32631 24735
rect 34069 24701 34103 24735
rect 10977 24633 11011 24667
rect 15117 24633 15151 24667
rect 1777 24565 1811 24599
rect 7941 24565 7975 24599
rect 8493 24565 8527 24599
rect 20913 24565 20947 24599
rect 28917 24565 28951 24599
rect 31217 24565 31251 24599
rect 9689 24361 9723 24395
rect 11161 24361 11195 24395
rect 11805 24361 11839 24395
rect 31953 24361 31987 24395
rect 34161 24361 34195 24395
rect 7849 24293 7883 24327
rect 14381 24293 14415 24327
rect 9321 24225 9355 24259
rect 12633 24225 12667 24259
rect 20085 24225 20119 24259
rect 24961 24225 24995 24259
rect 30481 24225 30515 24259
rect 32413 24225 32447 24259
rect 35173 24225 35207 24259
rect 1593 24157 1627 24191
rect 7297 24157 7331 24191
rect 7757 24157 7791 24191
rect 9137 24157 9171 24191
rect 11069 24157 11103 24191
rect 11713 24157 11747 24191
rect 12449 24157 12483 24191
rect 13369 24157 13403 24191
rect 14289 24157 14323 24191
rect 30205 24157 30239 24191
rect 34897 24157 34931 24191
rect 37473 24157 37507 24191
rect 37749 24157 37783 24191
rect 20361 24089 20395 24123
rect 24685 24089 24719 24123
rect 24777 24089 24811 24123
rect 32689 24089 32723 24123
rect 1777 24021 1811 24055
rect 7113 24021 7147 24055
rect 13461 24021 13495 24055
rect 21833 24021 21867 24055
rect 36645 24021 36679 24055
rect 29377 23817 29411 23851
rect 37565 23817 37599 23851
rect 11897 23749 11931 23783
rect 19533 23749 19567 23783
rect 21281 23749 21315 23783
rect 23673 23749 23707 23783
rect 13369 23681 13403 23715
rect 17049 23681 17083 23715
rect 19257 23681 19291 23715
rect 23397 23681 23431 23715
rect 27629 23681 27663 23715
rect 29837 23681 29871 23715
rect 34437 23681 34471 23715
rect 36461 23681 36495 23715
rect 37473 23681 37507 23715
rect 10977 23613 11011 23647
rect 11805 23613 11839 23647
rect 12265 23613 12299 23647
rect 17325 23613 17359 23647
rect 25421 23613 25455 23647
rect 27905 23613 27939 23647
rect 30113 23613 30147 23647
rect 34713 23613 34747 23647
rect 13461 23477 13495 23511
rect 18797 23477 18831 23511
rect 31585 23477 31619 23511
rect 9505 23273 9539 23307
rect 12449 23273 12483 23307
rect 15577 23273 15611 23307
rect 20729 23137 20763 23171
rect 23397 23137 23431 23171
rect 24041 23137 24075 23171
rect 30481 23137 30515 23171
rect 31493 23137 31527 23171
rect 33517 23137 33551 23171
rect 34897 23137 34931 23171
rect 9137 23069 9171 23103
rect 9321 23069 9355 23103
rect 11529 23069 11563 23103
rect 12357 23069 12391 23103
rect 15761 23069 15795 23103
rect 20453 23069 20487 23103
rect 25237 23069 25271 23103
rect 29745 23069 29779 23103
rect 37565 23069 37599 23103
rect 23489 23001 23523 23035
rect 25513 23001 25547 23035
rect 31769 23001 31803 23035
rect 35173 23001 35207 23035
rect 11621 22933 11655 22967
rect 22201 22933 22235 22967
rect 26985 22933 27019 22967
rect 36645 22933 36679 22967
rect 37657 22933 37691 22967
rect 31677 22729 31711 22763
rect 36553 22729 36587 22763
rect 12357 22661 12391 22695
rect 12449 22661 12483 22695
rect 14013 22661 14047 22695
rect 18797 22661 18831 22695
rect 23949 22661 23983 22695
rect 24501 22661 24535 22695
rect 25697 22661 25731 22695
rect 27445 22661 27479 22695
rect 1685 22593 1719 22627
rect 9137 22593 9171 22627
rect 10241 22593 10275 22627
rect 10977 22593 11011 22627
rect 15853 22593 15887 22627
rect 25421 22593 25455 22627
rect 26341 22593 26375 22627
rect 27169 22593 27203 22627
rect 29929 22593 29963 22627
rect 34345 22593 34379 22627
rect 34805 22593 34839 22627
rect 38025 22593 38059 22627
rect 8309 22525 8343 22559
rect 8953 22525 8987 22559
rect 13369 22525 13403 22559
rect 13921 22525 13955 22559
rect 14933 22525 14967 22559
rect 18521 22525 18555 22559
rect 23857 22525 23891 22559
rect 26433 22525 26467 22559
rect 30205 22525 30239 22559
rect 32321 22525 32355 22559
rect 32597 22525 32631 22559
rect 35081 22525 35115 22559
rect 1869 22457 1903 22491
rect 9321 22457 9355 22491
rect 10333 22457 10367 22491
rect 20269 22457 20303 22491
rect 28917 22457 28951 22491
rect 38209 22457 38243 22491
rect 11069 22389 11103 22423
rect 15945 22389 15979 22423
rect 29561 22389 29595 22423
rect 9229 22185 9263 22219
rect 15853 22185 15887 22219
rect 26144 22185 26178 22219
rect 37473 22185 37507 22219
rect 11621 22049 11655 22083
rect 12081 22049 12115 22083
rect 15393 22049 15427 22083
rect 24961 22049 24995 22083
rect 25881 22049 25915 22083
rect 28273 22049 28307 22083
rect 32597 22049 32631 22083
rect 34897 22049 34931 22083
rect 36645 22049 36679 22083
rect 1961 21981 1995 22015
rect 8217 21981 8251 22015
rect 9137 21981 9171 22015
rect 10885 21981 10919 22015
rect 16037 21981 16071 22015
rect 24869 21981 24903 22015
rect 28089 21981 28123 22015
rect 29009 21981 29043 22015
rect 37381 21983 37415 22017
rect 38301 21981 38335 22015
rect 11713 21913 11747 21947
rect 14381 21913 14415 21947
rect 14473 21913 14507 21947
rect 32873 21913 32907 21947
rect 35173 21913 35207 21947
rect 1777 21845 1811 21879
rect 8309 21845 8343 21879
rect 10977 21845 11011 21879
rect 27629 21845 27663 21879
rect 29101 21845 29135 21879
rect 34345 21845 34379 21879
rect 38117 21845 38151 21879
rect 14749 21641 14783 21675
rect 15393 21641 15427 21675
rect 23489 21641 23523 21675
rect 24501 21641 24535 21675
rect 25145 21641 25179 21675
rect 10149 21573 10183 21607
rect 26433 21573 26467 21607
rect 27997 21573 28031 21607
rect 28917 21573 28951 21607
rect 1593 21505 1627 21539
rect 8217 21505 8251 21539
rect 10701 21505 10735 21539
rect 14657 21505 14691 21539
rect 15301 21505 15335 21539
rect 23397 21505 23431 21539
rect 24409 21505 24443 21539
rect 25053 21505 25087 21539
rect 25697 21505 25731 21539
rect 26341 21505 26375 21539
rect 27629 21505 27663 21539
rect 34897 21505 34931 21539
rect 37657 21505 37691 21539
rect 10057 21437 10091 21471
rect 25789 21437 25823 21471
rect 28825 21437 28859 21471
rect 35173 21437 35207 21471
rect 38117 21437 38151 21471
rect 29377 21369 29411 21403
rect 1777 21301 1811 21335
rect 8309 21301 8343 21335
rect 36645 21301 36679 21335
rect 37473 21301 37507 21335
rect 1593 21097 1627 21131
rect 20637 21097 20671 21131
rect 22201 21097 22235 21131
rect 25881 21097 25915 21131
rect 26525 21097 26559 21131
rect 32229 21097 32263 21131
rect 33977 21097 34011 21131
rect 35909 21097 35943 21131
rect 23949 21029 23983 21063
rect 25237 21029 25271 21063
rect 17509 20961 17543 20995
rect 21373 20961 21407 20995
rect 28181 20961 28215 20995
rect 28457 20961 28491 20995
rect 30665 20961 30699 20995
rect 30941 20961 30975 20995
rect 36553 20961 36587 20995
rect 37289 20961 37323 20995
rect 37565 20961 37599 20995
rect 1777 20893 1811 20927
rect 16497 20893 16531 20927
rect 20545 20893 20579 20927
rect 21189 20893 21223 20927
rect 22109 20893 22143 20927
rect 25789 20893 25823 20927
rect 26433 20893 26467 20927
rect 27077 20893 27111 20927
rect 29745 20893 29779 20927
rect 32137 20893 32171 20927
rect 33241 20893 33275 20927
rect 33885 20893 33919 20927
rect 35173 20893 35207 20927
rect 35817 20893 35851 20927
rect 36461 20893 36495 20927
rect 17233 20825 17267 20859
rect 17325 20825 17359 20859
rect 23386 20825 23420 20859
rect 23482 20825 23516 20859
rect 24685 20825 24719 20859
rect 24777 20825 24811 20859
rect 27353 20825 27387 20859
rect 28273 20825 28307 20859
rect 30757 20825 30791 20859
rect 33333 20825 33367 20859
rect 37381 20825 37415 20859
rect 16589 20757 16623 20791
rect 29837 20757 29871 20791
rect 35265 20757 35299 20791
rect 6653 20553 6687 20587
rect 21281 20553 21315 20587
rect 23857 20553 23891 20587
rect 25053 20553 25087 20587
rect 28917 20553 28951 20587
rect 29561 20553 29595 20587
rect 33057 20553 33091 20587
rect 35541 20553 35575 20587
rect 36185 20553 36219 20587
rect 38209 20553 38243 20587
rect 16957 20485 16991 20519
rect 17049 20485 17083 20519
rect 26157 20485 26191 20519
rect 27445 20485 27479 20519
rect 30849 20485 30883 20519
rect 34069 20485 34103 20519
rect 6837 20417 6871 20451
rect 7481 20417 7515 20451
rect 18429 20417 18463 20451
rect 21189 20417 21223 20451
rect 22661 20417 22695 20451
rect 23765 20417 23799 20451
rect 24961 20417 24995 20451
rect 26065 20417 26099 20451
rect 28825 20417 28859 20451
rect 29469 20417 29503 20451
rect 32321 20417 32355 20451
rect 32965 20417 32999 20451
rect 35449 20417 35483 20451
rect 36093 20417 36127 20451
rect 36737 20417 36771 20451
rect 38025 20417 38059 20451
rect 14657 20349 14691 20383
rect 17877 20349 17911 20383
rect 23213 20349 23247 20383
rect 27353 20349 27387 20383
rect 27629 20349 27663 20383
rect 30757 20349 30791 20383
rect 31769 20349 31803 20383
rect 33977 20349 34011 20383
rect 34253 20349 34287 20383
rect 7297 20281 7331 20315
rect 18521 20213 18555 20247
rect 32413 20213 32447 20247
rect 36829 20213 36863 20247
rect 23029 20009 23063 20043
rect 23673 20009 23707 20043
rect 26157 20009 26191 20043
rect 28825 20009 28859 20043
rect 20085 19941 20119 19975
rect 14565 19873 14599 19907
rect 14841 19873 14875 19907
rect 24685 19873 24719 19907
rect 27445 19873 27479 19907
rect 28181 19873 28215 19907
rect 29745 19873 29779 19907
rect 29929 19873 29963 19907
rect 31585 19873 31619 19907
rect 33885 19873 33919 19907
rect 34989 19873 35023 19907
rect 35265 19873 35299 19907
rect 36461 19873 36495 19907
rect 38117 19873 38151 19907
rect 20637 19805 20671 19839
rect 21557 19805 21591 19839
rect 21649 19805 21683 19839
rect 22937 19805 22971 19839
rect 23581 19805 23615 19839
rect 24593 19805 24627 19839
rect 26065 19805 26099 19839
rect 28089 19805 28123 19839
rect 28733 19805 28767 19839
rect 32045 19805 32079 19839
rect 36277 19805 36311 19839
rect 11805 19737 11839 19771
rect 11897 19737 11931 19771
rect 12817 19737 12851 19771
rect 14657 19737 14691 19771
rect 19533 19737 19567 19771
rect 19625 19737 19659 19771
rect 26709 19737 26743 19771
rect 32229 19737 32263 19771
rect 35081 19737 35115 19771
rect 13277 19669 13311 19703
rect 20729 19669 20763 19703
rect 21373 19465 21407 19499
rect 26249 19465 26283 19499
rect 13093 19397 13127 19431
rect 13185 19397 13219 19431
rect 16957 19397 16991 19431
rect 17049 19397 17083 19431
rect 19257 19397 19291 19431
rect 22201 19397 22235 19431
rect 25605 19397 25639 19431
rect 27261 19397 27295 19431
rect 29929 19397 29963 19431
rect 30665 19397 30699 19431
rect 31585 19397 31619 19431
rect 34161 19397 34195 19431
rect 34805 19397 34839 19431
rect 36277 19397 36311 19431
rect 1869 19329 1903 19363
rect 9781 19329 9815 19363
rect 9873 19329 9907 19363
rect 20637 19329 20671 19363
rect 21281 19329 21315 19363
rect 25513 19329 25547 19363
rect 26157 19329 26191 19363
rect 27169 19329 27203 19363
rect 27997 19329 28031 19363
rect 28917 19329 28951 19363
rect 29193 19329 29227 19363
rect 29837 19329 29871 19363
rect 32321 19329 32355 19363
rect 36185 19329 36219 19363
rect 37749 19329 37783 19363
rect 1593 19261 1627 19295
rect 13737 19261 13771 19295
rect 19165 19261 19199 19295
rect 19441 19261 19475 19295
rect 20729 19261 20763 19295
rect 22109 19261 22143 19295
rect 28273 19261 28307 19295
rect 30573 19261 30607 19295
rect 32505 19261 32539 19295
rect 34713 19261 34747 19295
rect 34989 19261 35023 19295
rect 37473 19261 37507 19295
rect 17509 19193 17543 19227
rect 22661 19193 22695 19227
rect 1777 18921 1811 18955
rect 13645 18921 13679 18955
rect 18429 18921 18463 18955
rect 19533 18921 19567 18955
rect 29837 18921 29871 18955
rect 31125 18921 31159 18955
rect 31769 18921 31803 18955
rect 33701 18921 33735 18955
rect 36921 18921 36955 18955
rect 38209 18921 38243 18955
rect 15117 18853 15151 18887
rect 32413 18853 32447 18887
rect 37565 18853 37599 18887
rect 14565 18785 14599 18819
rect 16589 18785 16623 18819
rect 17601 18785 17635 18819
rect 25881 18785 25915 18819
rect 35633 18785 35667 18819
rect 1961 18717 1995 18751
rect 11805 18717 11839 18751
rect 13553 18717 13587 18751
rect 18337 18717 18371 18751
rect 19441 18717 19475 18751
rect 25145 18717 25179 18751
rect 27445 18717 27479 18751
rect 28549 18717 28583 18751
rect 29745 18717 29779 18751
rect 30389 18717 30423 18751
rect 31033 18717 31067 18751
rect 31677 18719 31711 18753
rect 32321 18717 32355 18751
rect 32965 18717 32999 18751
rect 33609 18717 33643 18751
rect 36829 18717 36863 18751
rect 37473 18717 37507 18751
rect 38117 18717 38151 18751
rect 10609 18649 10643 18683
rect 10701 18649 10735 18683
rect 11253 18649 11287 18683
rect 14657 18649 14691 18683
rect 16681 18649 16715 18683
rect 25973 18649 26007 18683
rect 26893 18649 26927 18683
rect 27905 18649 27939 18683
rect 33057 18649 33091 18683
rect 35357 18649 35391 18683
rect 35449 18649 35483 18683
rect 11897 18581 11931 18615
rect 25237 18581 25271 18615
rect 28641 18581 28675 18615
rect 30481 18581 30515 18615
rect 1593 18377 1627 18411
rect 16037 18377 16071 18411
rect 17509 18377 17543 18411
rect 28457 18377 28491 18411
rect 29101 18377 29135 18411
rect 31585 18377 31619 18411
rect 32413 18377 32447 18411
rect 34345 18377 34379 18411
rect 34989 18377 35023 18411
rect 35633 18377 35667 18411
rect 36277 18377 36311 18411
rect 37473 18377 37507 18411
rect 12357 18309 12391 18343
rect 12449 18309 12483 18343
rect 14473 18309 14507 18343
rect 19809 18309 19843 18343
rect 19901 18309 19935 18343
rect 20821 18309 20855 18343
rect 27353 18309 27387 18343
rect 30021 18309 30055 18343
rect 30113 18309 30147 18343
rect 33701 18309 33735 18343
rect 1777 18241 1811 18275
rect 14381 18241 14415 18275
rect 15945 18241 15979 18275
rect 17417 18241 17451 18275
rect 24777 18241 24811 18275
rect 26249 18241 26283 18275
rect 28365 18241 28399 18275
rect 29009 18241 29043 18275
rect 31493 18241 31527 18275
rect 32321 18241 32355 18275
rect 32965 18241 32999 18275
rect 33609 18241 33643 18275
rect 34253 18241 34287 18275
rect 34897 18241 34931 18275
rect 35541 18241 35575 18275
rect 36185 18241 36219 18275
rect 37657 18241 37691 18275
rect 38117 18241 38151 18275
rect 13369 18173 13403 18207
rect 25329 18173 25363 18207
rect 27261 18173 27295 18207
rect 27537 18173 27571 18207
rect 30389 18173 30423 18207
rect 38209 18105 38243 18139
rect 26341 18037 26375 18071
rect 33057 18037 33091 18071
rect 4077 17833 4111 17867
rect 17785 17833 17819 17867
rect 29837 17833 29871 17867
rect 35633 17833 35667 17867
rect 36921 17833 36955 17867
rect 37565 17833 37599 17867
rect 18429 17765 18463 17799
rect 30481 17765 30515 17799
rect 34989 17765 35023 17799
rect 10241 17697 10275 17731
rect 12081 17697 12115 17731
rect 20913 17697 20947 17731
rect 22937 17697 22971 17731
rect 27445 17697 27479 17731
rect 31585 17697 31619 17731
rect 31953 17697 31987 17731
rect 33977 17697 34011 17731
rect 38209 17697 38243 17731
rect 4261 17629 4295 17663
rect 11253 17629 11287 17663
rect 17693 17629 17727 17663
rect 18337 17629 18371 17663
rect 19441 17629 19475 17663
rect 20085 17629 20119 17663
rect 21557 17629 21591 17663
rect 26709 17629 26743 17663
rect 28089 17629 28123 17663
rect 28549 17629 28583 17663
rect 29745 17629 29779 17663
rect 30389 17629 30423 17663
rect 34897 17629 34931 17663
rect 35541 17629 35575 17663
rect 36185 17629 36219 17663
rect 36829 17629 36863 17663
rect 37473 17629 37507 17663
rect 38117 17629 38151 17663
rect 9965 17561 9999 17595
rect 10057 17561 10091 17595
rect 12173 17561 12207 17595
rect 12725 17561 12759 17595
rect 19533 17561 19567 17595
rect 21005 17561 21039 17595
rect 22661 17561 22695 17595
rect 22753 17561 22787 17595
rect 27514 17561 27548 17595
rect 28641 17561 28675 17595
rect 31677 17561 31711 17595
rect 33149 17561 33183 17595
rect 33241 17561 33275 17595
rect 11069 17493 11103 17527
rect 20177 17493 20211 17527
rect 26801 17493 26835 17527
rect 36277 17493 36311 17527
rect 13093 17289 13127 17323
rect 17509 17289 17543 17323
rect 20177 17289 20211 17323
rect 21373 17289 21407 17323
rect 27261 17289 27295 17323
rect 30849 17289 30883 17323
rect 9229 17221 9263 17255
rect 10149 17221 10183 17255
rect 10241 17221 10275 17255
rect 14289 17221 14323 17255
rect 28273 17221 28307 17255
rect 29377 17221 29411 17255
rect 29469 17221 29503 17255
rect 31585 17221 31619 17255
rect 32689 17221 32723 17255
rect 34253 17221 34287 17255
rect 35817 17221 35851 17255
rect 37657 17221 37691 17255
rect 1869 17153 1903 17187
rect 9137 17153 9171 17187
rect 12633 17153 12667 17187
rect 13277 17153 13311 17187
rect 14197 17153 14231 17187
rect 17417 17153 17451 17187
rect 20085 17153 20119 17187
rect 21281 17153 21315 17187
rect 22293 17153 22327 17187
rect 25421 17153 25455 17187
rect 27169 17153 27203 17187
rect 31493 17153 31527 17187
rect 1593 17085 1627 17119
rect 10977 17085 11011 17119
rect 23305 17085 23339 17119
rect 23489 17085 23523 17119
rect 28181 17085 28215 17119
rect 28457 17085 28491 17119
rect 29653 17085 29687 17119
rect 32597 17085 32631 17119
rect 32873 17085 32907 17119
rect 34161 17085 34195 17119
rect 34437 17085 34471 17119
rect 35725 17085 35759 17119
rect 36001 17085 36035 17119
rect 37565 17085 37599 17119
rect 38209 17085 38243 17119
rect 22109 17017 22143 17051
rect 23949 17017 23983 17051
rect 12449 16949 12483 16983
rect 25513 16949 25547 16983
rect 22385 16745 22419 16779
rect 27077 16745 27111 16779
rect 29837 16745 29871 16779
rect 20821 16677 20855 16711
rect 28641 16677 28675 16711
rect 15945 16609 15979 16643
rect 16957 16609 16991 16643
rect 23029 16609 23063 16643
rect 25513 16609 25547 16643
rect 35817 16609 35851 16643
rect 36369 16609 36403 16643
rect 10149 16541 10183 16575
rect 12633 16541 12667 16575
rect 17417 16541 17451 16575
rect 19901 16541 19935 16575
rect 21557 16541 21591 16575
rect 22293 16541 22327 16575
rect 26985 16541 27019 16575
rect 29745 16541 29779 16575
rect 30389 16541 30423 16575
rect 30481 16541 30515 16575
rect 31033 16541 31067 16575
rect 31125 16541 31159 16575
rect 31677 16541 31711 16575
rect 32321 16541 32355 16575
rect 32965 16541 32999 16575
rect 33609 16541 33643 16575
rect 34897 16541 34931 16575
rect 37381 16541 37415 16575
rect 38025 16541 38059 16575
rect 10241 16473 10275 16507
rect 16037 16473 16071 16507
rect 19993 16473 20027 16507
rect 20637 16473 20671 16507
rect 23121 16473 23155 16507
rect 24041 16473 24075 16507
rect 25605 16473 25639 16507
rect 26525 16473 26559 16507
rect 28089 16473 28123 16507
rect 28181 16473 28215 16507
rect 33057 16473 33091 16507
rect 35909 16473 35943 16507
rect 38117 16473 38151 16507
rect 12449 16405 12483 16439
rect 17509 16405 17543 16439
rect 21373 16405 21407 16439
rect 31769 16405 31803 16439
rect 32413 16405 32447 16439
rect 33701 16405 33735 16439
rect 34989 16405 35023 16439
rect 37473 16405 37507 16439
rect 10977 16201 11011 16235
rect 19533 16201 19567 16235
rect 29009 16201 29043 16235
rect 29653 16201 29687 16235
rect 35817 16201 35851 16235
rect 36461 16201 36495 16235
rect 12541 16133 12575 16167
rect 13461 16133 13495 16167
rect 14381 16133 14415 16167
rect 17049 16133 17083 16167
rect 22753 16133 22787 16167
rect 32505 16133 32539 16167
rect 34069 16133 34103 16167
rect 35173 16133 35207 16167
rect 37749 16133 37783 16167
rect 1593 16065 1627 16099
rect 10885 16065 10919 16099
rect 19441 16065 19475 16099
rect 20269 16065 20303 16099
rect 20729 16065 20763 16099
rect 28273 16065 28307 16099
rect 28917 16065 28951 16099
rect 29561 16065 29595 16099
rect 30205 16065 30239 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 35081 16065 35115 16099
rect 35725 16065 35759 16099
rect 36369 16065 36403 16099
rect 10241 15997 10275 16031
rect 12449 15997 12483 16031
rect 14289 15997 14323 16031
rect 14565 15997 14599 16031
rect 16957 15997 16991 16031
rect 17233 15997 17267 16031
rect 22662 15997 22696 16031
rect 22937 15997 22971 16031
rect 32413 15997 32447 16031
rect 33333 15997 33367 16031
rect 33977 15997 34011 16031
rect 34621 15997 34655 16031
rect 37657 15997 37691 16031
rect 38301 15997 38335 16031
rect 1777 15861 1811 15895
rect 20085 15861 20119 15895
rect 20821 15861 20855 15895
rect 28365 15861 28399 15895
rect 30297 15861 30331 15895
rect 31769 15861 31803 15895
rect 14381 15657 14415 15691
rect 19809 15657 19843 15691
rect 28825 15657 28859 15691
rect 33885 15657 33919 15691
rect 34989 15657 35023 15691
rect 37381 15657 37415 15691
rect 11345 15589 11379 15623
rect 30113 15589 30147 15623
rect 30941 15589 30975 15623
rect 33241 15589 33275 15623
rect 10241 15521 10275 15555
rect 10425 15521 10459 15555
rect 28089 15521 28123 15555
rect 29929 15521 29963 15555
rect 32689 15521 32723 15555
rect 35909 15521 35943 15555
rect 11529 15453 11563 15487
rect 13001 15453 13035 15487
rect 14289 15453 14323 15487
rect 18153 15453 18187 15487
rect 19993 15453 20027 15487
rect 20637 15453 20671 15487
rect 21465 15453 21499 15487
rect 25237 15453 25271 15487
rect 26433 15453 26467 15487
rect 27997 15453 28031 15487
rect 29745 15453 29779 15487
rect 30849 15453 30883 15487
rect 31677 15453 31711 15487
rect 33793 15453 33827 15487
rect 34897 15453 34931 15487
rect 37565 15453 37599 15487
rect 38025 15453 38059 15487
rect 20729 15385 20763 15419
rect 28733 15385 28767 15419
rect 32781 15385 32815 15419
rect 36001 15385 36035 15419
rect 36553 15385 36587 15419
rect 10885 15317 10919 15351
rect 12817 15317 12851 15351
rect 18245 15317 18279 15351
rect 21281 15317 21315 15351
rect 25053 15317 25087 15351
rect 26525 15317 26559 15351
rect 31493 15317 31527 15351
rect 38209 15317 38243 15351
rect 10793 15113 10827 15147
rect 11713 15113 11747 15147
rect 14933 15113 14967 15147
rect 26525 15113 26559 15147
rect 35633 15113 35667 15147
rect 37565 15113 37599 15147
rect 38209 15113 38243 15147
rect 13277 15045 13311 15079
rect 22109 15045 22143 15079
rect 22937 15045 22971 15079
rect 27353 15045 27387 15079
rect 29193 15045 29227 15079
rect 32505 15045 32539 15079
rect 9597 14977 9631 15011
rect 10701 14977 10735 15011
rect 11897 14977 11931 15011
rect 17325 14977 17359 15011
rect 20361 14977 20395 15011
rect 20545 14977 20579 15011
rect 22017 14977 22051 15011
rect 26433 14977 26467 15011
rect 30573 14977 30607 15011
rect 31401 14977 31435 15011
rect 33057 14977 33091 15011
rect 34161 14977 34195 15011
rect 34897 14977 34931 15011
rect 35541 14977 35575 15011
rect 36185 14977 36219 15011
rect 37473 14977 37507 15011
rect 38117 14977 38151 15011
rect 13185 14909 13219 14943
rect 13461 14909 13495 14943
rect 14289 14909 14323 14943
rect 14473 14909 14507 14943
rect 22845 14909 22879 14943
rect 23857 14909 23891 14943
rect 27261 14909 27295 14943
rect 27629 14909 27663 14943
rect 29101 14909 29135 14943
rect 29745 14909 29779 14943
rect 32413 14909 32447 14943
rect 33517 14909 33551 14943
rect 34989 14909 35023 14943
rect 9689 14841 9723 14875
rect 20729 14841 20763 14875
rect 17417 14773 17451 14807
rect 30665 14773 30699 14807
rect 31217 14773 31251 14807
rect 34253 14773 34287 14807
rect 36277 14773 36311 14807
rect 14381 14569 14415 14603
rect 28273 14569 28307 14603
rect 31125 14569 31159 14603
rect 32045 14569 32079 14603
rect 34989 14569 35023 14603
rect 36369 14569 36403 14603
rect 37841 14569 37875 14603
rect 14933 14501 14967 14535
rect 37197 14501 37231 14535
rect 17049 14433 17083 14467
rect 17877 14433 17911 14467
rect 25329 14433 25363 14467
rect 26985 14433 27019 14467
rect 27261 14433 27295 14467
rect 31677 14433 31711 14467
rect 31861 14433 31895 14467
rect 33609 14433 33643 14467
rect 36185 14433 36219 14467
rect 1593 14365 1627 14399
rect 14289 14365 14323 14399
rect 15117 14365 15151 14399
rect 18705 14365 18739 14399
rect 22477 14365 22511 14399
rect 28181 14365 28215 14399
rect 28825 14365 28859 14399
rect 29745 14365 29779 14399
rect 30389 14365 30423 14399
rect 31033 14365 31067 14399
rect 34897 14365 34931 14399
rect 36001 14365 36035 14399
rect 37105 14365 37139 14399
rect 37749 14365 37783 14399
rect 17141 14297 17175 14331
rect 25053 14297 25087 14331
rect 25145 14297 25179 14331
rect 27077 14297 27111 14331
rect 33333 14297 33367 14331
rect 33425 14297 33459 14331
rect 1777 14229 1811 14263
rect 18521 14229 18555 14263
rect 22569 14229 22603 14263
rect 28917 14229 28951 14263
rect 29837 14229 29871 14263
rect 30481 14229 30515 14263
rect 1593 14025 1627 14059
rect 14381 14025 14415 14059
rect 19257 14025 19291 14059
rect 22201 14025 22235 14059
rect 38209 14025 38243 14059
rect 13369 13957 13403 13991
rect 17141 13957 17175 13991
rect 17233 13957 17267 13991
rect 23397 13957 23431 13991
rect 23489 13957 23523 13991
rect 25697 13957 25731 13991
rect 25789 13957 25823 13991
rect 27813 13957 27847 13991
rect 29193 13957 29227 13991
rect 30849 13957 30883 13991
rect 33977 13957 34011 13991
rect 35541 13957 35575 13991
rect 36461 13957 36495 13991
rect 37565 13957 37599 13991
rect 1777 13889 1811 13923
rect 10701 13889 10735 13923
rect 14565 13889 14599 13923
rect 15209 13889 15243 13923
rect 19901 13889 19935 13923
rect 20821 13889 20855 13923
rect 22109 13889 22143 13923
rect 27169 13889 27203 13923
rect 28549 13889 28583 13923
rect 28733 13889 28767 13923
rect 29745 13889 29779 13923
rect 32321 13889 32355 13923
rect 37473 13889 37507 13923
rect 38117 13889 38151 13923
rect 10793 13821 10827 13855
rect 13277 13821 13311 13855
rect 13737 13821 13771 13855
rect 17969 13821 18003 13855
rect 18613 13821 18647 13855
rect 18797 13821 18831 13855
rect 23673 13821 23707 13855
rect 26157 13821 26191 13855
rect 27353 13821 27387 13855
rect 29837 13821 29871 13855
rect 30757 13821 30791 13855
rect 31677 13821 31711 13855
rect 32413 13821 32447 13855
rect 33149 13821 33183 13855
rect 33885 13821 33919 13855
rect 34161 13821 34195 13855
rect 35449 13821 35483 13855
rect 15025 13753 15059 13787
rect 19717 13685 19751 13719
rect 20913 13685 20947 13719
rect 14933 13481 14967 13515
rect 17877 13481 17911 13515
rect 19441 13481 19475 13515
rect 20729 13481 20763 13515
rect 26801 13481 26835 13515
rect 32873 13481 32907 13515
rect 34161 13481 34195 13515
rect 34989 13481 35023 13515
rect 36461 13481 36495 13515
rect 37289 13481 37323 13515
rect 25605 13413 25639 13447
rect 26249 13413 26283 13447
rect 32137 13413 32171 13447
rect 33425 13413 33459 13447
rect 13277 13345 13311 13379
rect 14565 13345 14599 13379
rect 20085 13345 20119 13379
rect 20269 13345 20303 13379
rect 36277 13345 36311 13379
rect 14749 13277 14783 13311
rect 17785 13277 17819 13311
rect 19625 13277 19659 13311
rect 22845 13277 22879 13311
rect 26157 13277 26191 13311
rect 26985 13277 27019 13311
rect 27445 13277 27479 13311
rect 32321 13277 32355 13311
rect 32781 13277 32815 13311
rect 33609 13277 33643 13311
rect 34069 13277 34103 13311
rect 34897 13277 34931 13311
rect 36093 13277 36127 13311
rect 37197 13277 37231 13311
rect 38025 13277 38059 13311
rect 25053 13209 25087 13243
rect 25145 13209 25179 13243
rect 12265 13141 12299 13175
rect 22937 13141 22971 13175
rect 27537 13141 27571 13175
rect 38209 13141 38243 13175
rect 6929 12937 6963 12971
rect 9321 12937 9355 12971
rect 12817 12937 12851 12971
rect 15025 12937 15059 12971
rect 20269 12937 20303 12971
rect 26433 12937 26467 12971
rect 29377 12937 29411 12971
rect 32321 12937 32355 12971
rect 32965 12937 32999 12971
rect 34989 12937 35023 12971
rect 35633 12937 35667 12971
rect 36277 12937 36311 12971
rect 18337 12869 18371 12903
rect 18429 12869 18463 12903
rect 37749 12869 37783 12903
rect 1593 12801 1627 12835
rect 7113 12801 7147 12835
rect 9229 12801 9263 12835
rect 12173 12801 12207 12835
rect 14933 12801 14967 12835
rect 19993 12801 20027 12835
rect 22937 12801 22971 12835
rect 26617 12801 26651 12835
rect 29285 12801 29319 12835
rect 31033 12801 31067 12835
rect 32505 12801 32539 12835
rect 33149 12801 33183 12835
rect 33609 12801 33643 12835
rect 34253 12801 34287 12835
rect 34897 12801 34931 12835
rect 35541 12801 35575 12835
rect 36185 12801 36219 12835
rect 12357 12733 12391 12767
rect 18613 12733 18647 12767
rect 37657 12733 37691 12767
rect 37933 12733 37967 12767
rect 31125 12665 31159 12699
rect 33701 12665 33735 12699
rect 1777 12597 1811 12631
rect 22753 12597 22787 12631
rect 34345 12597 34379 12631
rect 12449 12393 12483 12427
rect 20085 12393 20119 12427
rect 28273 12393 28307 12427
rect 33425 12393 33459 12427
rect 34253 12393 34287 12427
rect 35357 12393 35391 12427
rect 36645 12393 36679 12427
rect 35909 12325 35943 12359
rect 17601 12257 17635 12291
rect 22661 12257 22695 12291
rect 22845 12257 22879 12291
rect 26801 12257 26835 12291
rect 37289 12257 37323 12291
rect 37565 12257 37599 12291
rect 11989 12189 12023 12223
rect 12633 12189 12667 12223
rect 13461 12189 13495 12223
rect 19993 12189 20027 12223
rect 28181 12189 28215 12223
rect 33333 12189 33367 12223
rect 34161 12189 34195 12223
rect 35265 12189 35299 12223
rect 36093 12189 36127 12223
rect 36553 12189 36587 12223
rect 16957 12121 16991 12155
rect 17049 12121 17083 12155
rect 26893 12121 26927 12155
rect 27445 12121 27479 12155
rect 37381 12121 37415 12155
rect 11805 12053 11839 12087
rect 13553 12053 13587 12087
rect 23305 12053 23339 12087
rect 9597 11849 9631 11883
rect 14749 11849 14783 11883
rect 16957 11849 16991 11883
rect 19533 11849 19567 11883
rect 21465 11849 21499 11883
rect 23949 11849 23983 11883
rect 34897 11849 34931 11883
rect 35449 11849 35483 11883
rect 37565 11849 37599 11883
rect 25237 11781 25271 11815
rect 26341 11781 26375 11815
rect 36277 11781 36311 11815
rect 36369 11781 36403 11815
rect 9505 11713 9539 11747
rect 14657 11713 14691 11747
rect 16865 11713 16899 11747
rect 17509 11713 17543 11747
rect 18797 11713 18831 11747
rect 19441 11713 19475 11747
rect 23857 11713 23891 11747
rect 26249 11713 26283 11747
rect 33517 11713 33551 11747
rect 34345 11713 34379 11747
rect 34805 11713 34839 11747
rect 37473 11713 37507 11747
rect 38301 11713 38335 11747
rect 20821 11645 20855 11679
rect 21005 11645 21039 11679
rect 22753 11645 22787 11679
rect 22937 11645 22971 11679
rect 25145 11645 25179 11679
rect 25421 11645 25455 11679
rect 18889 11577 18923 11611
rect 33609 11577 33643 11611
rect 36829 11577 36863 11611
rect 38117 11577 38151 11611
rect 17601 11509 17635 11543
rect 23121 11509 23155 11543
rect 34161 11509 34195 11543
rect 17417 11305 17451 11339
rect 22845 11305 22879 11339
rect 34161 11305 34195 11339
rect 36737 11305 36771 11339
rect 1593 11237 1627 11271
rect 35357 11237 35391 11271
rect 9229 11169 9263 11203
rect 19533 11169 19567 11203
rect 21097 11169 21131 11203
rect 29193 11169 29227 11203
rect 37749 11169 37783 11203
rect 1777 11101 1811 11135
rect 9137 11101 9171 11135
rect 16405 11101 16439 11135
rect 17325 11101 17359 11135
rect 21925 11101 21959 11135
rect 23029 11101 23063 11135
rect 32045 11101 32079 11135
rect 34345 11101 34379 11135
rect 35541 11101 35575 11135
rect 36001 11101 36035 11135
rect 36645 11101 36679 11135
rect 16497 11033 16531 11067
rect 19625 11033 19659 11067
rect 20177 11033 20211 11067
rect 28181 11033 28215 11067
rect 28273 11033 28307 11067
rect 32137 11033 32171 11067
rect 36093 11033 36127 11067
rect 21741 10965 21775 10999
rect 1593 10761 1627 10795
rect 20821 10761 20855 10795
rect 32597 10761 32631 10795
rect 35909 10761 35943 10795
rect 36645 10761 36679 10795
rect 13001 10693 13035 10727
rect 17049 10693 17083 10727
rect 17601 10693 17635 10727
rect 34529 10693 34563 10727
rect 1777 10625 1811 10659
rect 21005 10625 21039 10659
rect 25053 10625 25087 10659
rect 28825 10625 28859 10659
rect 32505 10625 32539 10659
rect 34437 10625 34471 10659
rect 35265 10625 35299 10659
rect 36093 10625 36127 10659
rect 36553 10625 36587 10659
rect 38025 10625 38059 10659
rect 12909 10557 12943 10591
rect 13461 10557 13495 10591
rect 16957 10557 16991 10591
rect 24409 10557 24443 10591
rect 35357 10557 35391 10591
rect 25145 10421 25179 10455
rect 28917 10421 28951 10455
rect 38209 10421 38243 10455
rect 7941 10217 7975 10251
rect 25881 10217 25915 10251
rect 36737 10217 36771 10251
rect 37841 10149 37875 10183
rect 21741 10081 21775 10115
rect 24685 10081 24719 10115
rect 24961 10081 24995 10115
rect 7849 10013 7883 10047
rect 9505 10013 9539 10047
rect 19717 10013 19751 10047
rect 21925 10013 21959 10047
rect 25789 10013 25823 10047
rect 36185 10013 36219 10047
rect 36645 10013 36679 10047
rect 37749 10013 37783 10047
rect 24777 9945 24811 9979
rect 9597 9877 9631 9911
rect 19809 9877 19843 9911
rect 21005 9877 21039 9911
rect 22385 9877 22419 9911
rect 36001 9877 36035 9911
rect 4813 9605 4847 9639
rect 9137 9605 9171 9639
rect 22109 9605 22143 9639
rect 25421 9605 25455 9639
rect 30389 9605 30423 9639
rect 31309 9605 31343 9639
rect 36737 9605 36771 9639
rect 4721 9537 4755 9571
rect 6929 9537 6963 9571
rect 9045 9537 9079 9571
rect 18981 9537 19015 9571
rect 20821 9537 20855 9571
rect 22017 9537 22051 9571
rect 25329 9537 25363 9571
rect 27445 9537 27479 9571
rect 38025 9537 38059 9571
rect 21005 9469 21039 9503
rect 30297 9469 30331 9503
rect 19073 9401 19107 9435
rect 37841 9401 37875 9435
rect 7021 9333 7055 9367
rect 21189 9333 21223 9367
rect 27537 9333 27571 9367
rect 1593 9129 1627 9163
rect 20453 9129 20487 9163
rect 1777 8925 1811 8959
rect 18705 8925 18739 8959
rect 19993 8925 20027 8959
rect 20637 8925 20671 8959
rect 28089 8925 28123 8959
rect 38025 8925 38059 8959
rect 18797 8789 18831 8823
rect 19809 8789 19843 8823
rect 27905 8789 27939 8823
rect 38209 8789 38243 8823
rect 19257 8585 19291 8619
rect 25237 8585 25271 8619
rect 38117 8585 38151 8619
rect 7113 8449 7147 8483
rect 9229 8449 9263 8483
rect 19441 8449 19475 8483
rect 25145 8449 25179 8483
rect 37657 8449 37691 8483
rect 38301 8449 38335 8483
rect 6929 8313 6963 8347
rect 9321 8313 9355 8347
rect 37473 8313 37507 8347
rect 10977 8041 11011 8075
rect 2237 7905 2271 7939
rect 1593 7837 1627 7871
rect 10885 7837 10919 7871
rect 29009 7837 29043 7871
rect 38025 7837 38059 7871
rect 1777 7701 1811 7735
rect 28825 7701 28859 7735
rect 38209 7701 38243 7735
rect 38117 7497 38151 7531
rect 1869 7361 1903 7395
rect 17785 7361 17819 7395
rect 33149 7361 33183 7395
rect 38301 7361 38335 7395
rect 1593 7293 1627 7327
rect 17601 7157 17635 7191
rect 32965 7157 32999 7191
rect 7941 6273 7975 6307
rect 7757 6069 7791 6103
rect 8401 5865 8435 5899
rect 1869 5729 1903 5763
rect 1593 5661 1627 5695
rect 8309 5661 8343 5695
rect 29929 5661 29963 5695
rect 38025 5661 38059 5695
rect 29745 5525 29779 5559
rect 38209 5525 38243 5559
rect 1593 4777 1627 4811
rect 1777 4573 1811 4607
rect 32597 4573 32631 4607
rect 38301 4573 38335 4607
rect 32413 4437 32447 4471
rect 1777 4097 1811 4131
rect 36737 4097 36771 4131
rect 38025 4097 38059 4131
rect 1593 3961 1627 3995
rect 36829 3893 36863 3927
rect 38209 3893 38243 3927
rect 2329 3689 2363 3723
rect 36829 3689 36863 3723
rect 37749 3553 37783 3587
rect 1593 3485 1627 3519
rect 2513 3485 2547 3519
rect 37013 3485 37047 3519
rect 37473 3485 37507 3519
rect 1777 3349 1811 3383
rect 35541 3145 35575 3179
rect 36737 3145 36771 3179
rect 2145 3009 2179 3043
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 3985 3009 4019 3043
rect 16313 3009 16347 3043
rect 17049 3009 17083 3043
rect 33057 3009 33091 3043
rect 35725 3009 35759 3043
rect 36921 3009 36955 3043
rect 37473 3009 37507 3043
rect 2697 2805 2731 2839
rect 4169 2805 4203 2839
rect 16129 2805 16163 2839
rect 16865 2805 16899 2839
rect 32873 2805 32907 2839
rect 37657 2805 37691 2839
rect 2973 2601 3007 2635
rect 6561 2601 6595 2635
rect 7205 2601 7239 2635
rect 8401 2601 8435 2635
rect 14289 2601 14323 2635
rect 19441 2601 19475 2635
rect 20315 2601 20349 2635
rect 23305 2601 23339 2635
rect 24593 2601 24627 2635
rect 27813 2601 27847 2635
rect 29745 2601 29779 2635
rect 35081 2601 35115 2635
rect 2329 2533 2363 2567
rect 5273 2533 5307 2567
rect 22017 2533 22051 2567
rect 27169 2533 27203 2567
rect 36093 2533 36127 2567
rect 4261 2465 4295 2499
rect 10609 2465 10643 2499
rect 26065 2465 26099 2499
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 3157 2397 3191 2431
rect 3985 2397 4019 2431
rect 5457 2397 5491 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 8585 2397 8619 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 13185 2397 13219 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 18153 2397 18187 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 22201 2397 22235 2431
rect 22845 2397 22879 2431
rect 23489 2397 23523 2431
rect 24777 2397 24811 2431
rect 25789 2397 25823 2431
rect 27353 2397 27387 2431
rect 27997 2397 28031 2431
rect 29929 2397 29963 2431
rect 30389 2397 30423 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 35909 2397 35943 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 34989 2329 35023 2363
rect 1777 2261 1811 2295
rect 9781 2261 9815 2295
rect 13001 2261 13035 2295
rect 15117 2261 15151 2295
rect 16221 2261 16255 2295
rect 17049 2261 17083 2295
rect 18337 2261 18371 2295
rect 22661 2261 22695 2295
rect 30573 2261 30607 2295
rect 31309 2261 31343 2295
rect 32505 2261 32539 2295
rect 33793 2261 33827 2295
rect 36829 2261 36863 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 19334 37680 19340 37732
rect 19392 37720 19398 37732
rect 20346 37720 20352 37732
rect 19392 37692 20352 37720
rect 19392 37680 19398 37692
rect 20346 37680 20352 37692
rect 20404 37680 20410 37732
rect 17218 37612 17224 37664
rect 17276 37652 17282 37664
rect 27890 37652 27896 37664
rect 17276 37624 27896 37652
rect 17276 37612 17282 37624
rect 27890 37612 27896 37624
rect 27948 37612 27954 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 7742 37408 7748 37460
rect 7800 37448 7806 37460
rect 17218 37448 17224 37460
rect 7800 37420 17224 37448
rect 7800 37408 7806 37420
rect 17218 37408 17224 37420
rect 17276 37408 17282 37460
rect 19686 37451 19744 37457
rect 19686 37448 19698 37451
rect 18800 37420 19698 37448
rect 18800 37392 18828 37420
rect 19686 37417 19698 37420
rect 19732 37448 19744 37451
rect 20254 37448 20260 37460
rect 19732 37420 20260 37448
rect 19732 37417 19744 37420
rect 19686 37411 19744 37417
rect 20254 37408 20260 37420
rect 20312 37408 20318 37460
rect 658 37340 664 37392
rect 716 37380 722 37392
rect 4614 37380 4620 37392
rect 716 37352 4620 37380
rect 716 37340 722 37352
rect 4614 37340 4620 37352
rect 4672 37340 4678 37392
rect 8389 37383 8447 37389
rect 8389 37349 8401 37383
rect 8435 37349 8447 37383
rect 8389 37343 8447 37349
rect 10413 37383 10471 37389
rect 10413 37349 10425 37383
rect 10459 37380 10471 37383
rect 15194 37380 15200 37392
rect 10459 37352 15200 37380
rect 10459 37349 10471 37352
rect 10413 37343 10471 37349
rect 1578 37312 1584 37324
rect 1539 37284 1584 37312
rect 1578 37272 1584 37284
rect 1636 37272 1642 37324
rect 5166 37312 5172 37324
rect 5127 37284 5172 37312
rect 5166 37272 5172 37284
rect 5224 37272 5230 37324
rect 5810 37272 5816 37324
rect 5868 37312 5874 37324
rect 6549 37315 6607 37321
rect 6549 37312 6561 37315
rect 5868 37284 6561 37312
rect 5868 37272 5874 37284
rect 6549 37281 6561 37284
rect 6595 37281 6607 37315
rect 6549 37275 6607 37281
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 1946 37244 1952 37256
rect 1903 37216 1952 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 1946 37204 1952 37216
rect 2004 37204 2010 37256
rect 2869 37247 2927 37253
rect 2869 37213 2881 37247
rect 2915 37244 2927 37247
rect 3786 37244 3792 37256
rect 2915 37216 3792 37244
rect 2915 37213 2927 37216
rect 2869 37207 2927 37213
rect 3786 37204 3792 37216
rect 3844 37204 3850 37256
rect 3973 37247 4031 37253
rect 3973 37213 3985 37247
rect 4019 37244 4031 37247
rect 4062 37244 4068 37256
rect 4019 37216 4068 37244
rect 4019 37213 4031 37216
rect 3973 37207 4031 37213
rect 4062 37204 4068 37216
rect 4120 37204 4126 37256
rect 5442 37244 5448 37256
rect 5403 37216 5448 37244
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 6638 37204 6644 37256
rect 6696 37244 6702 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6696 37216 6837 37244
rect 6696 37204 6702 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 8404 37244 8432 37343
rect 15194 37340 15200 37352
rect 15252 37340 15258 37392
rect 18414 37380 18420 37392
rect 18375 37352 18420 37380
rect 18414 37340 18420 37352
rect 18472 37340 18478 37392
rect 18782 37380 18788 37392
rect 18743 37352 18788 37380
rect 18782 37340 18788 37352
rect 18840 37340 18846 37392
rect 23385 37383 23443 37389
rect 23385 37349 23397 37383
rect 23431 37349 23443 37383
rect 23385 37343 23443 37349
rect 10226 37312 10232 37324
rect 9784 37284 10232 37312
rect 8478 37244 8484 37256
rect 8404 37216 8484 37244
rect 6825 37207 6883 37213
rect 8478 37204 8484 37216
rect 8536 37204 8542 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37244 8631 37247
rect 9784 37244 9812 37284
rect 10226 37272 10232 37284
rect 10284 37272 10290 37324
rect 11606 37312 11612 37324
rect 11072 37284 11612 37312
rect 8619 37216 9812 37244
rect 9861 37247 9919 37253
rect 8619 37213 8631 37216
rect 8573 37207 8631 37213
rect 9861 37213 9873 37247
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 5074 37136 5080 37188
rect 5132 37176 5138 37188
rect 9122 37176 9128 37188
rect 5132 37148 9128 37176
rect 5132 37136 5138 37148
rect 9122 37136 9128 37148
rect 9180 37136 9186 37188
rect 9876 37176 9904 37207
rect 10042 37204 10048 37256
rect 10100 37244 10106 37256
rect 10321 37247 10379 37253
rect 10321 37244 10333 37247
rect 10100 37216 10333 37244
rect 10100 37204 10106 37216
rect 10321 37213 10333 37216
rect 10367 37213 10379 37247
rect 11072 37244 11100 37284
rect 11606 37272 11612 37284
rect 11664 37272 11670 37324
rect 11790 37312 11796 37324
rect 11751 37284 11796 37312
rect 11790 37272 11796 37284
rect 11848 37272 11854 37324
rect 12250 37272 12256 37324
rect 12308 37312 12314 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 12308 37284 12357 37312
rect 12308 37272 12314 37284
rect 12345 37281 12357 37284
rect 12391 37281 12403 37315
rect 12345 37275 12403 37281
rect 15473 37315 15531 37321
rect 15473 37281 15485 37315
rect 15519 37312 15531 37315
rect 16114 37312 16120 37324
rect 15519 37284 16120 37312
rect 15519 37281 15531 37284
rect 15473 37275 15531 37281
rect 16114 37272 16120 37284
rect 16172 37272 16178 37324
rect 16482 37272 16488 37324
rect 16540 37312 16546 37324
rect 22922 37312 22928 37324
rect 16540 37284 20944 37312
rect 22883 37284 22928 37312
rect 16540 37272 16546 37284
rect 10321 37207 10379 37213
rect 10428 37216 11100 37244
rect 11149 37247 11207 37253
rect 10428 37176 10456 37216
rect 11149 37213 11161 37247
rect 11195 37213 11207 37247
rect 11698 37244 11704 37256
rect 11659 37216 11704 37244
rect 11149 37207 11207 37213
rect 9508 37148 9812 37176
rect 9876 37148 10456 37176
rect 11164 37176 11192 37207
rect 11698 37204 11704 37216
rect 11756 37204 11762 37256
rect 12434 37244 12440 37256
rect 11808 37216 12440 37244
rect 11808 37176 11836 37216
rect 12434 37204 12440 37216
rect 12492 37204 12498 37256
rect 12621 37247 12679 37253
rect 12621 37213 12633 37247
rect 12667 37244 12679 37247
rect 12894 37244 12900 37256
rect 12667 37216 12900 37244
rect 12667 37213 12679 37216
rect 12621 37207 12679 37213
rect 12894 37204 12900 37216
rect 12952 37204 12958 37256
rect 14737 37247 14795 37253
rect 14737 37213 14749 37247
rect 14783 37213 14795 37247
rect 14737 37207 14795 37213
rect 15749 37247 15807 37253
rect 15749 37213 15761 37247
rect 15795 37244 15807 37247
rect 16666 37244 16672 37256
rect 15795 37216 16672 37244
rect 15795 37213 15807 37216
rect 15749 37207 15807 37213
rect 13630 37176 13636 37188
rect 11164 37148 11836 37176
rect 11900 37148 13636 37176
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2832 37080 3065 37108
rect 2832 37068 2838 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 3053 37071 3111 37077
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3936 37080 4169 37108
rect 3936 37068 3942 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4157 37071 4215 37077
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 9508 37108 9536 37148
rect 9674 37108 9680 37120
rect 5868 37080 9536 37108
rect 9635 37080 9680 37108
rect 5868 37068 5874 37080
rect 9674 37068 9680 37080
rect 9732 37068 9738 37120
rect 9784 37108 9812 37148
rect 10226 37108 10232 37120
rect 9784 37080 10232 37108
rect 10226 37068 10232 37080
rect 10284 37068 10290 37120
rect 10965 37111 11023 37117
rect 10965 37077 10977 37111
rect 11011 37108 11023 37111
rect 11900 37108 11928 37148
rect 13630 37136 13636 37148
rect 13688 37136 13694 37188
rect 11011 37080 11928 37108
rect 11011 37077 11023 37080
rect 10965 37071 11023 37077
rect 11974 37068 11980 37120
rect 12032 37108 12038 37120
rect 14752 37108 14780 37207
rect 16666 37204 16672 37216
rect 16724 37204 16730 37256
rect 18233 37247 18291 37253
rect 18233 37244 18245 37247
rect 17788 37216 18245 37244
rect 17788 37188 17816 37216
rect 18233 37213 18245 37216
rect 18279 37213 18291 37247
rect 18233 37207 18291 37213
rect 18322 37204 18328 37256
rect 18380 37244 18386 37256
rect 18380 37216 19288 37244
rect 18380 37204 18386 37216
rect 15010 37136 15016 37188
rect 15068 37176 15074 37188
rect 16945 37179 17003 37185
rect 16945 37176 16957 37179
rect 15068 37148 16957 37176
rect 15068 37136 15074 37148
rect 16945 37145 16957 37148
rect 16991 37145 17003 37179
rect 16945 37139 17003 37145
rect 17037 37179 17095 37185
rect 17037 37145 17049 37179
rect 17083 37145 17095 37179
rect 17037 37139 17095 37145
rect 12032 37080 14780 37108
rect 12032 37068 12038 37080
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 14921 37111 14979 37117
rect 14921 37108 14933 37111
rect 14884 37080 14933 37108
rect 14884 37068 14890 37080
rect 14921 37077 14933 37080
rect 14967 37077 14979 37111
rect 14921 37071 14979 37077
rect 15102 37068 15108 37120
rect 15160 37108 15166 37120
rect 16482 37108 16488 37120
rect 15160 37080 16488 37108
rect 15160 37068 15166 37080
rect 16482 37068 16488 37080
rect 16540 37068 16546 37120
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 17052 37108 17080 37139
rect 17770 37136 17776 37188
rect 17828 37136 17834 37188
rect 17957 37179 18015 37185
rect 17957 37145 17969 37179
rect 18003 37145 18015 37179
rect 17957 37139 18015 37145
rect 16632 37080 17080 37108
rect 16632 37068 16638 37080
rect 17218 37068 17224 37120
rect 17276 37108 17282 37120
rect 17972 37108 18000 37139
rect 18414 37136 18420 37188
rect 18472 37176 18478 37188
rect 19260 37176 19288 37216
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 19392 37216 19441 37244
rect 19392 37204 19398 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 20806 37204 20812 37256
rect 20864 37204 20870 37256
rect 20916 37244 20944 37284
rect 22922 37272 22928 37284
rect 22980 37272 22986 37324
rect 23400 37312 23428 37343
rect 23124 37284 23428 37312
rect 25133 37315 25191 37321
rect 20990 37244 20996 37256
rect 20916 37216 20996 37244
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21324 37216 22201 37244
rect 21324 37204 21330 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 22612 37216 22753 37244
rect 22612 37204 22618 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 23124 37176 23152 37284
rect 25133 37281 25145 37315
rect 25179 37312 25191 37315
rect 25498 37312 25504 37324
rect 25179 37284 25504 37312
rect 25179 37281 25191 37284
rect 25133 37275 25191 37281
rect 25498 37272 25504 37284
rect 25556 37272 25562 37324
rect 25774 37272 25780 37324
rect 25832 37312 25838 37324
rect 25832 37284 26372 37312
rect 25832 37272 25838 37284
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23569 37247 23627 37253
rect 23569 37244 23581 37247
rect 23256 37216 23581 37244
rect 23256 37204 23262 37216
rect 23569 37213 23581 37216
rect 23615 37213 23627 37247
rect 23569 37207 23627 37213
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 24857 37247 24915 37253
rect 24857 37244 24869 37247
rect 24820 37216 24869 37244
rect 24820 37204 24826 37216
rect 24857 37213 24869 37216
rect 24903 37213 24915 37247
rect 24857 37207 24915 37213
rect 26234 37204 26240 37256
rect 26292 37204 26298 37256
rect 26344 37244 26372 37284
rect 26988 37284 27292 37312
rect 26988 37244 27016 37284
rect 26344 37216 27016 37244
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 27120 37216 27169 37244
rect 27120 37204 27126 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27264 37244 27292 37284
rect 29638 37272 29644 37324
rect 29696 37312 29702 37324
rect 29733 37315 29791 37321
rect 29733 37312 29745 37315
rect 29696 37284 29745 37312
rect 29696 37272 29702 37284
rect 29733 37281 29745 37284
rect 29779 37281 29791 37315
rect 29733 37275 29791 37281
rect 32677 37315 32735 37321
rect 32677 37281 32689 37315
rect 32723 37312 32735 37315
rect 34054 37312 34060 37324
rect 32723 37284 34060 37312
rect 32723 37281 32735 37284
rect 32677 37275 32735 37281
rect 34054 37272 34060 37284
rect 34112 37272 34118 37324
rect 35158 37312 35164 37324
rect 35119 37284 35164 37312
rect 35158 37272 35164 37284
rect 35216 37272 35222 37324
rect 37458 37312 37464 37324
rect 37419 37284 37464 37312
rect 37458 37272 37464 37284
rect 37516 37272 37522 37324
rect 28077 37247 28135 37253
rect 28077 37244 28089 37247
rect 27264 37216 28089 37244
rect 27157 37207 27215 37213
rect 28077 37213 28089 37216
rect 28123 37213 28135 37247
rect 28077 37207 28135 37213
rect 28721 37247 28779 37253
rect 28721 37213 28733 37247
rect 28767 37213 28779 37247
rect 30006 37244 30012 37256
rect 29967 37216 30012 37244
rect 28721 37207 28779 37213
rect 18472 37148 19196 37176
rect 19260 37148 20116 37176
rect 18472 37136 18478 37148
rect 18966 37108 18972 37120
rect 17276 37080 18972 37108
rect 17276 37068 17282 37080
rect 18966 37068 18972 37080
rect 19024 37068 19030 37120
rect 19168 37108 19196 37148
rect 19978 37108 19984 37120
rect 19168 37080 19984 37108
rect 19978 37068 19984 37080
rect 20036 37068 20042 37120
rect 20088 37108 20116 37148
rect 21008 37148 23152 37176
rect 21008 37108 21036 37148
rect 26418 37136 26424 37188
rect 26476 37176 26482 37188
rect 26476 37148 27384 37176
rect 26476 37136 26482 37148
rect 21174 37108 21180 37120
rect 20088 37080 21036 37108
rect 21135 37080 21180 37108
rect 21174 37068 21180 37080
rect 21232 37068 21238 37120
rect 22002 37108 22008 37120
rect 21963 37080 22008 37108
rect 22002 37068 22008 37080
rect 22060 37068 22066 37120
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 27356 37117 27384 37148
rect 27706 37136 27712 37188
rect 27764 37176 27770 37188
rect 28736 37176 28764 37207
rect 30006 37204 30012 37216
rect 30064 37204 30070 37256
rect 31205 37247 31263 37253
rect 31205 37213 31217 37247
rect 31251 37213 31263 37247
rect 31205 37207 31263 37213
rect 27764 37148 28764 37176
rect 27764 37136 27770 37148
rect 28994 37136 29000 37188
rect 29052 37176 29058 37188
rect 31220 37176 31248 37207
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 32272 37216 32413 37244
rect 32272 37204 32278 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 34514 37204 34520 37256
rect 34572 37244 34578 37256
rect 34977 37247 35035 37253
rect 34977 37244 34989 37247
rect 34572 37216 34989 37244
rect 34572 37204 34578 37216
rect 34977 37213 34989 37216
rect 35023 37213 35035 37247
rect 36170 37244 36176 37256
rect 36131 37216 36176 37244
rect 34977 37207 35035 37213
rect 36170 37204 36176 37216
rect 36228 37204 36234 37256
rect 37737 37247 37795 37253
rect 37737 37213 37749 37247
rect 37783 37244 37795 37247
rect 39666 37244 39672 37256
rect 37783 37216 39672 37244
rect 37783 37213 37795 37216
rect 37737 37207 37795 37213
rect 39666 37204 39672 37216
rect 39724 37204 39730 37256
rect 29052 37148 31248 37176
rect 29052 37136 29058 37148
rect 33134 37136 33140 37188
rect 33192 37136 33198 37188
rect 26605 37111 26663 37117
rect 26605 37108 26617 37111
rect 22152 37080 26617 37108
rect 22152 37068 22158 37080
rect 26605 37077 26617 37080
rect 26651 37077 26663 37111
rect 26605 37071 26663 37077
rect 27341 37111 27399 37117
rect 27341 37077 27353 37111
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 27614 37068 27620 37120
rect 27672 37108 27678 37120
rect 27893 37111 27951 37117
rect 27893 37108 27905 37111
rect 27672 37080 27905 37108
rect 27672 37068 27678 37080
rect 27893 37077 27905 37080
rect 27939 37077 27951 37111
rect 27893 37071 27951 37077
rect 28537 37111 28595 37117
rect 28537 37077 28549 37111
rect 28583 37108 28595 37111
rect 30282 37108 30288 37120
rect 28583 37080 30288 37108
rect 28583 37077 28595 37080
rect 28537 37071 28595 37077
rect 30282 37068 30288 37080
rect 30340 37068 30346 37120
rect 31018 37108 31024 37120
rect 30979 37080 31024 37108
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 34146 37108 34152 37120
rect 34107 37080 34152 37108
rect 34146 37068 34152 37080
rect 34204 37068 34210 37120
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 36136 37080 36369 37108
rect 36136 37068 36142 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3326 36904 3332 36916
rect 1780 36876 3332 36904
rect 1670 36836 1676 36848
rect 1631 36808 1676 36836
rect 1670 36796 1676 36808
rect 1728 36796 1734 36848
rect 1780 36845 1808 36876
rect 3326 36864 3332 36876
rect 3384 36864 3390 36916
rect 3789 36907 3847 36913
rect 3789 36873 3801 36907
rect 3835 36904 3847 36907
rect 5074 36904 5080 36916
rect 3835 36876 5080 36904
rect 3835 36873 3847 36876
rect 3789 36867 3847 36873
rect 5074 36864 5080 36876
rect 5132 36864 5138 36916
rect 5169 36907 5227 36913
rect 5169 36873 5181 36907
rect 5215 36904 5227 36907
rect 8662 36904 8668 36916
rect 5215 36876 8668 36904
rect 5215 36873 5227 36876
rect 5169 36867 5227 36873
rect 8662 36864 8668 36876
rect 8720 36864 8726 36916
rect 9030 36864 9036 36916
rect 9088 36864 9094 36916
rect 9214 36864 9220 36916
rect 9272 36904 9278 36916
rect 11974 36904 11980 36916
rect 9272 36876 11980 36904
rect 9272 36864 9278 36876
rect 11974 36864 11980 36876
rect 12032 36864 12038 36916
rect 12345 36907 12403 36913
rect 12345 36873 12357 36907
rect 12391 36904 12403 36907
rect 13446 36904 13452 36916
rect 12391 36876 13452 36904
rect 12391 36873 12403 36876
rect 12345 36867 12403 36873
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 13538 36864 13544 36916
rect 13596 36904 13602 36916
rect 13817 36907 13875 36913
rect 13817 36904 13829 36907
rect 13596 36876 13829 36904
rect 13596 36864 13602 36876
rect 13817 36873 13829 36876
rect 13863 36873 13875 36907
rect 13817 36867 13875 36873
rect 13906 36864 13912 36916
rect 13964 36904 13970 36916
rect 22002 36904 22008 36916
rect 13964 36876 22008 36904
rect 13964 36864 13970 36876
rect 22002 36864 22008 36876
rect 22060 36864 22066 36916
rect 25866 36904 25872 36916
rect 22756 36876 23704 36904
rect 25827 36876 25872 36904
rect 1765 36839 1823 36845
rect 1765 36805 1777 36839
rect 1811 36805 1823 36839
rect 1765 36799 1823 36805
rect 2314 36796 2320 36848
rect 2372 36836 2378 36848
rect 7098 36836 7104 36848
rect 2372 36808 2774 36836
rect 2372 36796 2378 36808
rect 2746 36768 2774 36808
rect 5368 36808 7104 36836
rect 3329 36771 3387 36777
rect 3329 36768 3341 36771
rect 2746 36740 3341 36768
rect 3329 36737 3341 36740
rect 3375 36737 3387 36771
rect 3329 36731 3387 36737
rect 3418 36728 3424 36780
rect 3476 36768 3482 36780
rect 5368 36777 5396 36808
rect 7098 36796 7104 36808
rect 7156 36796 7162 36848
rect 9048 36836 9076 36864
rect 7852 36808 9076 36836
rect 9125 36839 9183 36845
rect 3973 36771 4031 36777
rect 3973 36768 3985 36771
rect 3476 36740 3985 36768
rect 3476 36728 3482 36740
rect 3973 36737 3985 36740
rect 4019 36737 4031 36771
rect 3973 36731 4031 36737
rect 4709 36771 4767 36777
rect 4709 36737 4721 36771
rect 4755 36737 4767 36771
rect 4709 36731 4767 36737
rect 5353 36771 5411 36777
rect 5353 36737 5365 36771
rect 5399 36737 5411 36771
rect 5353 36731 5411 36737
rect 5997 36771 6055 36777
rect 5997 36737 6009 36771
rect 6043 36737 6055 36771
rect 7006 36768 7012 36780
rect 6967 36740 7012 36768
rect 5997 36731 6055 36737
rect 2682 36700 2688 36712
rect 2643 36672 2688 36700
rect 2682 36660 2688 36672
rect 2740 36660 2746 36712
rect 4724 36700 4752 36731
rect 6012 36700 6040 36731
rect 7006 36728 7012 36740
rect 7064 36728 7070 36780
rect 7852 36777 7880 36808
rect 9125 36805 9137 36839
rect 9171 36836 9183 36839
rect 11146 36836 11152 36848
rect 9171 36808 11152 36836
rect 9171 36805 9183 36808
rect 9125 36799 9183 36805
rect 11146 36796 11152 36808
rect 11204 36796 11210 36848
rect 15286 36796 15292 36848
rect 15344 36836 15350 36848
rect 15381 36839 15439 36845
rect 15381 36836 15393 36839
rect 15344 36808 15393 36836
rect 15344 36796 15350 36808
rect 15381 36805 15393 36808
rect 15427 36805 15439 36839
rect 20070 36836 20076 36848
rect 19642 36808 20076 36836
rect 15381 36799 15439 36805
rect 20070 36796 20076 36808
rect 20128 36796 20134 36848
rect 20162 36796 20168 36848
rect 20220 36836 20226 36848
rect 22756 36836 22784 36876
rect 23569 36839 23627 36845
rect 23569 36836 23581 36839
rect 20220 36808 22784 36836
rect 22940 36808 23581 36836
rect 20220 36796 20226 36808
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36737 7895 36771
rect 7837 36731 7895 36737
rect 8389 36771 8447 36777
rect 8389 36737 8401 36771
rect 8435 36737 8447 36771
rect 9030 36768 9036 36780
rect 8991 36740 9036 36768
rect 8389 36731 8447 36737
rect 8294 36700 8300 36712
rect 4724 36672 5948 36700
rect 6012 36672 8300 36700
rect 4525 36635 4583 36641
rect 4525 36601 4537 36635
rect 4571 36632 4583 36635
rect 5626 36632 5632 36644
rect 4571 36604 5632 36632
rect 4571 36601 4583 36604
rect 4525 36595 4583 36601
rect 5626 36592 5632 36604
rect 5684 36592 5690 36644
rect 3142 36564 3148 36576
rect 3103 36536 3148 36564
rect 3142 36524 3148 36536
rect 3200 36524 3206 36576
rect 5810 36564 5816 36576
rect 5771 36536 5816 36564
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 5920 36564 5948 36672
rect 8294 36660 8300 36672
rect 8352 36660 8358 36712
rect 8404 36700 8432 36731
rect 9030 36728 9036 36740
rect 9088 36728 9094 36780
rect 10226 36728 10232 36780
rect 10284 36768 10290 36780
rect 10505 36771 10563 36777
rect 10505 36768 10517 36771
rect 10284 36740 10517 36768
rect 10284 36728 10290 36740
rect 10505 36737 10517 36740
rect 10551 36737 10563 36771
rect 10505 36731 10563 36737
rect 10870 36728 10876 36780
rect 10928 36768 10934 36780
rect 10965 36771 11023 36777
rect 10965 36768 10977 36771
rect 10928 36740 10977 36768
rect 10928 36728 10934 36740
rect 10965 36737 10977 36740
rect 11011 36737 11023 36771
rect 11885 36771 11943 36777
rect 11885 36768 11897 36771
rect 10965 36731 11023 36737
rect 11072 36740 11897 36768
rect 9677 36703 9735 36709
rect 8404 36672 9628 36700
rect 7101 36635 7159 36641
rect 7101 36601 7113 36635
rect 7147 36632 7159 36635
rect 8570 36632 8576 36644
rect 7147 36604 8432 36632
rect 8531 36604 8576 36632
rect 7147 36601 7159 36604
rect 7101 36595 7159 36601
rect 7466 36564 7472 36576
rect 5920 36536 7472 36564
rect 7466 36524 7472 36536
rect 7524 36524 7530 36576
rect 7650 36564 7656 36576
rect 7611 36536 7656 36564
rect 7650 36524 7656 36536
rect 7708 36524 7714 36576
rect 8404 36564 8432 36604
rect 8570 36592 8576 36604
rect 8628 36592 8634 36644
rect 8846 36564 8852 36576
rect 8404 36536 8852 36564
rect 8846 36524 8852 36536
rect 8904 36524 8910 36576
rect 9600 36564 9628 36672
rect 9677 36669 9689 36703
rect 9723 36669 9735 36703
rect 9677 36663 9735 36669
rect 9692 36632 9720 36663
rect 9766 36660 9772 36712
rect 9824 36700 9830 36712
rect 11072 36700 11100 36740
rect 11885 36737 11897 36740
rect 11931 36737 11943 36771
rect 11885 36731 11943 36737
rect 12989 36771 13047 36777
rect 12989 36737 13001 36771
rect 13035 36737 13047 36771
rect 13630 36768 13636 36780
rect 13591 36740 13636 36768
rect 12989 36731 13047 36737
rect 11698 36700 11704 36712
rect 9824 36672 11100 36700
rect 11659 36672 11704 36700
rect 9824 36660 9830 36672
rect 11698 36660 11704 36672
rect 11756 36660 11762 36712
rect 13004 36700 13032 36731
rect 13630 36728 13636 36740
rect 13688 36728 13694 36780
rect 13722 36728 13728 36780
rect 13780 36768 13786 36780
rect 14369 36771 14427 36777
rect 14369 36768 14381 36771
rect 13780 36740 14381 36768
rect 13780 36728 13786 36740
rect 14369 36737 14381 36740
rect 14415 36737 14427 36771
rect 14369 36731 14427 36737
rect 16853 36771 16911 36777
rect 16853 36737 16865 36771
rect 16899 36768 16911 36771
rect 17862 36768 17868 36780
rect 16899 36740 17868 36768
rect 16899 36737 16911 36740
rect 16853 36731 16911 36737
rect 17862 36728 17868 36740
rect 17920 36728 17926 36780
rect 20990 36728 20996 36780
rect 21048 36768 21054 36780
rect 22738 36768 22744 36780
rect 21048 36740 22744 36768
rect 21048 36728 21054 36740
rect 22738 36728 22744 36740
rect 22796 36728 22802 36780
rect 13906 36700 13912 36712
rect 13004 36672 13912 36700
rect 13906 36660 13912 36672
rect 13964 36660 13970 36712
rect 15289 36703 15347 36709
rect 15289 36669 15301 36703
rect 15335 36700 15347 36703
rect 15378 36700 15384 36712
rect 15335 36672 15384 36700
rect 15335 36669 15347 36672
rect 15289 36663 15347 36669
rect 15378 36660 15384 36672
rect 15436 36660 15442 36712
rect 16298 36700 16304 36712
rect 16211 36672 16304 36700
rect 16298 36660 16304 36672
rect 16356 36700 16362 36712
rect 17129 36703 17187 36709
rect 16356 36672 16988 36700
rect 16356 36660 16362 36672
rect 9692 36604 11192 36632
rect 10134 36564 10140 36576
rect 9600 36536 10140 36564
rect 10134 36524 10140 36536
rect 10192 36524 10198 36576
rect 10318 36564 10324 36576
rect 10279 36536 10324 36564
rect 10318 36524 10324 36536
rect 10376 36524 10382 36576
rect 11054 36564 11060 36576
rect 11015 36536 11060 36564
rect 11054 36524 11060 36536
rect 11112 36524 11118 36576
rect 11164 36564 11192 36604
rect 12434 36592 12440 36644
rect 12492 36632 12498 36644
rect 12492 36604 12940 36632
rect 12492 36592 12498 36604
rect 12526 36564 12532 36576
rect 11164 36536 12532 36564
rect 12526 36524 12532 36536
rect 12584 36524 12590 36576
rect 12618 36524 12624 36576
rect 12676 36564 12682 36576
rect 12805 36567 12863 36573
rect 12805 36564 12817 36567
rect 12676 36536 12817 36564
rect 12676 36524 12682 36536
rect 12805 36533 12817 36536
rect 12851 36533 12863 36567
rect 12912 36564 12940 36604
rect 16666 36592 16672 36644
rect 16724 36632 16730 36644
rect 16850 36632 16856 36644
rect 16724 36604 16856 36632
rect 16724 36592 16730 36604
rect 16850 36592 16856 36604
rect 16908 36592 16914 36644
rect 16960 36632 16988 36672
rect 17129 36669 17141 36703
rect 17175 36700 17187 36703
rect 17678 36700 17684 36712
rect 17175 36672 17684 36700
rect 17175 36669 17187 36672
rect 17129 36663 17187 36669
rect 17678 36660 17684 36672
rect 17736 36660 17742 36712
rect 18138 36700 18144 36712
rect 18099 36672 18144 36700
rect 18138 36660 18144 36672
rect 18196 36660 18202 36712
rect 18414 36700 18420 36712
rect 18375 36672 18420 36700
rect 18414 36660 18420 36672
rect 18472 36700 18478 36712
rect 19426 36700 19432 36712
rect 18472 36672 19432 36700
rect 18472 36660 18478 36672
rect 19426 36660 19432 36672
rect 19484 36660 19490 36712
rect 20346 36700 20352 36712
rect 20307 36672 20352 36700
rect 20346 36660 20352 36672
rect 20404 36660 20410 36712
rect 20438 36660 20444 36712
rect 20496 36700 20502 36712
rect 20625 36703 20683 36709
rect 20625 36700 20637 36703
rect 20496 36672 20637 36700
rect 20496 36660 20502 36672
rect 20625 36669 20637 36672
rect 20671 36669 20683 36703
rect 20625 36663 20683 36669
rect 21358 36660 21364 36712
rect 21416 36700 21422 36712
rect 22940 36700 22968 36808
rect 23569 36805 23581 36808
rect 23615 36805 23627 36839
rect 23676 36836 23704 36876
rect 25866 36864 25872 36876
rect 25924 36864 25930 36916
rect 31018 36904 31024 36916
rect 26528 36876 31024 36904
rect 23676 36808 24058 36836
rect 23569 36799 23627 36805
rect 24854 36728 24860 36780
rect 24912 36768 24918 36780
rect 25777 36771 25835 36777
rect 24912 36740 25728 36768
rect 24912 36728 24918 36740
rect 21416 36672 22968 36700
rect 23293 36703 23351 36709
rect 21416 36660 21422 36672
rect 23293 36669 23305 36703
rect 23339 36700 23351 36703
rect 23339 36672 23428 36700
rect 23339 36669 23351 36672
rect 23293 36663 23351 36669
rect 17218 36632 17224 36644
rect 16960 36604 17224 36632
rect 17218 36592 17224 36604
rect 17276 36592 17282 36644
rect 19702 36592 19708 36644
rect 19760 36632 19766 36644
rect 20714 36632 20720 36644
rect 19760 36604 20720 36632
rect 19760 36592 19766 36604
rect 20714 36592 20720 36604
rect 20772 36592 20778 36644
rect 14369 36567 14427 36573
rect 14369 36564 14381 36567
rect 12912 36536 14381 36564
rect 12805 36527 12863 36533
rect 14369 36533 14381 36536
rect 14415 36533 14427 36567
rect 14369 36527 14427 36533
rect 14826 36524 14832 36576
rect 14884 36564 14890 36576
rect 17770 36564 17776 36576
rect 14884 36536 17776 36564
rect 14884 36524 14890 36536
rect 17770 36524 17776 36536
rect 17828 36524 17834 36576
rect 18230 36524 18236 36576
rect 18288 36564 18294 36576
rect 19889 36567 19947 36573
rect 19889 36564 19901 36567
rect 18288 36536 19901 36564
rect 18288 36524 18294 36536
rect 19889 36533 19901 36536
rect 19935 36564 19947 36567
rect 23290 36564 23296 36576
rect 19935 36536 23296 36564
rect 19935 36533 19947 36536
rect 19889 36527 19947 36533
rect 23290 36524 23296 36536
rect 23348 36524 23354 36576
rect 23400 36564 23428 36672
rect 23934 36660 23940 36712
rect 23992 36700 23998 36712
rect 25317 36703 25375 36709
rect 23992 36672 24624 36700
rect 23992 36660 23998 36672
rect 24596 36632 24624 36672
rect 25317 36669 25329 36703
rect 25363 36700 25375 36703
rect 25406 36700 25412 36712
rect 25363 36672 25412 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 25700 36700 25728 36740
rect 25777 36737 25789 36771
rect 25823 36768 25835 36771
rect 26528 36768 26556 36876
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 32306 36864 32312 36916
rect 32364 36904 32370 36916
rect 32493 36907 32551 36913
rect 32493 36904 32505 36907
rect 32364 36876 32505 36904
rect 32364 36864 32370 36876
rect 32493 36873 32505 36876
rect 32539 36873 32551 36907
rect 32493 36867 32551 36873
rect 32858 36864 32864 36916
rect 32916 36904 32922 36916
rect 33229 36907 33287 36913
rect 33229 36904 33241 36907
rect 32916 36876 33241 36904
rect 32916 36864 32922 36876
rect 33229 36873 33241 36876
rect 33275 36873 33287 36907
rect 36722 36904 36728 36916
rect 33229 36867 33287 36873
rect 34348 36876 36728 36904
rect 27982 36836 27988 36848
rect 27540 36808 27988 36836
rect 25823 36740 26556 36768
rect 26605 36771 26663 36777
rect 25823 36737 25835 36740
rect 25777 36731 25835 36737
rect 26605 36737 26617 36771
rect 26651 36737 26663 36771
rect 26605 36731 26663 36737
rect 26620 36700 26648 36731
rect 25700 36672 26648 36700
rect 26142 36632 26148 36644
rect 24596 36604 26148 36632
rect 26142 36592 26148 36604
rect 26200 36592 26206 36644
rect 26234 36592 26240 36644
rect 26292 36632 26298 36644
rect 27540 36632 27568 36808
rect 27982 36796 27988 36808
rect 28040 36796 28046 36848
rect 30193 36839 30251 36845
rect 30193 36836 30205 36839
rect 29472 36808 30205 36836
rect 28994 36728 29000 36780
rect 29052 36728 29058 36780
rect 27617 36703 27675 36709
rect 27617 36669 27629 36703
rect 27663 36700 27675 36703
rect 27890 36700 27896 36712
rect 27663 36672 27752 36700
rect 27851 36672 27896 36700
rect 27663 36669 27675 36672
rect 27617 36663 27675 36669
rect 26292 36604 27568 36632
rect 26292 36592 26298 36604
rect 27724 36576 27752 36672
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 27982 36660 27988 36712
rect 28040 36700 28046 36712
rect 29472 36700 29500 36808
rect 30193 36805 30205 36808
rect 30239 36805 30251 36839
rect 33870 36836 33876 36848
rect 30193 36799 30251 36805
rect 31726 36808 33876 36836
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 30101 36771 30159 36777
rect 30101 36768 30113 36771
rect 29604 36740 30113 36768
rect 29604 36728 29610 36740
rect 30101 36737 30113 36740
rect 30147 36737 30159 36771
rect 30101 36731 30159 36737
rect 28040 36672 29500 36700
rect 29641 36703 29699 36709
rect 28040 36660 28046 36672
rect 29641 36669 29653 36703
rect 29687 36669 29699 36703
rect 30116 36700 30144 36731
rect 30282 36728 30288 36780
rect 30340 36768 30346 36780
rect 31113 36771 31171 36777
rect 31113 36768 31125 36771
rect 30340 36740 31125 36768
rect 30340 36728 30346 36740
rect 31113 36737 31125 36740
rect 31159 36737 31171 36771
rect 31113 36731 31171 36737
rect 31573 36771 31631 36777
rect 31573 36737 31585 36771
rect 31619 36768 31631 36771
rect 31726 36768 31754 36808
rect 33870 36796 33876 36808
rect 33928 36796 33934 36848
rect 32306 36768 32312 36780
rect 31619 36740 31754 36768
rect 32267 36740 32312 36768
rect 31619 36737 31631 36740
rect 31573 36731 31631 36737
rect 31588 36700 31616 36731
rect 32306 36728 32312 36740
rect 32364 36728 32370 36780
rect 33042 36768 33048 36780
rect 33003 36740 33048 36768
rect 33042 36728 33048 36740
rect 33100 36728 33106 36780
rect 33965 36771 34023 36777
rect 33965 36737 33977 36771
rect 34011 36768 34023 36771
rect 34348 36768 34376 36876
rect 36722 36864 36728 36876
rect 36780 36864 36786 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37645 36907 37703 36913
rect 37645 36904 37657 36907
rect 37424 36876 37657 36904
rect 37424 36864 37430 36876
rect 37645 36873 37657 36876
rect 37691 36873 37703 36907
rect 37645 36867 37703 36873
rect 35710 36796 35716 36848
rect 35768 36796 35774 36848
rect 34011 36740 34376 36768
rect 36725 36771 36783 36777
rect 34011 36737 34023 36740
rect 33965 36731 34023 36737
rect 36725 36737 36737 36771
rect 36771 36737 36783 36771
rect 36725 36731 36783 36737
rect 37461 36771 37519 36777
rect 37461 36737 37473 36771
rect 37507 36737 37519 36771
rect 37461 36731 37519 36737
rect 30116 36672 31616 36700
rect 29641 36663 29699 36669
rect 23566 36564 23572 36576
rect 23400 36536 23572 36564
rect 23566 36524 23572 36536
rect 23624 36564 23630 36576
rect 24762 36564 24768 36576
rect 23624 36536 24768 36564
rect 23624 36524 23630 36536
rect 24762 36524 24768 36536
rect 24820 36524 24826 36576
rect 26418 36564 26424 36576
rect 26379 36536 26424 36564
rect 26418 36524 26424 36536
rect 26476 36524 26482 36576
rect 27706 36524 27712 36576
rect 27764 36524 27770 36576
rect 27890 36524 27896 36576
rect 27948 36564 27954 36576
rect 29656 36564 29684 36663
rect 32214 36660 32220 36712
rect 32272 36700 32278 36712
rect 34422 36700 34428 36712
rect 32272 36672 34428 36700
rect 32272 36660 32278 36672
rect 34422 36660 34428 36672
rect 34480 36660 34486 36712
rect 34698 36700 34704 36712
rect 34659 36672 34704 36700
rect 34698 36660 34704 36672
rect 34756 36660 34762 36712
rect 36740 36700 36768 36731
rect 35866 36672 36768 36700
rect 35866 36644 35894 36672
rect 30929 36635 30987 36641
rect 30929 36601 30941 36635
rect 30975 36632 30987 36635
rect 30975 36604 33916 36632
rect 30975 36601 30987 36604
rect 30929 36595 30987 36601
rect 31662 36564 31668 36576
rect 27948 36536 29684 36564
rect 31623 36536 31668 36564
rect 27948 36524 27954 36536
rect 31662 36524 31668 36536
rect 31720 36524 31726 36576
rect 33778 36564 33784 36576
rect 33739 36536 33784 36564
rect 33778 36524 33784 36536
rect 33836 36524 33842 36576
rect 33888 36564 33916 36604
rect 35802 36592 35808 36644
rect 35860 36604 35894 36644
rect 37476 36632 37504 36731
rect 36004 36604 37504 36632
rect 35860 36592 35866 36604
rect 36004 36564 36032 36604
rect 33888 36536 36032 36564
rect 36170 36524 36176 36576
rect 36228 36564 36234 36576
rect 36814 36564 36820 36576
rect 36228 36536 36273 36564
rect 36775 36536 36820 36564
rect 36228 36524 36234 36536
rect 36814 36524 36820 36536
rect 36872 36524 36878 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 3786 36320 3792 36372
rect 3844 36360 3850 36372
rect 7101 36363 7159 36369
rect 7101 36360 7113 36363
rect 3844 36332 7113 36360
rect 3844 36320 3850 36332
rect 7101 36329 7113 36332
rect 7147 36329 7159 36363
rect 7101 36323 7159 36329
rect 8481 36363 8539 36369
rect 8481 36329 8493 36363
rect 8527 36360 8539 36363
rect 11698 36360 11704 36372
rect 8527 36332 11704 36360
rect 8527 36329 8539 36332
rect 8481 36323 8539 36329
rect 11698 36320 11704 36332
rect 11756 36320 11762 36372
rect 11882 36320 11888 36372
rect 11940 36360 11946 36372
rect 20438 36360 20444 36372
rect 11940 36332 20444 36360
rect 11940 36320 11946 36332
rect 20438 36320 20444 36332
rect 20496 36320 20502 36372
rect 20714 36320 20720 36372
rect 20772 36360 20778 36372
rect 26418 36360 26424 36372
rect 20772 36332 26424 36360
rect 20772 36320 20778 36332
rect 26418 36320 26424 36332
rect 26476 36320 26482 36372
rect 27614 36320 27620 36372
rect 27672 36360 27678 36372
rect 28997 36363 29055 36369
rect 27672 36332 28304 36360
rect 27672 36320 27678 36332
rect 7837 36295 7895 36301
rect 7837 36261 7849 36295
rect 7883 36292 7895 36295
rect 9766 36292 9772 36304
rect 7883 36264 9772 36292
rect 7883 36261 7895 36264
rect 7837 36255 7895 36261
rect 9766 36252 9772 36264
rect 9824 36252 9830 36304
rect 10134 36292 10140 36304
rect 10095 36264 10140 36292
rect 10134 36252 10140 36264
rect 10192 36252 10198 36304
rect 10318 36252 10324 36304
rect 10376 36292 10382 36304
rect 14826 36292 14832 36304
rect 10376 36264 14832 36292
rect 10376 36252 10382 36264
rect 14826 36252 14832 36264
rect 14884 36252 14890 36304
rect 14921 36295 14979 36301
rect 14921 36261 14933 36295
rect 14967 36292 14979 36295
rect 26326 36292 26332 36304
rect 14967 36264 19564 36292
rect 26287 36264 26332 36292
rect 14967 36261 14979 36264
rect 14921 36255 14979 36261
rect 2682 36224 2688 36236
rect 2643 36196 2688 36224
rect 2682 36184 2688 36196
rect 2740 36224 2746 36236
rect 3418 36224 3424 36236
rect 2740 36196 3424 36224
rect 2740 36184 2746 36196
rect 3418 36184 3424 36196
rect 3476 36184 3482 36236
rect 7006 36224 7012 36236
rect 6012 36196 7012 36224
rect 1762 36156 1768 36168
rect 1723 36128 1768 36156
rect 1762 36116 1768 36128
rect 1820 36116 1826 36168
rect 4157 36159 4215 36165
rect 4157 36125 4169 36159
rect 4203 36156 4215 36159
rect 4614 36156 4620 36168
rect 4203 36128 4620 36156
rect 4203 36125 4215 36128
rect 4157 36119 4215 36125
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 6012 36165 6040 36196
rect 7006 36184 7012 36196
rect 7064 36184 7070 36236
rect 7466 36184 7472 36236
rect 7524 36224 7530 36236
rect 8294 36224 8300 36236
rect 7524 36196 8300 36224
rect 7524 36184 7530 36196
rect 8294 36184 8300 36196
rect 8352 36184 8358 36236
rect 10502 36224 10508 36236
rect 8404 36196 10508 36224
rect 5997 36159 6055 36165
rect 5997 36125 6009 36159
rect 6043 36125 6055 36159
rect 6454 36156 6460 36168
rect 6415 36128 6460 36156
rect 5997 36119 6055 36125
rect 6454 36116 6460 36128
rect 6512 36116 6518 36168
rect 7285 36159 7343 36165
rect 7285 36125 7297 36159
rect 7331 36156 7343 36159
rect 7558 36156 7564 36168
rect 7331 36128 7564 36156
rect 7331 36125 7343 36128
rect 7285 36119 7343 36125
rect 7558 36116 7564 36128
rect 7616 36116 7622 36168
rect 7742 36156 7748 36168
rect 7703 36128 7748 36156
rect 7742 36116 7748 36128
rect 7800 36116 7806 36168
rect 8404 36165 8432 36196
rect 10502 36184 10508 36196
rect 10560 36184 10566 36236
rect 10781 36227 10839 36233
rect 10781 36224 10793 36227
rect 10612 36196 10793 36224
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36125 8447 36159
rect 9306 36156 9312 36168
rect 9267 36128 9312 36156
rect 8389 36119 8447 36125
rect 9306 36116 9312 36128
rect 9364 36116 9370 36168
rect 10042 36156 10048 36168
rect 9955 36128 10048 36156
rect 10042 36116 10048 36128
rect 10100 36156 10106 36168
rect 10318 36156 10324 36168
rect 10100 36128 10324 36156
rect 10100 36116 10106 36128
rect 10318 36116 10324 36128
rect 10376 36116 10382 36168
rect 10410 36116 10416 36168
rect 10468 36156 10474 36168
rect 10612 36156 10640 36196
rect 10781 36193 10793 36196
rect 10827 36193 10839 36227
rect 10781 36187 10839 36193
rect 12526 36184 12532 36236
rect 12584 36224 12590 36236
rect 12805 36227 12863 36233
rect 12805 36224 12817 36227
rect 12584 36196 12817 36224
rect 12584 36184 12590 36196
rect 12805 36193 12817 36196
rect 12851 36193 12863 36227
rect 13446 36224 13452 36236
rect 13407 36196 13452 36224
rect 12805 36187 12863 36193
rect 13446 36184 13452 36196
rect 13504 36224 13510 36236
rect 15565 36227 15623 36233
rect 15565 36224 15577 36227
rect 13504 36196 15577 36224
rect 13504 36184 13510 36196
rect 15565 36193 15577 36196
rect 15611 36193 15623 36227
rect 15565 36187 15623 36193
rect 16761 36227 16819 36233
rect 16761 36193 16773 36227
rect 16807 36224 16819 36227
rect 16942 36224 16948 36236
rect 16807 36196 16948 36224
rect 16807 36193 16819 36196
rect 16761 36187 16819 36193
rect 16942 36184 16948 36196
rect 17000 36184 17006 36236
rect 17126 36184 17132 36236
rect 17184 36224 17190 36236
rect 19334 36224 19340 36236
rect 17184 36196 19340 36224
rect 17184 36184 17190 36196
rect 19334 36184 19340 36196
rect 19392 36184 19398 36236
rect 19536 36224 19564 36264
rect 26326 36252 26332 36264
rect 26384 36252 26390 36304
rect 20162 36224 20168 36236
rect 19536 36196 20168 36224
rect 20162 36184 20168 36196
rect 20220 36184 20226 36236
rect 21729 36227 21787 36233
rect 21729 36193 21741 36227
rect 21775 36224 21787 36227
rect 23566 36224 23572 36236
rect 21775 36196 23572 36224
rect 21775 36193 21787 36196
rect 21729 36187 21787 36193
rect 23566 36184 23572 36196
rect 23624 36184 23630 36236
rect 26789 36227 26847 36233
rect 26789 36193 26801 36227
rect 26835 36224 26847 36227
rect 27706 36224 27712 36236
rect 26835 36196 27712 36224
rect 26835 36193 26847 36196
rect 26789 36187 26847 36193
rect 27706 36184 27712 36196
rect 27764 36184 27770 36236
rect 10468 36128 10640 36156
rect 12989 36159 13047 36165
rect 10468 36116 10474 36128
rect 12989 36125 13001 36159
rect 13035 36125 13047 36159
rect 14826 36156 14832 36168
rect 14787 36128 14832 36156
rect 12989 36119 13047 36125
rect 2406 36088 2412 36100
rect 2367 36060 2412 36088
rect 2406 36048 2412 36060
rect 2464 36048 2470 36100
rect 2498 36048 2504 36100
rect 2556 36088 2562 36100
rect 9214 36088 9220 36100
rect 2556 36060 2601 36088
rect 5828 36060 9220 36088
rect 2556 36048 2562 36060
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 3878 36020 3884 36032
rect 1627 35992 3884 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 3878 35980 3884 35992
rect 3936 35980 3942 36032
rect 3973 36023 4031 36029
rect 3973 35989 3985 36023
rect 4019 36020 4031 36023
rect 5718 36020 5724 36032
rect 4019 35992 5724 36020
rect 4019 35989 4031 35992
rect 3973 35983 4031 35989
rect 5718 35980 5724 35992
rect 5776 35980 5782 36032
rect 5828 36029 5856 36060
rect 9214 36048 9220 36060
rect 9272 36048 9278 36100
rect 9401 36091 9459 36097
rect 9401 36057 9413 36091
rect 9447 36088 9459 36091
rect 10594 36088 10600 36100
rect 9447 36060 10600 36088
rect 9447 36057 9459 36060
rect 9401 36051 9459 36057
rect 10594 36048 10600 36060
rect 10652 36048 10658 36100
rect 10873 36091 10931 36097
rect 10873 36057 10885 36091
rect 10919 36088 10931 36091
rect 10962 36088 10968 36100
rect 10919 36060 10968 36088
rect 10919 36057 10931 36060
rect 10873 36051 10931 36057
rect 10962 36048 10968 36060
rect 11020 36048 11026 36100
rect 11698 36048 11704 36100
rect 11756 36088 11762 36100
rect 11793 36091 11851 36097
rect 11793 36088 11805 36091
rect 11756 36060 11805 36088
rect 11756 36048 11762 36060
rect 11793 36057 11805 36060
rect 11839 36088 11851 36091
rect 12066 36088 12072 36100
rect 11839 36060 12072 36088
rect 11839 36057 11851 36060
rect 11793 36051 11851 36057
rect 12066 36048 12072 36060
rect 12124 36048 12130 36100
rect 12158 36048 12164 36100
rect 12216 36088 12222 36100
rect 13004 36088 13032 36119
rect 14826 36116 14832 36128
rect 14884 36116 14890 36168
rect 18230 36156 18236 36168
rect 17604 36128 17908 36156
rect 18191 36128 18236 36156
rect 12216 36060 13032 36088
rect 12216 36048 12222 36060
rect 15654 36048 15660 36100
rect 15712 36088 15718 36100
rect 16206 36088 16212 36100
rect 15712 36060 15757 36088
rect 16167 36060 16212 36088
rect 15712 36048 15718 36060
rect 16206 36048 16212 36060
rect 16264 36048 16270 36100
rect 16298 36048 16304 36100
rect 16356 36088 16362 36100
rect 16853 36091 16911 36097
rect 16853 36088 16865 36091
rect 16356 36060 16865 36088
rect 16356 36048 16362 36060
rect 16853 36057 16865 36060
rect 16899 36057 16911 36091
rect 17604 36088 17632 36128
rect 17770 36088 17776 36100
rect 16853 36051 16911 36057
rect 16960 36060 17632 36088
rect 17731 36060 17776 36088
rect 5813 36023 5871 36029
rect 5813 35989 5825 36023
rect 5859 35989 5871 36023
rect 5813 35983 5871 35989
rect 6549 36023 6607 36029
rect 6549 35989 6561 36023
rect 6595 36020 6607 36023
rect 7466 36020 7472 36032
rect 6595 35992 7472 36020
rect 6595 35989 6607 35992
rect 6549 35983 6607 35989
rect 7466 35980 7472 35992
rect 7524 35980 7530 36032
rect 7834 35980 7840 36032
rect 7892 36020 7898 36032
rect 10410 36020 10416 36032
rect 7892 35992 10416 36020
rect 7892 35980 7898 35992
rect 10410 35980 10416 35992
rect 10468 35980 10474 36032
rect 15286 35980 15292 36032
rect 15344 36020 15350 36032
rect 16960 36020 16988 36060
rect 17770 36048 17776 36060
rect 17828 36048 17834 36100
rect 17880 36088 17908 36128
rect 18230 36116 18236 36128
rect 18288 36116 18294 36168
rect 19242 36116 19248 36168
rect 19300 36156 19306 36168
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 19300 36128 19441 36156
rect 19300 36116 19306 36128
rect 19429 36125 19441 36128
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 28276 36156 28304 36332
rect 28997 36329 29009 36363
rect 29043 36360 29055 36363
rect 33042 36360 33048 36372
rect 29043 36332 33048 36360
rect 29043 36329 29055 36332
rect 28997 36323 29055 36329
rect 33042 36320 33048 36332
rect 33100 36320 33106 36372
rect 33778 36320 33784 36372
rect 33836 36360 33842 36372
rect 37918 36360 37924 36372
rect 33836 36332 37924 36360
rect 33836 36320 33842 36332
rect 37918 36320 37924 36332
rect 37976 36320 37982 36372
rect 28442 36252 28448 36304
rect 28500 36292 28506 36304
rect 29546 36292 29552 36304
rect 28500 36264 29552 36292
rect 28500 36252 28506 36264
rect 29546 36252 29552 36264
rect 29604 36252 29610 36304
rect 33870 36252 33876 36304
rect 33928 36292 33934 36304
rect 37550 36292 37556 36304
rect 33928 36264 35020 36292
rect 37511 36264 37556 36292
rect 33928 36252 33934 36264
rect 29733 36227 29791 36233
rect 29733 36193 29745 36227
rect 29779 36224 29791 36227
rect 32214 36224 32220 36236
rect 29779 36196 32220 36224
rect 29779 36193 29791 36196
rect 29733 36187 29791 36193
rect 32214 36184 32220 36196
rect 32272 36184 32278 36236
rect 34422 36184 34428 36236
rect 34480 36224 34486 36236
rect 34885 36227 34943 36233
rect 34885 36224 34897 36227
rect 34480 36196 34897 36224
rect 34480 36184 34486 36196
rect 34885 36193 34897 36196
rect 34931 36193 34943 36227
rect 34992 36224 35020 36264
rect 37550 36252 37556 36264
rect 37608 36252 37614 36304
rect 35802 36224 35808 36236
rect 34992 36196 35808 36224
rect 34885 36187 34943 36193
rect 35802 36184 35808 36196
rect 35860 36184 35866 36236
rect 29181 36159 29239 36165
rect 29181 36156 29193 36159
rect 28276 36128 29193 36156
rect 24581 36119 24639 36125
rect 29181 36125 29193 36128
rect 29227 36125 29239 36159
rect 29181 36119 29239 36125
rect 19610 36088 19616 36100
rect 17880 36060 19616 36088
rect 19610 36048 19616 36060
rect 19668 36048 19674 36100
rect 19705 36091 19763 36097
rect 19705 36057 19717 36091
rect 19751 36057 19763 36091
rect 19705 36051 19763 36057
rect 15344 35992 16988 36020
rect 15344 35980 15350 35992
rect 17034 35980 17040 36032
rect 17092 36020 17098 36032
rect 18325 36023 18383 36029
rect 18325 36020 18337 36023
rect 17092 35992 18337 36020
rect 17092 35980 17098 35992
rect 18325 35989 18337 35992
rect 18371 35989 18383 36023
rect 19720 36020 19748 36051
rect 20714 36048 20720 36100
rect 20772 36048 20778 36100
rect 21008 36060 21312 36088
rect 20530 36020 20536 36032
rect 19720 35992 20536 36020
rect 18325 35983 18383 35989
rect 20530 35980 20536 35992
rect 20588 35980 20594 36032
rect 20622 35980 20628 36032
rect 20680 36020 20686 36032
rect 21008 36020 21036 36060
rect 21174 36020 21180 36032
rect 20680 35992 21036 36020
rect 21135 35992 21180 36020
rect 20680 35980 20686 35992
rect 21174 35980 21180 35992
rect 21232 35980 21238 36032
rect 21284 36020 21312 36060
rect 21910 36048 21916 36100
rect 21968 36088 21974 36100
rect 22005 36091 22063 36097
rect 22005 36088 22017 36091
rect 21968 36060 22017 36088
rect 21968 36048 21974 36060
rect 22005 36057 22017 36060
rect 22051 36057 22063 36091
rect 22005 36051 22063 36057
rect 22296 36060 22494 36088
rect 22296 36020 22324 36060
rect 23290 36048 23296 36100
rect 23348 36088 23354 36100
rect 24596 36088 24624 36119
rect 37182 36116 37188 36168
rect 37240 36156 37246 36168
rect 37369 36159 37427 36165
rect 37369 36156 37381 36159
rect 37240 36128 37381 36156
rect 37240 36116 37246 36128
rect 37369 36125 37381 36128
rect 37415 36125 37427 36159
rect 38010 36156 38016 36168
rect 37971 36128 38016 36156
rect 37369 36119 37427 36125
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 24762 36088 24768 36100
rect 23348 36060 23612 36088
rect 24596 36060 24768 36088
rect 23348 36048 23354 36060
rect 23474 36020 23480 36032
rect 21284 35992 22324 36020
rect 23435 35992 23480 36020
rect 23474 35980 23480 35992
rect 23532 35980 23538 36032
rect 23584 36020 23612 36060
rect 24762 36048 24768 36060
rect 24820 36048 24826 36100
rect 24854 36048 24860 36100
rect 24912 36088 24918 36100
rect 24912 36060 25268 36088
rect 24912 36048 24918 36060
rect 24946 36020 24952 36032
rect 23584 35992 24952 36020
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 25240 36020 25268 36060
rect 25314 36048 25320 36100
rect 25372 36048 25378 36100
rect 26142 36048 26148 36100
rect 26200 36088 26206 36100
rect 27065 36091 27123 36097
rect 27065 36088 27077 36091
rect 26200 36060 27077 36088
rect 26200 36048 26206 36060
rect 27065 36057 27077 36060
rect 27111 36057 27123 36091
rect 27065 36051 27123 36057
rect 27798 36048 27804 36100
rect 27856 36048 27862 36100
rect 28350 36048 28356 36100
rect 28408 36088 28414 36100
rect 28408 36060 29868 36088
rect 28408 36048 28414 36060
rect 27890 36020 27896 36032
rect 25240 35992 27896 36020
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 28074 35980 28080 36032
rect 28132 36020 28138 36032
rect 28537 36023 28595 36029
rect 28537 36020 28549 36023
rect 28132 35992 28549 36020
rect 28132 35980 28138 35992
rect 28537 35989 28549 35992
rect 28583 35989 28595 36023
rect 29840 36020 29868 36060
rect 29914 36048 29920 36100
rect 29972 36088 29978 36100
rect 30009 36091 30067 36097
rect 30009 36088 30021 36091
rect 29972 36060 30021 36088
rect 29972 36048 29978 36060
rect 30009 36057 30021 36060
rect 30055 36057 30067 36091
rect 30009 36051 30067 36057
rect 30466 36048 30472 36100
rect 30524 36048 30530 36100
rect 31754 36088 31760 36100
rect 31312 36060 31760 36088
rect 31312 36020 31340 36060
rect 31754 36048 31760 36060
rect 31812 36048 31818 36100
rect 32493 36091 32551 36097
rect 32493 36057 32505 36091
rect 32539 36057 32551 36091
rect 34514 36088 34520 36100
rect 33718 36060 34520 36088
rect 32493 36051 32551 36057
rect 29840 35992 31340 36020
rect 28537 35983 28595 35989
rect 31386 35980 31392 36032
rect 31444 36020 31450 36032
rect 32508 36020 32536 36051
rect 34514 36048 34520 36060
rect 34572 36048 34578 36100
rect 34606 36048 34612 36100
rect 34664 36088 34670 36100
rect 35161 36091 35219 36097
rect 35161 36088 35173 36091
rect 34664 36060 35173 36088
rect 34664 36048 34670 36060
rect 35161 36057 35173 36060
rect 35207 36057 35219 36091
rect 36814 36088 36820 36100
rect 36386 36060 36820 36088
rect 35161 36051 35219 36057
rect 33962 36020 33968 36032
rect 31444 35992 32536 36020
rect 33923 35992 33968 36020
rect 31444 35980 31450 35992
rect 33962 35980 33968 35992
rect 34020 35980 34026 36032
rect 35176 36020 35204 36051
rect 36814 36048 36820 36060
rect 36872 36048 36878 36100
rect 35894 36020 35900 36032
rect 35176 35992 35900 36020
rect 35894 35980 35900 35992
rect 35952 35980 35958 36032
rect 35986 35980 35992 36032
rect 36044 36020 36050 36032
rect 36633 36023 36691 36029
rect 36633 36020 36645 36023
rect 36044 35992 36645 36020
rect 36044 35980 36050 35992
rect 36633 35989 36645 35992
rect 36679 35989 36691 36023
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 36633 35983 36691 35989
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 3326 35816 3332 35828
rect 3287 35788 3332 35816
rect 3326 35776 3332 35788
rect 3384 35776 3390 35828
rect 12986 35816 12992 35828
rect 9784 35788 12992 35816
rect 1670 35748 1676 35760
rect 1631 35720 1676 35748
rect 1670 35708 1676 35720
rect 1728 35708 1734 35760
rect 1762 35708 1768 35760
rect 1820 35748 1826 35760
rect 2682 35748 2688 35760
rect 1820 35720 1865 35748
rect 2643 35720 2688 35748
rect 1820 35708 1826 35720
rect 2682 35708 2688 35720
rect 2740 35708 2746 35760
rect 7837 35751 7895 35757
rect 7837 35717 7849 35751
rect 7883 35748 7895 35751
rect 8570 35748 8576 35760
rect 7883 35720 8576 35748
rect 7883 35717 7895 35720
rect 7837 35711 7895 35717
rect 8570 35708 8576 35720
rect 8628 35708 8634 35760
rect 3234 35680 3240 35692
rect 3195 35652 3240 35680
rect 3234 35640 3240 35652
rect 3292 35640 3298 35692
rect 9784 35689 9812 35788
rect 12986 35776 12992 35788
rect 13044 35776 13050 35828
rect 13081 35819 13139 35825
rect 13081 35785 13093 35819
rect 13127 35816 13139 35819
rect 13446 35816 13452 35828
rect 13127 35788 13452 35816
rect 13127 35785 13139 35788
rect 13081 35779 13139 35785
rect 13446 35776 13452 35788
rect 13504 35776 13510 35828
rect 13538 35776 13544 35828
rect 13596 35816 13602 35828
rect 13596 35788 15424 35816
rect 13596 35776 13602 35788
rect 10318 35708 10324 35760
rect 10376 35748 10382 35760
rect 10597 35751 10655 35757
rect 10597 35748 10609 35751
rect 10376 35720 10609 35748
rect 10376 35708 10382 35720
rect 10597 35717 10609 35720
rect 10643 35717 10655 35751
rect 10597 35711 10655 35717
rect 11606 35708 11612 35760
rect 11664 35748 11670 35760
rect 15286 35748 15292 35760
rect 11664 35720 15292 35748
rect 11664 35708 11670 35720
rect 15286 35708 15292 35720
rect 15344 35708 15350 35760
rect 9769 35683 9827 35689
rect 9769 35649 9781 35683
rect 9815 35649 9827 35683
rect 9769 35643 9827 35649
rect 11238 35640 11244 35692
rect 11296 35680 11302 35692
rect 11793 35683 11851 35689
rect 11793 35680 11805 35683
rect 11296 35652 11805 35680
rect 11296 35640 11302 35652
rect 11793 35649 11805 35652
rect 11839 35680 11851 35683
rect 12066 35680 12072 35692
rect 11839 35652 12072 35680
rect 11839 35649 11851 35652
rect 11793 35643 11851 35649
rect 12066 35640 12072 35652
rect 12124 35640 12130 35692
rect 12434 35680 12440 35692
rect 12395 35652 12440 35680
rect 12434 35640 12440 35652
rect 12492 35640 12498 35692
rect 13814 35640 13820 35692
rect 13872 35680 13878 35692
rect 14093 35683 14151 35689
rect 14093 35680 14105 35683
rect 13872 35652 14105 35680
rect 13872 35640 13878 35652
rect 14093 35649 14105 35652
rect 14139 35680 14151 35683
rect 14737 35683 14795 35689
rect 14737 35680 14749 35683
rect 14139 35652 14749 35680
rect 14139 35649 14151 35652
rect 14093 35643 14151 35649
rect 14737 35649 14749 35652
rect 14783 35680 14795 35683
rect 14826 35680 14832 35692
rect 14783 35652 14832 35680
rect 14783 35649 14795 35652
rect 14737 35643 14795 35649
rect 14826 35640 14832 35652
rect 14884 35640 14890 35692
rect 15396 35689 15424 35788
rect 16206 35776 16212 35828
rect 16264 35816 16270 35828
rect 16264 35788 17632 35816
rect 16264 35776 16270 35788
rect 17034 35748 17040 35760
rect 16995 35720 17040 35748
rect 17034 35708 17040 35720
rect 17092 35708 17098 35760
rect 17604 35757 17632 35788
rect 17770 35776 17776 35828
rect 17828 35816 17834 35828
rect 27522 35816 27528 35828
rect 17828 35788 27528 35816
rect 17828 35776 17834 35788
rect 27522 35776 27528 35788
rect 27580 35776 27586 35828
rect 33962 35816 33968 35828
rect 28276 35788 33968 35816
rect 17589 35751 17647 35757
rect 17589 35717 17601 35751
rect 17635 35717 17647 35751
rect 17589 35711 17647 35717
rect 18417 35751 18475 35757
rect 18417 35717 18429 35751
rect 18463 35748 18475 35751
rect 18506 35748 18512 35760
rect 18463 35720 18512 35748
rect 18463 35717 18475 35720
rect 18417 35711 18475 35717
rect 18506 35708 18512 35720
rect 18564 35708 18570 35760
rect 19426 35708 19432 35760
rect 19484 35708 19490 35760
rect 28276 35757 28304 35788
rect 33962 35776 33968 35788
rect 34020 35816 34026 35828
rect 34330 35816 34336 35828
rect 34020 35788 34336 35816
rect 34020 35776 34026 35788
rect 34330 35776 34336 35788
rect 34388 35776 34394 35828
rect 35621 35819 35679 35825
rect 35621 35785 35633 35819
rect 35667 35816 35679 35819
rect 35710 35816 35716 35828
rect 35667 35788 35716 35816
rect 35667 35785 35679 35788
rect 35621 35779 35679 35785
rect 35710 35776 35716 35788
rect 35768 35776 35774 35828
rect 36722 35776 36728 35828
rect 36780 35816 36786 35828
rect 36817 35819 36875 35825
rect 36817 35816 36829 35819
rect 36780 35788 36829 35816
rect 36780 35776 36786 35788
rect 36817 35785 36829 35788
rect 36863 35785 36875 35819
rect 36817 35779 36875 35785
rect 28261 35751 28319 35757
rect 19720 35720 25622 35748
rect 15381 35683 15439 35689
rect 15381 35649 15393 35683
rect 15427 35649 15439 35683
rect 15381 35643 15439 35649
rect 16301 35683 16359 35689
rect 16301 35649 16313 35683
rect 16347 35680 16359 35683
rect 16758 35680 16764 35692
rect 16347 35652 16764 35680
rect 16347 35649 16359 35652
rect 16301 35643 16359 35649
rect 16758 35640 16764 35652
rect 16816 35640 16822 35692
rect 18138 35680 18144 35692
rect 18099 35652 18144 35680
rect 18138 35640 18144 35652
rect 18196 35640 18202 35692
rect 7009 35615 7067 35621
rect 7009 35581 7021 35615
rect 7055 35612 7067 35615
rect 7745 35615 7803 35621
rect 7745 35612 7757 35615
rect 7055 35584 7757 35612
rect 7055 35581 7067 35584
rect 7009 35575 7067 35581
rect 7745 35581 7757 35584
rect 7791 35581 7803 35615
rect 7745 35575 7803 35581
rect 8757 35615 8815 35621
rect 8757 35581 8769 35615
rect 8803 35581 8815 35615
rect 8757 35575 8815 35581
rect 8772 35476 8800 35575
rect 8846 35572 8852 35624
rect 8904 35612 8910 35624
rect 10505 35615 10563 35621
rect 10505 35612 10517 35615
rect 8904 35584 10517 35612
rect 8904 35572 8910 35584
rect 10505 35581 10517 35584
rect 10551 35581 10563 35615
rect 10505 35575 10563 35581
rect 11146 35572 11152 35624
rect 11204 35612 11210 35624
rect 12621 35615 12679 35621
rect 12621 35612 12633 35615
rect 11204 35584 12633 35612
rect 11204 35572 11210 35584
rect 12621 35581 12633 35584
rect 12667 35581 12679 35615
rect 13906 35612 13912 35624
rect 12621 35575 12679 35581
rect 12728 35584 13912 35612
rect 9861 35547 9919 35553
rect 9861 35513 9873 35547
rect 9907 35544 9919 35547
rect 10962 35544 10968 35556
rect 9907 35516 10968 35544
rect 9907 35513 9919 35516
rect 9861 35507 9919 35513
rect 10962 35504 10968 35516
rect 11020 35504 11026 35556
rect 11057 35547 11115 35553
rect 11057 35513 11069 35547
rect 11103 35544 11115 35547
rect 11238 35544 11244 35556
rect 11103 35516 11244 35544
rect 11103 35513 11115 35516
rect 11057 35507 11115 35513
rect 11238 35504 11244 35516
rect 11296 35544 11302 35556
rect 12728 35544 12756 35584
rect 13906 35572 13912 35584
rect 13964 35572 13970 35624
rect 14185 35615 14243 35621
rect 14185 35581 14197 35615
rect 14231 35612 14243 35615
rect 16666 35612 16672 35624
rect 14231 35584 16672 35612
rect 14231 35581 14243 35584
rect 14185 35575 14243 35581
rect 16666 35572 16672 35584
rect 16724 35572 16730 35624
rect 16945 35615 17003 35621
rect 16945 35581 16957 35615
rect 16991 35612 17003 35615
rect 17770 35612 17776 35624
rect 16991 35584 17776 35612
rect 16991 35581 17003 35584
rect 16945 35575 17003 35581
rect 17770 35572 17776 35584
rect 17828 35572 17834 35624
rect 19720 35612 19748 35720
rect 28261 35717 28273 35751
rect 28307 35717 28319 35751
rect 28261 35711 28319 35717
rect 31386 35708 31392 35760
rect 31444 35748 31450 35760
rect 34698 35748 34704 35760
rect 31444 35720 34704 35748
rect 31444 35708 31450 35720
rect 34698 35708 34704 35720
rect 34756 35708 34762 35760
rect 20254 35640 20260 35692
rect 20312 35680 20318 35692
rect 24670 35680 24676 35692
rect 20312 35652 24676 35680
rect 20312 35640 20318 35652
rect 24670 35640 24676 35652
rect 24728 35640 24734 35692
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35680 27399 35683
rect 27614 35680 27620 35692
rect 27387 35652 27620 35680
rect 27387 35649 27399 35652
rect 27341 35643 27399 35649
rect 27614 35640 27620 35652
rect 27672 35640 27678 35692
rect 30282 35680 30288 35692
rect 17880 35584 19748 35612
rect 11296 35516 12756 35544
rect 11296 35504 11302 35516
rect 12802 35504 12808 35556
rect 12860 35544 12866 35556
rect 17880 35544 17908 35584
rect 24762 35572 24768 35624
rect 24820 35612 24826 35624
rect 24857 35615 24915 35621
rect 24857 35612 24869 35615
rect 24820 35584 24869 35612
rect 24820 35572 24826 35584
rect 24857 35581 24869 35584
rect 24903 35581 24915 35615
rect 25130 35612 25136 35624
rect 25091 35584 25136 35612
rect 24857 35575 24915 35581
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 27430 35612 27436 35624
rect 27391 35584 27436 35612
rect 27430 35572 27436 35584
rect 27488 35572 27494 35624
rect 27706 35572 27712 35624
rect 27764 35612 27770 35624
rect 27982 35612 27988 35624
rect 27764 35584 27988 35612
rect 27764 35572 27770 35584
rect 27982 35572 27988 35584
rect 28040 35572 28046 35624
rect 29380 35612 29408 35666
rect 30243 35652 30288 35680
rect 30282 35640 30288 35652
rect 30340 35640 30346 35692
rect 30377 35683 30435 35689
rect 30377 35649 30389 35683
rect 30423 35680 30435 35683
rect 30466 35680 30472 35692
rect 30423 35652 30472 35680
rect 30423 35649 30435 35652
rect 30377 35643 30435 35649
rect 30466 35640 30472 35652
rect 30524 35680 30530 35692
rect 30834 35680 30840 35692
rect 30524 35652 30840 35680
rect 30524 35640 30530 35652
rect 30834 35640 30840 35652
rect 30892 35640 30898 35692
rect 30926 35640 30932 35692
rect 30984 35680 30990 35692
rect 31205 35683 31263 35689
rect 31205 35680 31217 35683
rect 30984 35652 31217 35680
rect 30984 35640 30990 35652
rect 31205 35649 31217 35652
rect 31251 35649 31263 35683
rect 31205 35643 31263 35649
rect 32309 35683 32367 35689
rect 32309 35649 32321 35683
rect 32355 35649 32367 35683
rect 32309 35643 32367 35649
rect 34885 35683 34943 35689
rect 34885 35649 34897 35683
rect 34931 35680 34943 35683
rect 35529 35683 35587 35689
rect 35529 35680 35541 35683
rect 34931 35652 35541 35680
rect 34931 35649 34943 35652
rect 34885 35643 34943 35649
rect 35529 35649 35541 35652
rect 35575 35680 35587 35683
rect 35802 35680 35808 35692
rect 35575 35652 35808 35680
rect 35575 35649 35587 35652
rect 35529 35643 35587 35649
rect 32324 35612 32352 35643
rect 35802 35640 35808 35652
rect 35860 35640 35866 35692
rect 36725 35683 36783 35689
rect 36725 35649 36737 35683
rect 36771 35649 36783 35683
rect 36725 35643 36783 35649
rect 35434 35612 35440 35624
rect 28092 35584 29408 35612
rect 31036 35584 32352 35612
rect 32784 35584 35440 35612
rect 28092 35544 28120 35584
rect 31036 35553 31064 35584
rect 31021 35547 31079 35553
rect 12860 35516 17908 35544
rect 26160 35516 28120 35544
rect 29288 35516 30512 35544
rect 12860 35504 12866 35516
rect 11698 35476 11704 35488
rect 8772 35448 11704 35476
rect 11698 35436 11704 35448
rect 11756 35436 11762 35488
rect 11882 35476 11888 35488
rect 11843 35448 11888 35476
rect 11882 35436 11888 35448
rect 11940 35436 11946 35488
rect 12066 35436 12072 35488
rect 12124 35476 12130 35488
rect 13814 35476 13820 35488
rect 12124 35448 13820 35476
rect 12124 35436 12130 35448
rect 13814 35436 13820 35448
rect 13872 35436 13878 35488
rect 14826 35476 14832 35488
rect 14787 35448 14832 35476
rect 14826 35436 14832 35448
rect 14884 35436 14890 35488
rect 15470 35476 15476 35488
rect 15431 35448 15476 35476
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 16117 35479 16175 35485
rect 16117 35445 16129 35479
rect 16163 35476 16175 35479
rect 17218 35476 17224 35488
rect 16163 35448 17224 35476
rect 16163 35445 16175 35448
rect 16117 35439 16175 35445
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 19889 35479 19947 35485
rect 19889 35445 19901 35479
rect 19935 35476 19947 35479
rect 19978 35476 19984 35488
rect 19935 35448 19984 35476
rect 19935 35445 19947 35448
rect 19889 35439 19947 35445
rect 19978 35436 19984 35448
rect 20036 35436 20042 35488
rect 20990 35436 20996 35488
rect 21048 35476 21054 35488
rect 23842 35476 23848 35488
rect 21048 35448 23848 35476
rect 21048 35436 21054 35448
rect 23842 35436 23848 35448
rect 23900 35436 23906 35488
rect 24854 35436 24860 35488
rect 24912 35476 24918 35488
rect 26160 35476 26188 35516
rect 24912 35448 26188 35476
rect 24912 35436 24918 35448
rect 26510 35436 26516 35488
rect 26568 35476 26574 35488
rect 26605 35479 26663 35485
rect 26605 35476 26617 35479
rect 26568 35448 26617 35476
rect 26568 35436 26574 35448
rect 26605 35445 26617 35448
rect 26651 35445 26663 35479
rect 26605 35439 26663 35445
rect 27522 35436 27528 35488
rect 27580 35476 27586 35488
rect 29288 35476 29316 35516
rect 27580 35448 29316 35476
rect 27580 35436 27586 35448
rect 29362 35436 29368 35488
rect 29420 35476 29426 35488
rect 29733 35479 29791 35485
rect 29733 35476 29745 35479
rect 29420 35448 29745 35476
rect 29420 35436 29426 35448
rect 29733 35445 29745 35448
rect 29779 35445 29791 35479
rect 30484 35476 30512 35516
rect 31021 35513 31033 35547
rect 31067 35513 31079 35547
rect 32784 35544 32812 35584
rect 35434 35572 35440 35584
rect 35492 35572 35498 35624
rect 36740 35612 36768 35643
rect 36814 35640 36820 35692
rect 36872 35680 36878 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 36872 35652 38025 35680
rect 36872 35640 36878 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 38286 35612 38292 35624
rect 36740 35584 38292 35612
rect 38286 35572 38292 35584
rect 38344 35572 38350 35624
rect 31021 35507 31079 35513
rect 31128 35516 32812 35544
rect 31128 35476 31156 35516
rect 32858 35504 32864 35556
rect 32916 35544 32922 35556
rect 35986 35544 35992 35556
rect 32916 35516 35992 35544
rect 32916 35504 32922 35516
rect 35986 35504 35992 35516
rect 36044 35504 36050 35556
rect 30484 35448 31156 35476
rect 29733 35439 29791 35445
rect 31478 35436 31484 35488
rect 31536 35476 31542 35488
rect 32401 35479 32459 35485
rect 32401 35476 32413 35479
rect 31536 35448 32413 35476
rect 31536 35436 31542 35448
rect 32401 35445 32413 35448
rect 32447 35445 32459 35479
rect 32401 35439 32459 35445
rect 34698 35436 34704 35488
rect 34756 35476 34762 35488
rect 34977 35479 35035 35485
rect 34977 35476 34989 35479
rect 34756 35448 34989 35476
rect 34756 35436 34762 35448
rect 34977 35445 34989 35448
rect 35023 35445 35035 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 34977 35439 35035 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 7653 35275 7711 35281
rect 7653 35241 7665 35275
rect 7699 35272 7711 35275
rect 7834 35272 7840 35284
rect 7699 35244 7840 35272
rect 7699 35241 7711 35244
rect 7653 35235 7711 35241
rect 7834 35232 7840 35244
rect 7892 35232 7898 35284
rect 10318 35272 10324 35284
rect 10279 35244 10324 35272
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 11054 35272 11060 35284
rect 11015 35244 11060 35272
rect 11054 35232 11060 35244
rect 11112 35232 11118 35284
rect 13446 35272 13452 35284
rect 12636 35244 13452 35272
rect 6549 35207 6607 35213
rect 6549 35173 6561 35207
rect 6595 35204 6607 35207
rect 11701 35207 11759 35213
rect 6595 35176 9352 35204
rect 6595 35173 6607 35176
rect 6549 35167 6607 35173
rect 6638 35136 6644 35148
rect 4356 35108 6644 35136
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35068 1823 35071
rect 2866 35068 2872 35080
rect 1811 35040 2872 35068
rect 1811 35037 1823 35040
rect 1765 35031 1823 35037
rect 2866 35028 2872 35040
rect 2924 35028 2930 35080
rect 4356 35077 4384 35108
rect 6638 35096 6644 35108
rect 6696 35096 6702 35148
rect 8478 35136 8484 35148
rect 7576 35108 8484 35136
rect 4341 35071 4399 35077
rect 4341 35037 4353 35071
rect 4387 35037 4399 35071
rect 4341 35031 4399 35037
rect 5626 35028 5632 35080
rect 5684 35068 5690 35080
rect 7576 35077 7604 35108
rect 8478 35096 8484 35108
rect 8536 35096 8542 35148
rect 8846 35096 8852 35148
rect 8904 35136 8910 35148
rect 9324 35145 9352 35176
rect 11701 35173 11713 35207
rect 11747 35204 11759 35207
rect 12636 35204 12664 35244
rect 13446 35232 13452 35244
rect 13504 35232 13510 35284
rect 13630 35272 13636 35284
rect 13591 35244 13636 35272
rect 13630 35232 13636 35244
rect 13688 35232 13694 35284
rect 14734 35232 14740 35284
rect 14792 35272 14798 35284
rect 16574 35272 16580 35284
rect 14792 35244 16580 35272
rect 14792 35232 14798 35244
rect 16574 35232 16580 35244
rect 16632 35232 16638 35284
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18012 35244 22094 35272
rect 18012 35232 18018 35244
rect 21266 35204 21272 35216
rect 11747 35176 12664 35204
rect 12728 35176 21272 35204
rect 11747 35173 11759 35176
rect 11701 35167 11759 35173
rect 9125 35139 9183 35145
rect 9125 35136 9137 35139
rect 8904 35108 9137 35136
rect 8904 35096 8910 35108
rect 9125 35105 9137 35108
rect 9171 35105 9183 35139
rect 9125 35099 9183 35105
rect 9309 35139 9367 35145
rect 9309 35105 9321 35139
rect 9355 35105 9367 35139
rect 9309 35099 9367 35105
rect 11882 35096 11888 35148
rect 11940 35136 11946 35148
rect 12618 35136 12624 35148
rect 11940 35108 12624 35136
rect 11940 35096 11946 35108
rect 12618 35096 12624 35108
rect 12676 35096 12682 35148
rect 6733 35071 6791 35077
rect 6733 35068 6745 35071
rect 5684 35040 6745 35068
rect 5684 35028 5690 35040
rect 6733 35037 6745 35040
rect 6779 35037 6791 35071
rect 6733 35031 6791 35037
rect 7561 35071 7619 35077
rect 7561 35037 7573 35071
rect 7607 35037 7619 35071
rect 7561 35031 7619 35037
rect 8389 35071 8447 35077
rect 8389 35037 8401 35071
rect 8435 35068 8447 35071
rect 8662 35068 8668 35080
rect 8435 35040 8668 35068
rect 8435 35037 8447 35040
rect 8389 35031 8447 35037
rect 8662 35028 8668 35040
rect 8720 35028 8726 35080
rect 10229 35071 10287 35077
rect 10229 35037 10241 35071
rect 10275 35068 10287 35071
rect 10778 35068 10784 35080
rect 10275 35040 10784 35068
rect 10275 35037 10287 35040
rect 10229 35031 10287 35037
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 10962 35068 10968 35080
rect 10923 35040 10968 35068
rect 10962 35028 10968 35040
rect 11020 35028 11026 35080
rect 11609 35071 11667 35077
rect 11609 35037 11621 35071
rect 11655 35068 11667 35071
rect 11974 35068 11980 35080
rect 11655 35040 11980 35068
rect 11655 35037 11667 35040
rect 11609 35031 11667 35037
rect 11974 35028 11980 35040
rect 12032 35028 12038 35080
rect 12253 35071 12311 35077
rect 12253 35037 12265 35071
rect 12299 35037 12311 35071
rect 12253 35031 12311 35037
rect 6822 35000 6828 35012
rect 1596 34972 6828 35000
rect 1596 34941 1624 34972
rect 6822 34960 6828 34972
rect 6880 34960 6886 35012
rect 9416 34972 10640 35000
rect 9416 34944 9444 34972
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34901 1639 34935
rect 1581 34895 1639 34901
rect 2958 34892 2964 34944
rect 3016 34932 3022 34944
rect 4157 34935 4215 34941
rect 4157 34932 4169 34935
rect 3016 34904 4169 34932
rect 3016 34892 3022 34904
rect 4157 34901 4169 34904
rect 4203 34901 4215 34935
rect 4157 34895 4215 34901
rect 8481 34935 8539 34941
rect 8481 34901 8493 34935
rect 8527 34932 8539 34935
rect 9398 34932 9404 34944
rect 8527 34904 9404 34932
rect 8527 34901 8539 34904
rect 8481 34895 8539 34901
rect 9398 34892 9404 34904
rect 9456 34892 9462 34944
rect 9766 34932 9772 34944
rect 9727 34904 9772 34932
rect 9766 34892 9772 34904
rect 9824 34892 9830 34944
rect 10612 34932 10640 34972
rect 10870 34960 10876 35012
rect 10928 35000 10934 35012
rect 12268 35000 12296 35031
rect 10928 34972 12296 35000
rect 12345 35003 12403 35009
rect 10928 34960 10934 34972
rect 12345 34969 12357 35003
rect 12391 35000 12403 35003
rect 12728 35000 12756 35176
rect 21266 35164 21272 35176
rect 21324 35164 21330 35216
rect 22066 35204 22094 35244
rect 23842 35232 23848 35284
rect 23900 35272 23906 35284
rect 23900 35244 34192 35272
rect 23900 35232 23906 35244
rect 24854 35204 24860 35216
rect 22066 35176 24860 35204
rect 24854 35164 24860 35176
rect 24912 35164 24918 35216
rect 14553 35139 14611 35145
rect 14553 35136 14565 35139
rect 12391 34972 12756 35000
rect 12820 35108 14565 35136
rect 12391 34969 12403 34972
rect 12345 34963 12403 34969
rect 12158 34932 12164 34944
rect 10612 34904 12164 34932
rect 12158 34892 12164 34904
rect 12216 34932 12222 34944
rect 12820 34932 12848 35108
rect 14553 35105 14565 35108
rect 14599 35105 14611 35139
rect 14553 35099 14611 35105
rect 15470 35096 15476 35148
rect 15528 35136 15534 35148
rect 20714 35136 20720 35148
rect 15528 35108 20720 35136
rect 15528 35096 15534 35108
rect 20714 35096 20720 35108
rect 20772 35096 20778 35148
rect 24302 35096 24308 35148
rect 24360 35136 24366 35148
rect 24762 35136 24768 35148
rect 24360 35108 24768 35136
rect 24360 35096 24366 35108
rect 24762 35096 24768 35108
rect 24820 35136 24826 35148
rect 24949 35139 25007 35145
rect 24949 35136 24961 35139
rect 24820 35108 24961 35136
rect 24820 35096 24826 35108
rect 24949 35105 24961 35108
rect 24995 35136 25007 35139
rect 31478 35136 31484 35148
rect 24995 35108 26648 35136
rect 31439 35108 31484 35136
rect 24995 35105 25007 35108
rect 24949 35099 25007 35105
rect 12897 35071 12955 35077
rect 12897 35037 12909 35071
rect 12943 35068 12955 35071
rect 13262 35068 13268 35080
rect 12943 35040 13268 35068
rect 12943 35037 12955 35040
rect 12897 35031 12955 35037
rect 13262 35028 13268 35040
rect 13320 35028 13326 35080
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35068 13599 35071
rect 13814 35068 13820 35080
rect 13587 35040 13820 35068
rect 13587 35037 13599 35040
rect 13541 35031 13599 35037
rect 13814 35028 13820 35040
rect 13872 35028 13878 35080
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 15396 35040 16405 35068
rect 12989 35003 13047 35009
rect 12989 34969 13001 35003
rect 13035 35000 13047 35003
rect 14642 35000 14648 35012
rect 13035 34972 14504 35000
rect 14603 34972 14648 35000
rect 13035 34969 13047 34972
rect 12989 34963 13047 34969
rect 12216 34904 12848 34932
rect 12216 34892 12222 34904
rect 13446 34892 13452 34944
rect 13504 34932 13510 34944
rect 14366 34932 14372 34944
rect 13504 34904 14372 34932
rect 13504 34892 13510 34904
rect 14366 34892 14372 34904
rect 14424 34892 14430 34944
rect 14476 34932 14504 34972
rect 14642 34960 14648 34972
rect 14700 34960 14706 35012
rect 14918 34960 14924 35012
rect 14976 35000 14982 35012
rect 15396 35000 15424 35040
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 20806 35068 20812 35080
rect 16393 35031 16451 35037
rect 17788 35040 20812 35068
rect 15562 35000 15568 35012
rect 14976 34972 15424 35000
rect 15523 34972 15568 35000
rect 14976 34960 14982 34972
rect 15562 34960 15568 34972
rect 15620 34960 15626 35012
rect 16574 35000 16580 35012
rect 16535 34972 16580 35000
rect 16574 34960 16580 34972
rect 16632 34960 16638 35012
rect 16666 34960 16672 35012
rect 16724 35000 16730 35012
rect 17788 35000 17816 35040
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 26620 35012 26648 35108
rect 31478 35096 31484 35108
rect 31536 35096 31542 35148
rect 31846 35136 31852 35148
rect 31807 35108 31852 35136
rect 31846 35096 31852 35108
rect 31904 35096 31910 35148
rect 32214 35096 32220 35148
rect 32272 35136 32278 35148
rect 32585 35139 32643 35145
rect 32585 35136 32597 35139
rect 32272 35108 32597 35136
rect 32272 35096 32278 35108
rect 32585 35105 32597 35108
rect 32631 35136 32643 35139
rect 32950 35136 32956 35148
rect 32631 35108 32956 35136
rect 32631 35105 32643 35108
rect 32585 35099 32643 35105
rect 32950 35096 32956 35108
rect 33008 35096 33014 35148
rect 34164 35136 34192 35244
rect 34514 35232 34520 35284
rect 34572 35272 34578 35284
rect 34977 35275 35035 35281
rect 34977 35272 34989 35275
rect 34572 35244 34989 35272
rect 34572 35232 34578 35244
rect 34977 35241 34989 35244
rect 35023 35241 35035 35275
rect 34977 35235 35035 35241
rect 36725 35275 36783 35281
rect 36725 35241 36737 35275
rect 36771 35272 36783 35275
rect 36814 35272 36820 35284
rect 36771 35244 36820 35272
rect 36771 35241 36783 35244
rect 36725 35235 36783 35241
rect 36814 35232 36820 35244
rect 36872 35232 36878 35284
rect 37369 35275 37427 35281
rect 37369 35241 37381 35275
rect 37415 35272 37427 35275
rect 38010 35272 38016 35284
rect 37415 35244 38016 35272
rect 37415 35241 37427 35244
rect 37369 35235 37427 35241
rect 38010 35232 38016 35244
rect 38068 35232 38074 35284
rect 38197 35275 38255 35281
rect 38197 35241 38209 35275
rect 38243 35272 38255 35275
rect 39298 35272 39304 35284
rect 38243 35244 39304 35272
rect 38243 35241 38255 35244
rect 38197 35235 38255 35241
rect 39298 35232 39304 35244
rect 39356 35232 39362 35284
rect 34330 35164 34336 35216
rect 34388 35204 34394 35216
rect 34388 35176 35894 35204
rect 34388 35164 34394 35176
rect 34164 35108 34928 35136
rect 26786 35028 26792 35080
rect 26844 35068 26850 35080
rect 34900 35077 34928 35108
rect 27157 35071 27215 35077
rect 27157 35068 27169 35071
rect 26844 35040 27169 35068
rect 26844 35028 26850 35040
rect 27157 35037 27169 35040
rect 27203 35068 27215 35071
rect 34885 35071 34943 35077
rect 27203 35040 28994 35068
rect 27203 35037 27215 35040
rect 27157 35031 27215 35037
rect 16724 34972 17816 35000
rect 18233 35003 18291 35009
rect 16724 34960 16730 34972
rect 18233 34969 18245 35003
rect 18279 35000 18291 35003
rect 19150 35000 19156 35012
rect 18279 34972 19156 35000
rect 18279 34969 18291 34972
rect 18233 34963 18291 34969
rect 19150 34960 19156 34972
rect 19208 34960 19214 35012
rect 20622 34960 20628 35012
rect 20680 35000 20686 35012
rect 20993 35003 21051 35009
rect 20993 35000 21005 35003
rect 20680 34972 21005 35000
rect 20680 34960 20686 34972
rect 20993 34969 21005 34972
rect 21039 34969 21051 35003
rect 20993 34963 21051 34969
rect 21821 35003 21879 35009
rect 21821 34969 21833 35003
rect 21867 35000 21879 35003
rect 22002 35000 22008 35012
rect 21867 34972 22008 35000
rect 21867 34969 21879 34972
rect 21821 34963 21879 34969
rect 22002 34960 22008 34972
rect 22060 34960 22066 35012
rect 24946 34960 24952 35012
rect 25004 35000 25010 35012
rect 25225 35003 25283 35009
rect 25225 35000 25237 35003
rect 25004 34972 25237 35000
rect 25004 34960 25010 34972
rect 25225 34969 25237 34972
rect 25271 34969 25283 35003
rect 25225 34963 25283 34969
rect 26234 34960 26240 35012
rect 26292 34960 26298 35012
rect 26602 34960 26608 35012
rect 26660 35000 26666 35012
rect 27893 35003 27951 35009
rect 27893 35000 27905 35003
rect 26660 34972 27905 35000
rect 26660 34960 26666 34972
rect 27893 34969 27905 34972
rect 27939 34969 27951 35003
rect 28966 35000 28994 35040
rect 34885 35037 34897 35071
rect 34931 35037 34943 35071
rect 35866 35068 35894 35176
rect 36081 35071 36139 35077
rect 36081 35068 36093 35071
rect 35866 35040 36093 35068
rect 34885 35031 34943 35037
rect 36081 35037 36093 35040
rect 36127 35037 36139 35071
rect 36081 35031 36139 35037
rect 36446 35028 36452 35080
rect 36504 35068 36510 35080
rect 36909 35071 36967 35077
rect 36909 35068 36921 35071
rect 36504 35040 36921 35068
rect 36504 35028 36510 35040
rect 36909 35037 36921 35040
rect 36955 35037 36967 35071
rect 37550 35068 37556 35080
rect 37511 35040 37556 35068
rect 36909 35031 36967 35037
rect 37550 35028 37556 35040
rect 37608 35028 37614 35080
rect 37918 35028 37924 35080
rect 37976 35068 37982 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 37976 35040 38025 35068
rect 37976 35028 37982 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 29730 35000 29736 35012
rect 28966 34972 29736 35000
rect 27893 34963 27951 34969
rect 29730 34960 29736 34972
rect 29788 34960 29794 35012
rect 30558 35000 30564 35012
rect 30519 34972 30564 35000
rect 30558 34960 30564 34972
rect 30616 34960 30622 35012
rect 31570 34960 31576 35012
rect 31628 35000 31634 35012
rect 32858 35000 32864 35012
rect 31628 34972 31673 35000
rect 32819 34972 32864 35000
rect 31628 34960 31634 34972
rect 32858 34960 32864 34972
rect 32916 34960 32922 35012
rect 36814 35000 36820 35012
rect 34086 34972 36820 35000
rect 36814 34960 36820 34972
rect 36872 34960 36878 35012
rect 22554 34932 22560 34944
rect 14476 34904 22560 34932
rect 22554 34892 22560 34904
rect 22612 34892 22618 34944
rect 26694 34932 26700 34944
rect 26655 34904 26700 34932
rect 26694 34892 26700 34904
rect 26752 34892 26758 34944
rect 27430 34892 27436 34944
rect 27488 34932 27494 34944
rect 31018 34932 31024 34944
rect 27488 34904 31024 34932
rect 27488 34892 27494 34904
rect 31018 34892 31024 34904
rect 31076 34892 31082 34944
rect 34330 34932 34336 34944
rect 34291 34904 34336 34932
rect 34330 34892 34336 34904
rect 34388 34892 34394 34944
rect 36170 34932 36176 34944
rect 36131 34904 36176 34932
rect 36170 34892 36176 34904
rect 36228 34892 36234 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1762 34688 1768 34740
rect 1820 34728 1826 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 1820 34700 2421 34728
rect 1820 34688 1826 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 8662 34728 8668 34740
rect 2409 34691 2467 34697
rect 2746 34700 8668 34728
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 2317 34595 2375 34601
rect 2317 34561 2329 34595
rect 2363 34592 2375 34595
rect 2746 34592 2774 34700
rect 8662 34688 8668 34700
rect 8720 34688 8726 34740
rect 9766 34688 9772 34740
rect 9824 34728 9830 34740
rect 9824 34700 11468 34728
rect 9824 34688 9830 34700
rect 8478 34620 8484 34672
rect 8536 34660 8542 34672
rect 10686 34660 10692 34672
rect 8536 34632 10692 34660
rect 8536 34620 8542 34632
rect 10686 34620 10692 34632
rect 10744 34620 10750 34672
rect 11440 34660 11468 34700
rect 11974 34688 11980 34740
rect 12032 34728 12038 34740
rect 13262 34728 13268 34740
rect 12032 34700 13268 34728
rect 12032 34688 12038 34700
rect 13262 34688 13268 34700
rect 13320 34688 13326 34740
rect 13630 34688 13636 34740
rect 13688 34728 13694 34740
rect 14642 34728 14648 34740
rect 13688 34700 14648 34728
rect 13688 34688 13694 34700
rect 14642 34688 14648 34700
rect 14700 34688 14706 34740
rect 14826 34688 14832 34740
rect 14884 34728 14890 34740
rect 19610 34728 19616 34740
rect 14884 34700 19616 34728
rect 14884 34688 14890 34700
rect 19610 34688 19616 34700
rect 19668 34688 19674 34740
rect 21450 34728 21456 34740
rect 19720 34700 21456 34728
rect 11793 34663 11851 34669
rect 11793 34660 11805 34663
rect 11440 34632 11805 34660
rect 11793 34629 11805 34632
rect 11839 34629 11851 34663
rect 11793 34623 11851 34629
rect 11882 34620 11888 34672
rect 11940 34660 11946 34672
rect 13541 34663 13599 34669
rect 13541 34660 13553 34663
rect 11940 34632 11985 34660
rect 13004 34632 13553 34660
rect 11940 34620 11946 34632
rect 8294 34592 8300 34604
rect 2363 34564 2774 34592
rect 8255 34564 8300 34592
rect 2363 34561 2375 34564
rect 2317 34555 2375 34561
rect 8294 34552 8300 34564
rect 8352 34552 8358 34604
rect 8389 34595 8447 34601
rect 8389 34561 8401 34595
rect 8435 34592 8447 34595
rect 9585 34595 9643 34601
rect 9585 34592 9597 34595
rect 8435 34564 9597 34592
rect 8435 34561 8447 34564
rect 8389 34555 8447 34561
rect 9585 34561 9597 34564
rect 9631 34561 9643 34595
rect 9585 34555 9643 34561
rect 10965 34595 11023 34601
rect 10965 34561 10977 34595
rect 11011 34592 11023 34595
rect 11606 34592 11612 34604
rect 11011 34564 11612 34592
rect 11011 34561 11023 34564
rect 10965 34555 11023 34561
rect 11606 34552 11612 34564
rect 11664 34552 11670 34604
rect 8312 34524 8340 34552
rect 9214 34524 9220 34536
rect 8312 34496 9220 34524
rect 9214 34484 9220 34496
rect 9272 34484 9278 34536
rect 9398 34524 9404 34536
rect 9359 34496 9404 34524
rect 9398 34484 9404 34496
rect 9456 34484 9462 34536
rect 11057 34527 11115 34533
rect 11057 34493 11069 34527
rect 11103 34524 11115 34527
rect 11146 34524 11152 34536
rect 11103 34496 11152 34524
rect 11103 34493 11115 34496
rect 11057 34487 11115 34493
rect 11146 34484 11152 34496
rect 11204 34484 11210 34536
rect 13004 34524 13032 34632
rect 13541 34629 13553 34632
rect 13587 34629 13599 34663
rect 13541 34623 13599 34629
rect 13906 34620 13912 34672
rect 13964 34660 13970 34672
rect 14093 34663 14151 34669
rect 14093 34660 14105 34663
rect 13964 34632 14105 34660
rect 13964 34620 13970 34632
rect 14093 34629 14105 34632
rect 14139 34660 14151 34663
rect 14458 34660 14464 34672
rect 14139 34632 14464 34660
rect 14139 34629 14151 34632
rect 14093 34623 14151 34629
rect 14458 34620 14464 34632
rect 14516 34660 14522 34672
rect 15010 34660 15016 34672
rect 14516 34632 15016 34660
rect 14516 34620 14522 34632
rect 15010 34620 15016 34632
rect 15068 34620 15074 34672
rect 15749 34663 15807 34669
rect 15749 34629 15761 34663
rect 15795 34660 15807 34663
rect 17494 34660 17500 34672
rect 15795 34632 17500 34660
rect 15795 34629 15807 34632
rect 15749 34623 15807 34629
rect 17494 34620 17500 34632
rect 17552 34620 17558 34672
rect 14553 34595 14611 34601
rect 14553 34561 14565 34595
rect 14599 34561 14611 34595
rect 14553 34555 14611 34561
rect 14645 34595 14703 34601
rect 14645 34561 14657 34595
rect 14691 34592 14703 34595
rect 14734 34592 14740 34604
rect 14691 34564 14740 34592
rect 14691 34561 14703 34564
rect 14645 34555 14703 34561
rect 11256 34496 13032 34524
rect 13449 34527 13507 34533
rect 9766 34456 9772 34468
rect 9727 34428 9772 34456
rect 9766 34416 9772 34428
rect 9824 34416 9830 34468
rect 10962 34416 10968 34468
rect 11020 34456 11026 34468
rect 11256 34456 11284 34496
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13538 34524 13544 34536
rect 13495 34496 13544 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13538 34484 13544 34496
rect 13596 34484 13602 34536
rect 14568 34524 14596 34555
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 17218 34592 17224 34604
rect 17179 34564 17224 34592
rect 17218 34552 17224 34564
rect 17276 34552 17282 34604
rect 19720 34592 19748 34700
rect 21450 34688 21456 34700
rect 21508 34688 21514 34740
rect 21542 34688 21548 34740
rect 21600 34728 21606 34740
rect 21600 34700 24900 34728
rect 21600 34688 21606 34700
rect 19886 34620 19892 34672
rect 19944 34660 19950 34672
rect 19944 34632 20470 34660
rect 19944 34620 19950 34632
rect 21266 34620 21272 34672
rect 21324 34660 21330 34672
rect 24872 34660 24900 34700
rect 27982 34688 27988 34740
rect 28040 34728 28046 34740
rect 30558 34728 30564 34740
rect 28040 34700 30564 34728
rect 28040 34688 28046 34700
rect 21324 34632 22770 34660
rect 24872 34632 25070 34660
rect 21324 34620 21330 34632
rect 24302 34592 24308 34604
rect 19306 34564 19748 34592
rect 24263 34564 24308 34592
rect 15657 34527 15715 34533
rect 14568 34496 15608 34524
rect 12342 34456 12348 34468
rect 11020 34428 11284 34456
rect 12303 34428 12348 34456
rect 11020 34416 11026 34428
rect 12342 34416 12348 34428
rect 12400 34456 12406 34468
rect 13722 34456 13728 34468
rect 12400 34428 13728 34456
rect 12400 34416 12406 34428
rect 13722 34416 13728 34428
rect 13780 34416 13786 34468
rect 15580 34456 15608 34496
rect 15657 34493 15669 34527
rect 15703 34524 15715 34527
rect 15930 34524 15936 34536
rect 15703 34496 15936 34524
rect 15703 34493 15715 34496
rect 15657 34487 15715 34493
rect 15930 34484 15936 34496
rect 15988 34484 15994 34536
rect 19306 34524 19334 34564
rect 24302 34552 24308 34564
rect 24360 34552 24366 34604
rect 29288 34601 29316 34700
rect 30558 34688 30564 34700
rect 30616 34688 30622 34740
rect 32953 34731 33011 34737
rect 32953 34697 32965 34731
rect 32999 34728 33011 34731
rect 35345 34731 35403 34737
rect 35345 34728 35357 34731
rect 32999 34700 35357 34728
rect 32999 34697 33011 34700
rect 32953 34691 33011 34697
rect 35345 34697 35357 34700
rect 35391 34697 35403 34731
rect 36814 34728 36820 34740
rect 36775 34700 36820 34728
rect 35345 34691 35403 34697
rect 31478 34660 31484 34672
rect 30774 34632 31484 34660
rect 31478 34620 31484 34632
rect 31536 34620 31542 34672
rect 33410 34620 33416 34672
rect 33468 34660 33474 34672
rect 33468 34632 34284 34660
rect 33468 34620 33474 34632
rect 29273 34595 29331 34601
rect 29273 34561 29285 34595
rect 29319 34561 29331 34595
rect 29273 34555 29331 34561
rect 30834 34552 30840 34604
rect 30892 34592 30898 34604
rect 32309 34595 32367 34601
rect 32309 34592 32321 34595
rect 30892 34564 32321 34592
rect 30892 34552 30898 34564
rect 32309 34561 32321 34564
rect 32355 34561 32367 34595
rect 32309 34555 32367 34561
rect 33597 34595 33655 34601
rect 33597 34561 33609 34595
rect 33643 34592 33655 34595
rect 34146 34592 34152 34604
rect 33643 34564 34152 34592
rect 33643 34561 33655 34564
rect 33597 34555 33655 34561
rect 34146 34552 34152 34564
rect 34204 34552 34210 34604
rect 34256 34601 34284 34632
rect 34241 34595 34299 34601
rect 34241 34561 34253 34595
rect 34287 34561 34299 34595
rect 34241 34555 34299 34561
rect 16040 34496 19334 34524
rect 19705 34527 19763 34533
rect 16040 34456 16068 34496
rect 19705 34493 19717 34527
rect 19751 34524 19763 34527
rect 19981 34527 20039 34533
rect 19751 34496 19840 34524
rect 19751 34493 19763 34496
rect 19705 34487 19763 34493
rect 15580 34428 16068 34456
rect 16206 34416 16212 34468
rect 16264 34456 16270 34468
rect 16264 34428 16357 34456
rect 16264 34416 16270 34428
rect 18138 34416 18144 34468
rect 18196 34456 18202 34468
rect 19242 34456 19248 34468
rect 18196 34428 19248 34456
rect 18196 34416 18202 34428
rect 19242 34416 19248 34428
rect 19300 34416 19306 34468
rect 19610 34456 19616 34468
rect 19352 34428 19616 34456
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 10134 34348 10140 34400
rect 10192 34388 10198 34400
rect 16224 34388 16252 34416
rect 19352 34400 19380 34428
rect 19610 34416 19616 34428
rect 19668 34416 19674 34468
rect 10192 34360 16252 34388
rect 10192 34348 10198 34360
rect 17126 34348 17132 34400
rect 17184 34388 17190 34400
rect 17313 34391 17371 34397
rect 17313 34388 17325 34391
rect 17184 34360 17325 34388
rect 17184 34348 17190 34360
rect 17313 34357 17325 34360
rect 17359 34357 17371 34391
rect 17313 34351 17371 34357
rect 19334 34348 19340 34400
rect 19392 34348 19398 34400
rect 19426 34348 19432 34400
rect 19484 34388 19490 34400
rect 19812 34388 19840 34496
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20714 34524 20720 34536
rect 20027 34496 20720 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20714 34484 20720 34496
rect 20772 34484 20778 34536
rect 22002 34524 22008 34536
rect 21963 34496 22008 34524
rect 22002 34484 22008 34496
rect 22060 34484 22066 34536
rect 22278 34524 22284 34536
rect 22239 34496 22284 34524
rect 22278 34484 22284 34496
rect 22336 34484 22342 34536
rect 23750 34524 23756 34536
rect 23663 34496 23756 34524
rect 23750 34484 23756 34496
rect 23808 34524 23814 34536
rect 23934 34524 23940 34536
rect 23808 34496 23940 34524
rect 23808 34484 23814 34496
rect 23934 34484 23940 34496
rect 23992 34484 23998 34536
rect 24581 34527 24639 34533
rect 24581 34524 24593 34527
rect 24412 34496 24593 34524
rect 22020 34456 22048 34484
rect 24412 34456 24440 34496
rect 24581 34493 24593 34496
rect 24627 34493 24639 34527
rect 24581 34487 24639 34493
rect 24670 34484 24676 34536
rect 24728 34524 24734 34536
rect 26053 34527 26111 34533
rect 26053 34524 26065 34527
rect 24728 34496 26065 34524
rect 24728 34484 24734 34496
rect 26053 34493 26065 34496
rect 26099 34493 26111 34527
rect 29549 34527 29607 34533
rect 29549 34524 29561 34527
rect 26053 34487 26111 34493
rect 29380 34496 29561 34524
rect 21008 34428 22048 34456
rect 23308 34428 24440 34456
rect 21008 34388 21036 34428
rect 19484 34360 21036 34388
rect 19484 34348 19490 34360
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 23308 34388 23336 34428
rect 26510 34416 26516 34468
rect 26568 34456 26574 34468
rect 29380 34456 29408 34496
rect 29549 34493 29561 34496
rect 29595 34493 29607 34527
rect 29549 34487 29607 34493
rect 30742 34484 30748 34536
rect 30800 34524 30806 34536
rect 31294 34524 31300 34536
rect 30800 34496 31300 34524
rect 30800 34484 30806 34496
rect 31294 34484 31300 34496
rect 31352 34484 31358 34536
rect 32493 34527 32551 34533
rect 32493 34493 32505 34527
rect 32539 34524 32551 34527
rect 32539 34496 34100 34524
rect 32539 34493 32551 34496
rect 32493 34487 32551 34493
rect 33410 34456 33416 34468
rect 26568 34428 29408 34456
rect 33371 34428 33416 34456
rect 26568 34416 26574 34428
rect 33410 34416 33416 34428
rect 33468 34416 33474 34468
rect 34072 34465 34100 34496
rect 34606 34484 34612 34536
rect 34664 34524 34670 34536
rect 34701 34527 34759 34533
rect 34701 34524 34713 34527
rect 34664 34496 34713 34524
rect 34664 34484 34670 34496
rect 34701 34493 34713 34496
rect 34747 34493 34759 34527
rect 34701 34487 34759 34493
rect 34790 34484 34796 34536
rect 34848 34524 34854 34536
rect 34885 34527 34943 34533
rect 34885 34524 34897 34527
rect 34848 34496 34897 34524
rect 34848 34484 34854 34496
rect 34885 34493 34897 34496
rect 34931 34493 34943 34527
rect 35360 34524 35388 34691
rect 36814 34688 36820 34700
rect 36872 34688 36878 34740
rect 35618 34620 35624 34672
rect 35676 34660 35682 34672
rect 35676 34632 36768 34660
rect 35676 34620 35682 34632
rect 36740 34601 36768 34632
rect 36265 34595 36323 34601
rect 36265 34561 36277 34595
rect 36311 34561 36323 34595
rect 36265 34555 36323 34561
rect 36725 34595 36783 34601
rect 36725 34561 36737 34595
rect 36771 34561 36783 34595
rect 36725 34555 36783 34561
rect 38013 34595 38071 34601
rect 38013 34561 38025 34595
rect 38059 34592 38071 34595
rect 39022 34592 39028 34604
rect 38059 34564 39028 34592
rect 38059 34561 38071 34564
rect 38013 34555 38071 34561
rect 35894 34524 35900 34536
rect 35360 34496 35900 34524
rect 34885 34487 34943 34493
rect 35894 34484 35900 34496
rect 35952 34484 35958 34536
rect 36280 34524 36308 34555
rect 39022 34552 39028 34564
rect 39080 34552 39086 34604
rect 38654 34524 38660 34536
rect 36280 34496 38660 34524
rect 38654 34484 38660 34496
rect 38712 34484 38718 34536
rect 34057 34459 34115 34465
rect 34057 34425 34069 34459
rect 34103 34425 34115 34459
rect 34057 34419 34115 34425
rect 21140 34360 23336 34388
rect 21140 34348 21146 34360
rect 26418 34348 26424 34400
rect 26476 34388 26482 34400
rect 35618 34388 35624 34400
rect 26476 34360 35624 34388
rect 26476 34348 26482 34360
rect 35618 34348 35624 34360
rect 35676 34348 35682 34400
rect 36078 34388 36084 34400
rect 36039 34360 36084 34388
rect 36078 34348 36084 34360
rect 36136 34348 36142 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 8478 34184 8484 34196
rect 8439 34156 8484 34184
rect 8478 34144 8484 34156
rect 8536 34144 8542 34196
rect 10226 34144 10232 34196
rect 10284 34184 10290 34196
rect 11422 34184 11428 34196
rect 10284 34156 11428 34184
rect 10284 34144 10290 34156
rect 11422 34144 11428 34156
rect 11480 34144 11486 34196
rect 11517 34187 11575 34193
rect 11517 34153 11529 34187
rect 11563 34184 11575 34187
rect 13446 34184 13452 34196
rect 11563 34156 13452 34184
rect 11563 34153 11575 34156
rect 11517 34147 11575 34153
rect 13446 34144 13452 34156
rect 13504 34144 13510 34196
rect 13541 34187 13599 34193
rect 13541 34153 13553 34187
rect 13587 34184 13599 34187
rect 13630 34184 13636 34196
rect 13587 34156 13636 34184
rect 13587 34153 13599 34156
rect 13541 34147 13599 34153
rect 13630 34144 13636 34156
rect 13688 34144 13694 34196
rect 15562 34184 15568 34196
rect 13740 34156 15568 34184
rect 10873 34119 10931 34125
rect 10873 34085 10885 34119
rect 10919 34116 10931 34119
rect 12894 34116 12900 34128
rect 10919 34088 12900 34116
rect 10919 34085 10931 34088
rect 10873 34079 10931 34085
rect 12894 34076 12900 34088
rect 12952 34076 12958 34128
rect 12986 34076 12992 34128
rect 13044 34116 13050 34128
rect 13740 34116 13768 34156
rect 15562 34144 15568 34156
rect 15620 34144 15626 34196
rect 15654 34144 15660 34196
rect 15712 34184 15718 34196
rect 16485 34187 16543 34193
rect 16485 34184 16497 34187
rect 15712 34156 16497 34184
rect 15712 34144 15718 34156
rect 16485 34153 16497 34156
rect 16531 34153 16543 34187
rect 16485 34147 16543 34153
rect 16666 34144 16672 34196
rect 16724 34184 16730 34196
rect 19610 34184 19616 34196
rect 16724 34156 19616 34184
rect 16724 34144 16730 34156
rect 19610 34144 19616 34156
rect 19668 34144 19674 34196
rect 20254 34144 20260 34196
rect 20312 34184 20318 34196
rect 21082 34184 21088 34196
rect 20312 34156 21088 34184
rect 20312 34144 20318 34156
rect 21082 34144 21088 34156
rect 21140 34144 21146 34196
rect 26694 34184 26700 34196
rect 21652 34156 26700 34184
rect 13044 34088 13768 34116
rect 14645 34119 14703 34125
rect 13044 34076 13050 34088
rect 14645 34085 14657 34119
rect 14691 34116 14703 34119
rect 21542 34116 21548 34128
rect 14691 34088 21548 34116
rect 14691 34085 14703 34088
rect 14645 34079 14703 34085
rect 21542 34076 21548 34088
rect 21600 34076 21606 34128
rect 10042 34048 10048 34060
rect 9508 34020 10048 34048
rect 8389 33983 8447 33989
rect 8389 33949 8401 33983
rect 8435 33980 8447 33983
rect 9030 33980 9036 33992
rect 8435 33952 9036 33980
rect 8435 33949 8447 33952
rect 8389 33943 8447 33949
rect 9030 33940 9036 33952
rect 9088 33940 9094 33992
rect 9508 33989 9536 34020
rect 10042 34008 10048 34020
rect 10100 34008 10106 34060
rect 21652 34048 21680 34156
rect 26694 34144 26700 34156
rect 26752 34144 26758 34196
rect 34241 34187 34299 34193
rect 34241 34153 34253 34187
rect 34287 34184 34299 34187
rect 34790 34184 34796 34196
rect 34287 34156 34796 34184
rect 34287 34153 34299 34156
rect 34241 34147 34299 34153
rect 34790 34144 34796 34156
rect 34848 34144 34854 34196
rect 24029 34119 24087 34125
rect 13464 34020 16344 34048
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33949 9551 33983
rect 10134 33980 10140 33992
rect 10095 33952 10140 33980
rect 9493 33943 9551 33949
rect 10134 33940 10140 33952
rect 10192 33940 10198 33992
rect 10226 33940 10232 33992
rect 10284 33940 10290 33992
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33980 10839 33983
rect 10870 33980 10876 33992
rect 10827 33952 10876 33980
rect 10827 33949 10839 33952
rect 10781 33943 10839 33949
rect 10870 33940 10876 33952
rect 10928 33940 10934 33992
rect 11425 33983 11483 33989
rect 11425 33949 11437 33983
rect 11471 33980 11483 33983
rect 11790 33980 11796 33992
rect 11471 33952 11796 33980
rect 11471 33949 11483 33952
rect 11425 33943 11483 33949
rect 11790 33940 11796 33952
rect 11848 33940 11854 33992
rect 13464 33989 13492 34020
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 13814 33940 13820 33992
rect 13872 33980 13878 33992
rect 14553 33983 14611 33989
rect 14553 33980 14565 33983
rect 13872 33952 14565 33980
rect 13872 33940 13878 33952
rect 14553 33949 14565 33952
rect 14599 33949 14611 33983
rect 14553 33943 14611 33949
rect 9398 33872 9404 33924
rect 9456 33912 9462 33924
rect 10244 33912 10272 33940
rect 11974 33912 11980 33924
rect 9456 33884 11980 33912
rect 9456 33872 9462 33884
rect 11974 33872 11980 33884
rect 12032 33872 12038 33924
rect 12158 33912 12164 33924
rect 12119 33884 12164 33912
rect 12158 33872 12164 33884
rect 12216 33872 12222 33924
rect 12253 33915 12311 33921
rect 12253 33881 12265 33915
rect 12299 33881 12311 33915
rect 12802 33912 12808 33924
rect 12715 33884 12808 33912
rect 12253 33875 12311 33881
rect 3234 33804 3240 33856
rect 3292 33844 3298 33856
rect 8202 33844 8208 33856
rect 3292 33816 8208 33844
rect 3292 33804 3298 33816
rect 8202 33804 8208 33816
rect 8260 33804 8266 33856
rect 9582 33844 9588 33856
rect 9543 33816 9588 33844
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 9766 33804 9772 33856
rect 9824 33844 9830 33856
rect 10229 33847 10287 33853
rect 10229 33844 10241 33847
rect 9824 33816 10241 33844
rect 9824 33804 9830 33816
rect 10229 33813 10241 33816
rect 10275 33813 10287 33847
rect 10229 33807 10287 33813
rect 10318 33804 10324 33856
rect 10376 33844 10382 33856
rect 12268 33844 12296 33875
rect 12802 33872 12808 33884
rect 12860 33912 12866 33924
rect 12860 33884 13492 33912
rect 12860 33872 12866 33884
rect 10376 33816 12296 33844
rect 13464 33844 13492 33884
rect 13538 33872 13544 33924
rect 13596 33912 13602 33924
rect 15289 33915 15347 33921
rect 15289 33912 15301 33915
rect 13596 33884 15301 33912
rect 13596 33872 13602 33884
rect 15289 33881 15301 33884
rect 15335 33881 15347 33915
rect 15289 33875 15347 33881
rect 15378 33872 15384 33924
rect 15436 33912 15442 33924
rect 15933 33915 15991 33921
rect 15436 33884 15481 33912
rect 15436 33872 15442 33884
rect 15933 33881 15945 33915
rect 15979 33912 15991 33915
rect 16022 33912 16028 33924
rect 15979 33884 16028 33912
rect 15979 33881 15991 33884
rect 15933 33875 15991 33881
rect 15948 33844 15976 33875
rect 16022 33872 16028 33884
rect 16080 33872 16086 33924
rect 16316 33912 16344 34020
rect 16408 34020 21680 34048
rect 21836 34088 22094 34116
rect 16408 33989 16436 34020
rect 16393 33983 16451 33989
rect 16393 33949 16405 33983
rect 16439 33949 16451 33983
rect 16393 33943 16451 33949
rect 16482 33940 16488 33992
rect 16540 33980 16546 33992
rect 19518 33980 19524 33992
rect 16540 33952 19524 33980
rect 16540 33940 16546 33952
rect 19518 33940 19524 33952
rect 19576 33940 19582 33992
rect 19610 33940 19616 33992
rect 19668 33980 19674 33992
rect 21836 33980 21864 34088
rect 22066 34048 22094 34088
rect 24029 34085 24041 34119
rect 24075 34116 24087 34119
rect 25130 34116 25136 34128
rect 24075 34088 25136 34116
rect 24075 34085 24087 34088
rect 24029 34079 24087 34085
rect 24044 34048 24072 34079
rect 25130 34076 25136 34088
rect 25188 34076 25194 34128
rect 26602 34048 26608 34060
rect 22066 34020 24072 34048
rect 26563 34020 26608 34048
rect 26602 34008 26608 34020
rect 26660 34008 26666 34060
rect 26712 34048 26740 34144
rect 28184 34088 35894 34116
rect 26881 34051 26939 34057
rect 26881 34048 26893 34051
rect 26712 34020 26893 34048
rect 26881 34017 26893 34020
rect 26927 34017 26939 34051
rect 26881 34011 26939 34017
rect 19668 33952 21864 33980
rect 19668 33940 19674 33952
rect 22002 33940 22008 33992
rect 22060 33980 22066 33992
rect 22281 33983 22339 33989
rect 22281 33980 22293 33983
rect 22060 33952 22293 33980
rect 22060 33940 22066 33952
rect 22281 33949 22293 33952
rect 22327 33949 22339 33983
rect 22281 33943 22339 33949
rect 16316 33884 20116 33912
rect 13464 33816 15976 33844
rect 10376 33804 10382 33816
rect 17034 33804 17040 33856
rect 17092 33844 17098 33856
rect 19978 33844 19984 33856
rect 17092 33816 19984 33844
rect 17092 33804 17098 33816
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 20088 33844 20116 33884
rect 21450 33872 21456 33924
rect 21508 33912 21514 33924
rect 22557 33915 22615 33921
rect 22557 33912 22569 33915
rect 21508 33884 22569 33912
rect 21508 33872 21514 33884
rect 22557 33881 22569 33884
rect 22603 33881 22615 33915
rect 22557 33875 22615 33881
rect 23014 33872 23020 33924
rect 23072 33872 23078 33924
rect 24670 33872 24676 33924
rect 24728 33912 24734 33924
rect 25130 33912 25136 33924
rect 24728 33884 25136 33912
rect 24728 33872 24734 33884
rect 25130 33872 25136 33884
rect 25188 33912 25194 33924
rect 27154 33912 27160 33924
rect 25188 33884 27160 33912
rect 25188 33872 25194 33884
rect 27154 33872 27160 33884
rect 27212 33872 27218 33924
rect 27614 33872 27620 33924
rect 27672 33872 27678 33924
rect 24762 33844 24768 33856
rect 20088 33816 24768 33844
rect 24762 33804 24768 33816
rect 24820 33804 24826 33856
rect 24854 33804 24860 33856
rect 24912 33844 24918 33856
rect 28184 33844 28212 34088
rect 29730 34008 29736 34060
rect 29788 34048 29794 34060
rect 29788 34020 32812 34048
rect 29788 34008 29794 34020
rect 32784 33989 32812 34020
rect 34606 34008 34612 34060
rect 34664 34048 34670 34060
rect 34977 34051 35035 34057
rect 34977 34048 34989 34051
rect 34664 34020 34989 34048
rect 34664 34008 34670 34020
rect 34977 34017 34989 34020
rect 35023 34017 35035 34051
rect 35434 34048 35440 34060
rect 35395 34020 35440 34048
rect 34977 34011 35035 34017
rect 35434 34008 35440 34020
rect 35492 34008 35498 34060
rect 32769 33983 32827 33989
rect 32769 33949 32781 33983
rect 32815 33949 32827 33983
rect 34146 33980 34152 33992
rect 34107 33952 34152 33980
rect 32769 33943 32827 33949
rect 34146 33940 34152 33952
rect 34204 33940 34210 33992
rect 35866 33980 35894 34088
rect 36633 33983 36691 33989
rect 36633 33980 36645 33983
rect 35866 33952 36645 33980
rect 36633 33949 36645 33952
rect 36679 33949 36691 33983
rect 36633 33943 36691 33949
rect 31018 33872 31024 33924
rect 31076 33912 31082 33924
rect 31205 33915 31263 33921
rect 31205 33912 31217 33915
rect 31076 33884 31217 33912
rect 31076 33872 31082 33884
rect 31205 33881 31217 33884
rect 31251 33881 31263 33915
rect 31205 33875 31263 33881
rect 31297 33915 31355 33921
rect 31297 33881 31309 33915
rect 31343 33912 31355 33915
rect 31846 33912 31852 33924
rect 31343 33884 31754 33912
rect 31807 33884 31852 33912
rect 31343 33881 31355 33884
rect 31297 33875 31355 33881
rect 28350 33844 28356 33856
rect 24912 33816 28212 33844
rect 28311 33816 28356 33844
rect 24912 33804 24918 33816
rect 28350 33804 28356 33816
rect 28408 33804 28414 33856
rect 31726 33844 31754 33884
rect 31846 33872 31852 33884
rect 31904 33872 31910 33924
rect 32950 33872 32956 33924
rect 33008 33912 33014 33924
rect 33505 33915 33563 33921
rect 33505 33912 33517 33915
rect 33008 33884 33517 33912
rect 33008 33872 33014 33884
rect 33505 33881 33517 33884
rect 33551 33912 33563 33915
rect 34790 33912 34796 33924
rect 33551 33884 34796 33912
rect 33551 33881 33563 33884
rect 33505 33875 33563 33881
rect 34790 33872 34796 33884
rect 34848 33872 34854 33924
rect 35069 33915 35127 33921
rect 35069 33881 35081 33915
rect 35115 33881 35127 33915
rect 35069 33875 35127 33881
rect 32398 33844 32404 33856
rect 31726 33816 32404 33844
rect 32398 33804 32404 33816
rect 32456 33804 32462 33856
rect 33410 33804 33416 33856
rect 33468 33844 33474 33856
rect 35084 33844 35112 33875
rect 33468 33816 35112 33844
rect 33468 33804 33474 33816
rect 36354 33804 36360 33856
rect 36412 33844 36418 33856
rect 36725 33847 36783 33853
rect 36725 33844 36737 33847
rect 36412 33816 36737 33844
rect 36412 33804 36418 33816
rect 36725 33813 36737 33816
rect 36771 33813 36783 33847
rect 36725 33807 36783 33813
rect 36906 33804 36912 33856
rect 36964 33844 36970 33856
rect 37553 33847 37611 33853
rect 37553 33844 37565 33847
rect 36964 33816 37565 33844
rect 36964 33804 36970 33816
rect 37553 33813 37565 33816
rect 37599 33813 37611 33847
rect 37553 33807 37611 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 2498 33600 2504 33652
rect 2556 33640 2562 33652
rect 6825 33643 6883 33649
rect 6825 33640 6837 33643
rect 2556 33612 6837 33640
rect 2556 33600 2562 33612
rect 6825 33609 6837 33612
rect 6871 33609 6883 33643
rect 8570 33640 8576 33652
rect 8531 33612 8576 33640
rect 6825 33603 6883 33609
rect 8570 33600 8576 33612
rect 8628 33600 8634 33652
rect 9582 33600 9588 33652
rect 9640 33640 9646 33652
rect 15013 33643 15071 33649
rect 9640 33612 13952 33640
rect 9640 33600 9646 33612
rect 7466 33532 7472 33584
rect 7524 33572 7530 33584
rect 10318 33572 10324 33584
rect 7524 33544 9260 33572
rect 7524 33532 7530 33544
rect 6733 33507 6791 33513
rect 6733 33473 6745 33507
rect 6779 33504 6791 33507
rect 8294 33504 8300 33516
rect 6779 33476 8300 33504
rect 6779 33473 6791 33476
rect 6733 33467 6791 33473
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 8481 33507 8539 33513
rect 8481 33473 8493 33507
rect 8527 33473 8539 33507
rect 8481 33467 8539 33473
rect 8496 33368 8524 33467
rect 9232 33436 9260 33544
rect 9600 33544 10324 33572
rect 9398 33464 9404 33516
rect 9456 33504 9462 33516
rect 9600 33513 9628 33544
rect 10318 33532 10324 33544
rect 10376 33532 10382 33584
rect 10410 33532 10416 33584
rect 10468 33572 10474 33584
rect 11885 33575 11943 33581
rect 11885 33572 11897 33575
rect 10468 33544 11897 33572
rect 10468 33532 10474 33544
rect 11885 33541 11897 33544
rect 11931 33541 11943 33575
rect 11885 33535 11943 33541
rect 11974 33532 11980 33584
rect 12032 33572 12038 33584
rect 13924 33581 13952 33612
rect 15013 33609 15025 33643
rect 15059 33640 15071 33643
rect 16298 33640 16304 33652
rect 15059 33612 16304 33640
rect 15059 33609 15071 33612
rect 15013 33603 15071 33609
rect 16298 33600 16304 33612
rect 16356 33600 16362 33652
rect 16574 33600 16580 33652
rect 16632 33640 16638 33652
rect 17129 33643 17187 33649
rect 17129 33640 17141 33643
rect 16632 33612 17141 33640
rect 16632 33600 16638 33612
rect 17129 33609 17141 33612
rect 17175 33609 17187 33643
rect 17129 33603 17187 33609
rect 17236 33612 19748 33640
rect 13909 33575 13967 33581
rect 12032 33544 13124 33572
rect 12032 33532 12038 33544
rect 9493 33507 9551 33513
rect 9493 33504 9505 33507
rect 9456 33476 9505 33504
rect 9456 33464 9462 33476
rect 9493 33473 9505 33476
rect 9539 33473 9551 33507
rect 9493 33467 9551 33473
rect 9585 33507 9643 33513
rect 9585 33473 9597 33507
rect 9631 33473 9643 33507
rect 10134 33504 10140 33516
rect 10095 33476 10140 33504
rect 9585 33467 9643 33473
rect 10134 33464 10140 33476
rect 10192 33464 10198 33516
rect 10965 33507 11023 33513
rect 10965 33473 10977 33507
rect 11011 33504 11023 33507
rect 11054 33504 11060 33516
rect 11011 33476 11060 33504
rect 11011 33473 11023 33476
rect 10965 33467 11023 33473
rect 11054 33464 11060 33476
rect 11112 33464 11118 33516
rect 13096 33513 13124 33544
rect 13909 33541 13921 33575
rect 13955 33541 13967 33575
rect 14458 33572 14464 33584
rect 14419 33544 14464 33572
rect 13909 33535 13967 33541
rect 14458 33532 14464 33544
rect 14516 33532 14522 33584
rect 15657 33575 15715 33581
rect 15657 33541 15669 33575
rect 15703 33572 15715 33575
rect 16482 33572 16488 33584
rect 15703 33544 16488 33572
rect 15703 33541 15715 33544
rect 15657 33535 15715 33541
rect 16482 33532 16488 33544
rect 16540 33532 16546 33584
rect 13081 33507 13139 33513
rect 13081 33473 13093 33507
rect 13127 33473 13139 33507
rect 13081 33467 13139 33473
rect 14921 33507 14979 33513
rect 14921 33473 14933 33507
rect 14967 33504 14979 33507
rect 15010 33504 15016 33516
rect 14967 33476 15016 33504
rect 14967 33473 14979 33476
rect 14921 33467 14979 33473
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 15562 33504 15568 33516
rect 15523 33476 15568 33504
rect 15562 33464 15568 33476
rect 15620 33464 15626 33516
rect 17034 33504 17040 33516
rect 16995 33476 17040 33504
rect 17034 33464 17040 33476
rect 17092 33464 17098 33516
rect 11793 33439 11851 33445
rect 11793 33436 11805 33439
rect 9232 33408 11805 33436
rect 11793 33405 11805 33408
rect 11839 33405 11851 33439
rect 13814 33436 13820 33448
rect 11793 33399 11851 33405
rect 12268 33408 12664 33436
rect 13775 33408 13820 33436
rect 12268 33368 12296 33408
rect 8496 33340 12296 33368
rect 12345 33371 12403 33377
rect 12345 33337 12357 33371
rect 12391 33368 12403 33371
rect 12526 33368 12532 33380
rect 12391 33340 12532 33368
rect 12391 33337 12403 33340
rect 12345 33331 12403 33337
rect 12526 33328 12532 33340
rect 12584 33328 12590 33380
rect 12636 33368 12664 33408
rect 13814 33396 13820 33408
rect 13872 33396 13878 33448
rect 17236 33436 17264 33612
rect 19720 33504 19748 33612
rect 19978 33600 19984 33652
rect 20036 33640 20042 33652
rect 24670 33640 24676 33652
rect 20036 33612 24676 33640
rect 20036 33600 20042 33612
rect 24670 33600 24676 33612
rect 24728 33600 24734 33652
rect 24762 33600 24768 33652
rect 24820 33640 24826 33652
rect 31481 33643 31539 33649
rect 24820 33612 31432 33640
rect 24820 33600 24826 33612
rect 19794 33532 19800 33584
rect 19852 33572 19858 33584
rect 24854 33572 24860 33584
rect 19852 33544 24860 33572
rect 19852 33532 19858 33544
rect 24854 33532 24860 33544
rect 24912 33532 24918 33584
rect 25130 33532 25136 33584
rect 25188 33572 25194 33584
rect 25188 33544 25233 33572
rect 25188 33532 25194 33544
rect 25590 33532 25596 33584
rect 25648 33532 25654 33584
rect 31404 33513 31432 33612
rect 31481 33609 31493 33643
rect 31527 33640 31539 33643
rect 31570 33640 31576 33652
rect 31527 33612 31576 33640
rect 31527 33609 31539 33612
rect 31481 33603 31539 33609
rect 31570 33600 31576 33612
rect 31628 33600 31634 33652
rect 32398 33640 32404 33652
rect 32359 33612 32404 33640
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 35621 33643 35679 33649
rect 35621 33609 35633 33643
rect 35667 33640 35679 33643
rect 36446 33640 36452 33652
rect 35667 33612 36452 33640
rect 35667 33609 35679 33612
rect 35621 33603 35679 33609
rect 36446 33600 36452 33612
rect 36504 33600 36510 33652
rect 32858 33572 32864 33584
rect 32324 33544 32864 33572
rect 32324 33513 32352 33544
rect 32858 33532 32864 33544
rect 32916 33532 32922 33584
rect 34698 33572 34704 33584
rect 34454 33544 34704 33572
rect 34698 33532 34704 33544
rect 34756 33532 34762 33584
rect 31389 33507 31447 33513
rect 18138 33436 18144 33448
rect 14476 33408 17264 33436
rect 18099 33408 18144 33436
rect 14476 33368 14504 33408
rect 18138 33396 18144 33408
rect 18196 33396 18202 33448
rect 18417 33439 18475 33445
rect 18417 33405 18429 33439
rect 18463 33436 18475 33439
rect 18874 33436 18880 33448
rect 18463 33408 18880 33436
rect 18463 33405 18475 33408
rect 18417 33399 18475 33405
rect 18874 33396 18880 33408
rect 18932 33396 18938 33448
rect 18966 33396 18972 33448
rect 19024 33436 19030 33448
rect 19536 33436 19564 33490
rect 19720 33476 22094 33504
rect 20162 33436 20168 33448
rect 19024 33408 19472 33436
rect 19536 33408 20168 33436
rect 19024 33396 19030 33408
rect 12636 33340 14504 33368
rect 19444 33368 19472 33408
rect 20162 33396 20168 33408
rect 20220 33396 20226 33448
rect 19702 33368 19708 33380
rect 19444 33340 19708 33368
rect 19702 33328 19708 33340
rect 19760 33328 19766 33380
rect 19886 33368 19892 33380
rect 19847 33340 19892 33368
rect 19886 33328 19892 33340
rect 19944 33368 19950 33380
rect 20254 33368 20260 33380
rect 19944 33340 20260 33368
rect 19944 33328 19950 33340
rect 20254 33328 20260 33340
rect 20312 33328 20318 33380
rect 22066 33368 22094 33476
rect 31389 33473 31401 33507
rect 31435 33504 31447 33507
rect 32309 33507 32367 33513
rect 31435 33476 31754 33504
rect 31435 33473 31447 33476
rect 31389 33467 31447 33473
rect 24394 33396 24400 33448
rect 24452 33436 24458 33448
rect 24857 33439 24915 33445
rect 24857 33436 24869 33439
rect 24452 33408 24869 33436
rect 24452 33396 24458 33408
rect 24857 33405 24869 33408
rect 24903 33405 24915 33439
rect 26510 33436 26516 33448
rect 24857 33399 24915 33405
rect 24964 33408 26516 33436
rect 24964 33368 24992 33408
rect 26510 33396 26516 33408
rect 26568 33396 26574 33448
rect 22066 33340 24992 33368
rect 9858 33260 9864 33312
rect 9916 33300 9922 33312
rect 10229 33303 10287 33309
rect 10229 33300 10241 33303
rect 9916 33272 10241 33300
rect 9916 33260 9922 33272
rect 10229 33269 10241 33272
rect 10275 33269 10287 33303
rect 10229 33263 10287 33269
rect 11057 33303 11115 33309
rect 11057 33269 11069 33303
rect 11103 33300 11115 33303
rect 11974 33300 11980 33312
rect 11103 33272 11980 33300
rect 11103 33269 11115 33272
rect 11057 33263 11115 33269
rect 11974 33260 11980 33272
rect 12032 33260 12038 33312
rect 13173 33303 13231 33309
rect 13173 33269 13185 33303
rect 13219 33300 13231 33303
rect 13814 33300 13820 33312
rect 13219 33272 13820 33300
rect 13219 33269 13231 33272
rect 13173 33263 13231 33269
rect 13814 33260 13820 33272
rect 13872 33260 13878 33312
rect 17586 33260 17592 33312
rect 17644 33300 17650 33312
rect 26418 33300 26424 33312
rect 17644 33272 26424 33300
rect 17644 33260 17650 33272
rect 26418 33260 26424 33272
rect 26476 33260 26482 33312
rect 26602 33300 26608 33312
rect 26563 33272 26608 33300
rect 26602 33260 26608 33272
rect 26660 33260 26666 33312
rect 31726 33300 31754 33476
rect 32309 33473 32321 33507
rect 32355 33473 32367 33507
rect 32950 33504 32956 33516
rect 32911 33476 32956 33504
rect 32309 33467 32367 33473
rect 32950 33464 32956 33476
rect 33008 33464 33014 33516
rect 35526 33504 35532 33516
rect 35487 33476 35532 33504
rect 35526 33464 35532 33476
rect 35584 33464 35590 33516
rect 36354 33504 36360 33516
rect 36315 33476 36360 33504
rect 36354 33464 36360 33476
rect 36412 33464 36418 33516
rect 38102 33504 38108 33516
rect 38063 33476 38108 33504
rect 38102 33464 38108 33476
rect 38160 33464 38166 33516
rect 33229 33439 33287 33445
rect 33229 33436 33241 33439
rect 32324 33408 33241 33436
rect 32324 33380 32352 33408
rect 33229 33405 33241 33408
rect 33275 33405 33287 33439
rect 33229 33399 33287 33405
rect 34514 33396 34520 33448
rect 34572 33396 34578 33448
rect 32306 33328 32312 33380
rect 32364 33328 32370 33380
rect 34532 33368 34560 33396
rect 34256 33340 34560 33368
rect 38289 33371 38347 33377
rect 34256 33300 34284 33340
rect 38289 33337 38301 33371
rect 38335 33368 38347 33371
rect 38838 33368 38844 33380
rect 38335 33340 38844 33368
rect 38335 33337 38347 33340
rect 38289 33331 38347 33337
rect 38838 33328 38844 33340
rect 38896 33328 38902 33380
rect 31726 33272 34284 33300
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 34701 33303 34759 33309
rect 34701 33300 34713 33303
rect 34572 33272 34713 33300
rect 34572 33260 34578 33272
rect 34701 33269 34713 33272
rect 34747 33269 34759 33303
rect 34701 33263 34759 33269
rect 36173 33303 36231 33309
rect 36173 33269 36185 33303
rect 36219 33300 36231 33303
rect 38010 33300 38016 33312
rect 36219 33272 38016 33300
rect 36219 33269 36231 33272
rect 36173 33263 36231 33269
rect 38010 33260 38016 33272
rect 38068 33260 38074 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 12158 33096 12164 33108
rect 9232 33068 12164 33096
rect 1581 32895 1639 32901
rect 1581 32861 1593 32895
rect 1627 32892 1639 32895
rect 2958 32892 2964 32904
rect 1627 32864 2964 32892
rect 1627 32861 1639 32864
rect 1581 32855 1639 32861
rect 2958 32852 2964 32864
rect 3016 32852 3022 32904
rect 5718 32852 5724 32904
rect 5776 32892 5782 32904
rect 9232 32901 9260 33068
rect 12158 33056 12164 33068
rect 12216 33056 12222 33108
rect 12250 33056 12256 33108
rect 12308 33096 12314 33108
rect 15102 33096 15108 33108
rect 12308 33068 15108 33096
rect 12308 33056 12314 33068
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 15194 33056 15200 33108
rect 15252 33096 15258 33108
rect 15252 33068 20760 33096
rect 15252 33056 15258 33068
rect 10597 33031 10655 33037
rect 10597 32997 10609 33031
rect 10643 33028 10655 33031
rect 10962 33028 10968 33040
rect 10643 33000 10968 33028
rect 10643 32997 10655 33000
rect 10597 32991 10655 32997
rect 10962 32988 10968 33000
rect 11020 32988 11026 33040
rect 13998 33028 14004 33040
rect 11164 33000 14004 33028
rect 7193 32895 7251 32901
rect 7193 32892 7205 32895
rect 5776 32864 7205 32892
rect 5776 32852 5782 32864
rect 7193 32861 7205 32864
rect 7239 32861 7251 32895
rect 7193 32855 7251 32861
rect 8573 32895 8631 32901
rect 8573 32861 8585 32895
rect 8619 32861 8631 32895
rect 8573 32855 8631 32861
rect 9217 32895 9275 32901
rect 9217 32861 9229 32895
rect 9263 32861 9275 32895
rect 9217 32855 9275 32861
rect 7558 32784 7564 32836
rect 7616 32824 7622 32836
rect 8588 32824 8616 32855
rect 9674 32852 9680 32904
rect 9732 32892 9738 32904
rect 9861 32895 9919 32901
rect 9861 32892 9873 32895
rect 9732 32864 9873 32892
rect 9732 32852 9738 32864
rect 9861 32861 9873 32864
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 10505 32895 10563 32901
rect 10505 32861 10517 32895
rect 10551 32892 10563 32895
rect 10594 32892 10600 32904
rect 10551 32864 10600 32892
rect 10551 32861 10563 32864
rect 10505 32855 10563 32861
rect 10594 32852 10600 32864
rect 10652 32852 10658 32904
rect 11164 32901 11192 33000
rect 13998 32988 14004 33000
rect 14056 32988 14062 33040
rect 14918 32988 14924 33040
rect 14976 33028 14982 33040
rect 20732 33028 20760 33068
rect 20806 33056 20812 33108
rect 20864 33096 20870 33108
rect 21177 33099 21235 33105
rect 21177 33096 21189 33099
rect 20864 33068 21189 33096
rect 20864 33056 20870 33068
rect 21177 33065 21189 33068
rect 21223 33096 21235 33099
rect 21358 33096 21364 33108
rect 21223 33068 21364 33096
rect 21223 33065 21235 33068
rect 21177 33059 21235 33065
rect 21358 33056 21364 33068
rect 21416 33056 21422 33108
rect 22922 33056 22928 33108
rect 22980 33096 22986 33108
rect 34241 33099 34299 33105
rect 22980 33068 30880 33096
rect 22980 33056 22986 33068
rect 24486 33028 24492 33040
rect 14976 33000 19564 33028
rect 20732 33000 24492 33028
rect 14976 32988 14982 33000
rect 11514 32920 11520 32972
rect 11572 32960 11578 32972
rect 12161 32963 12219 32969
rect 12161 32960 12173 32963
rect 11572 32932 12173 32960
rect 11572 32920 11578 32932
rect 12161 32929 12173 32932
rect 12207 32929 12219 32963
rect 12161 32923 12219 32929
rect 15194 32920 15200 32972
rect 15252 32960 15258 32972
rect 16025 32963 16083 32969
rect 16025 32960 16037 32963
rect 15252 32932 16037 32960
rect 15252 32920 15258 32932
rect 16025 32929 16037 32932
rect 16071 32960 16083 32963
rect 17034 32960 17040 32972
rect 16071 32932 17040 32960
rect 16071 32929 16083 32932
rect 16025 32923 16083 32929
rect 17034 32920 17040 32932
rect 17092 32920 17098 32972
rect 17221 32963 17279 32969
rect 17221 32929 17233 32963
rect 17267 32960 17279 32963
rect 17494 32960 17500 32972
rect 17267 32932 17500 32960
rect 17267 32929 17279 32932
rect 17221 32923 17279 32929
rect 17494 32920 17500 32932
rect 17552 32920 17558 32972
rect 19426 32960 19432 32972
rect 19387 32932 19432 32960
rect 19426 32920 19432 32932
rect 19484 32920 19490 32972
rect 19536 32960 19564 33000
rect 24486 32988 24492 33000
rect 24544 32988 24550 33040
rect 19536 32932 22094 32960
rect 11149 32895 11207 32901
rect 11149 32861 11161 32895
rect 11195 32861 11207 32895
rect 11149 32855 11207 32861
rect 13262 32852 13268 32904
rect 13320 32892 13326 32904
rect 13541 32895 13599 32901
rect 13541 32892 13553 32895
rect 13320 32864 13553 32892
rect 13320 32852 13326 32864
rect 13541 32861 13553 32864
rect 13587 32892 13599 32895
rect 14369 32895 14427 32901
rect 14369 32892 14381 32895
rect 13587 32864 14381 32892
rect 13587 32861 13599 32864
rect 13541 32855 13599 32861
rect 14369 32861 14381 32864
rect 14415 32861 14427 32895
rect 15010 32892 15016 32904
rect 14971 32864 15016 32892
rect 14369 32855 14427 32861
rect 15010 32852 15016 32864
rect 15068 32852 15074 32904
rect 17129 32895 17187 32901
rect 17129 32861 17141 32895
rect 17175 32886 17187 32895
rect 18414 32892 18420 32904
rect 17328 32886 18420 32892
rect 17175 32864 18420 32886
rect 17175 32861 17356 32864
rect 17129 32858 17356 32861
rect 17129 32855 17187 32858
rect 18414 32852 18420 32864
rect 18472 32852 18478 32904
rect 22066 32892 22094 32932
rect 22738 32920 22744 32972
rect 22796 32960 22802 32972
rect 24857 32963 24915 32969
rect 24857 32960 24869 32963
rect 22796 32932 24869 32960
rect 22796 32920 22802 32932
rect 24857 32929 24869 32932
rect 24903 32960 24915 32963
rect 26602 32960 26608 32972
rect 24903 32932 26608 32960
rect 24903 32929 24915 32932
rect 24857 32923 24915 32929
rect 26602 32920 26608 32932
rect 26660 32920 26666 32972
rect 30558 32920 30564 32972
rect 30616 32960 30622 32972
rect 30745 32963 30803 32969
rect 30745 32960 30757 32963
rect 30616 32932 30757 32960
rect 30616 32920 30622 32932
rect 30745 32929 30757 32932
rect 30791 32929 30803 32963
rect 30852 32960 30880 33068
rect 34241 33065 34253 33099
rect 34287 33096 34299 33099
rect 34606 33096 34612 33108
rect 34287 33068 34612 33096
rect 34287 33065 34299 33068
rect 34241 33059 34299 33065
rect 34606 33056 34612 33068
rect 34664 33056 34670 33108
rect 36633 33099 36691 33105
rect 36633 33096 36645 33099
rect 34716 33068 36645 33096
rect 34146 32988 34152 33040
rect 34204 33028 34210 33040
rect 34716 33028 34744 33068
rect 36633 33065 36645 33068
rect 36679 33065 36691 33099
rect 36633 33059 36691 33065
rect 37461 33099 37519 33105
rect 37461 33065 37473 33099
rect 37507 33096 37519 33099
rect 37550 33096 37556 33108
rect 37507 33068 37556 33096
rect 37507 33065 37519 33068
rect 37461 33059 37519 33065
rect 37550 33056 37556 33068
rect 37608 33056 37614 33108
rect 34204 33000 34744 33028
rect 34204 32988 34210 33000
rect 33962 32960 33968 32972
rect 30852 32932 33968 32960
rect 30745 32923 30803 32929
rect 33962 32920 33968 32932
rect 34020 32960 34026 32972
rect 34020 32932 34192 32960
rect 34020 32920 34026 32932
rect 23750 32892 23756 32904
rect 22066 32864 23756 32892
rect 23750 32852 23756 32864
rect 23808 32852 23814 32904
rect 24394 32852 24400 32904
rect 24452 32892 24458 32904
rect 34164 32901 34192 32932
rect 34790 32920 34796 32972
rect 34848 32960 34854 32972
rect 34885 32963 34943 32969
rect 34885 32960 34897 32963
rect 34848 32932 34897 32960
rect 34848 32920 34854 32932
rect 34885 32929 34897 32932
rect 34931 32929 34943 32963
rect 34885 32923 34943 32929
rect 24581 32895 24639 32901
rect 24581 32892 24593 32895
rect 24452 32864 24593 32892
rect 24452 32852 24458 32864
rect 24581 32861 24593 32864
rect 24627 32861 24639 32895
rect 24581 32855 24639 32861
rect 34149 32895 34207 32901
rect 34149 32861 34161 32895
rect 34195 32861 34207 32895
rect 34149 32855 34207 32861
rect 37369 32895 37427 32901
rect 37369 32861 37381 32895
rect 37415 32892 37427 32895
rect 37826 32892 37832 32904
rect 37415 32864 37832 32892
rect 37415 32861 37427 32864
rect 37369 32855 37427 32861
rect 37826 32852 37832 32864
rect 37884 32852 37890 32904
rect 38010 32892 38016 32904
rect 37971 32864 38016 32892
rect 38010 32852 38016 32864
rect 38068 32852 38074 32904
rect 9766 32824 9772 32836
rect 7616 32796 8524 32824
rect 8588 32796 9772 32824
rect 7616 32784 7622 32796
rect 1762 32756 1768 32768
rect 1723 32728 1768 32756
rect 1762 32716 1768 32728
rect 1820 32716 1826 32768
rect 7282 32756 7288 32768
rect 7243 32728 7288 32756
rect 7282 32716 7288 32728
rect 7340 32716 7346 32768
rect 8386 32756 8392 32768
rect 8347 32728 8392 32756
rect 8386 32716 8392 32728
rect 8444 32716 8450 32768
rect 8496 32756 8524 32796
rect 9766 32784 9772 32796
rect 9824 32784 9830 32836
rect 9953 32827 10011 32833
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 11885 32827 11943 32833
rect 11885 32824 11897 32827
rect 9999 32796 11897 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 11885 32793 11897 32796
rect 11931 32793 11943 32827
rect 11885 32787 11943 32793
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 12032 32796 12077 32824
rect 12032 32784 12038 32796
rect 12158 32784 12164 32836
rect 12216 32824 12222 32836
rect 14458 32824 14464 32836
rect 12216 32796 14320 32824
rect 14419 32796 14464 32824
rect 12216 32784 12222 32796
rect 9309 32759 9367 32765
rect 9309 32756 9321 32759
rect 8496 32728 9321 32756
rect 9309 32725 9321 32728
rect 9355 32725 9367 32759
rect 9309 32719 9367 32725
rect 11241 32759 11299 32765
rect 11241 32725 11253 32759
rect 11287 32756 11299 32759
rect 12250 32756 12256 32768
rect 11287 32728 12256 32756
rect 11287 32725 11299 32728
rect 11241 32719 11299 32725
rect 12250 32716 12256 32728
rect 12308 32716 12314 32768
rect 13630 32756 13636 32768
rect 13591 32728 13636 32756
rect 13630 32716 13636 32728
rect 13688 32716 13694 32768
rect 14292 32756 14320 32796
rect 14458 32784 14464 32796
rect 14516 32784 14522 32836
rect 15838 32824 15844 32836
rect 14752 32796 15844 32824
rect 14752 32768 14780 32796
rect 15838 32784 15844 32796
rect 15896 32784 15902 32836
rect 16114 32784 16120 32836
rect 16172 32824 16178 32836
rect 16669 32827 16727 32833
rect 16172 32796 16217 32824
rect 16172 32784 16178 32796
rect 16669 32793 16681 32827
rect 16715 32824 16727 32827
rect 16758 32824 16764 32836
rect 16715 32796 16764 32824
rect 16715 32793 16727 32796
rect 16669 32787 16727 32793
rect 16758 32784 16764 32796
rect 16816 32784 16822 32836
rect 16850 32784 16856 32836
rect 16908 32824 16914 32836
rect 16908 32796 19380 32824
rect 16908 32784 16914 32796
rect 14734 32756 14740 32768
rect 14292 32728 14740 32756
rect 14734 32716 14740 32728
rect 14792 32716 14798 32768
rect 15105 32759 15163 32765
rect 15105 32725 15117 32759
rect 15151 32756 15163 32759
rect 18966 32756 18972 32768
rect 15151 32728 18972 32756
rect 15151 32725 15163 32728
rect 15105 32719 15163 32725
rect 18966 32716 18972 32728
rect 19024 32716 19030 32768
rect 19352 32756 19380 32796
rect 19426 32784 19432 32836
rect 19484 32824 19490 32836
rect 19705 32827 19763 32833
rect 19705 32824 19717 32827
rect 19484 32796 19717 32824
rect 19484 32784 19490 32796
rect 19705 32793 19717 32796
rect 19751 32793 19763 32827
rect 19705 32787 19763 32793
rect 20714 32784 20720 32836
rect 20772 32784 20778 32836
rect 22646 32784 22652 32836
rect 22704 32824 22710 32836
rect 24302 32824 24308 32836
rect 22704 32796 24308 32824
rect 22704 32784 22710 32796
rect 24302 32784 24308 32796
rect 24360 32784 24366 32836
rect 25498 32784 25504 32836
rect 25556 32784 25562 32836
rect 30650 32784 30656 32836
rect 30708 32824 30714 32836
rect 31021 32827 31079 32833
rect 31021 32824 31033 32827
rect 30708 32796 31033 32824
rect 30708 32784 30714 32796
rect 31021 32793 31033 32796
rect 31067 32793 31079 32827
rect 31021 32787 31079 32793
rect 31662 32784 31668 32836
rect 31720 32784 31726 32836
rect 33134 32784 33140 32836
rect 33192 32824 33198 32836
rect 35161 32827 35219 32833
rect 35161 32824 35173 32827
rect 33192 32796 35173 32824
rect 33192 32784 33198 32796
rect 35161 32793 35173 32796
rect 35207 32793 35219 32827
rect 38562 32824 38568 32836
rect 36386 32796 38568 32824
rect 35161 32787 35219 32793
rect 38562 32784 38568 32796
rect 38620 32784 38626 32836
rect 20438 32756 20444 32768
rect 19352 32728 20444 32756
rect 20438 32716 20444 32728
rect 20496 32716 20502 32768
rect 23934 32716 23940 32768
rect 23992 32756 23998 32768
rect 26329 32759 26387 32765
rect 26329 32756 26341 32759
rect 23992 32728 26341 32756
rect 23992 32716 23998 32728
rect 26329 32725 26341 32728
rect 26375 32725 26387 32759
rect 26329 32719 26387 32725
rect 32306 32716 32312 32768
rect 32364 32756 32370 32768
rect 32493 32759 32551 32765
rect 32493 32756 32505 32759
rect 32364 32728 32505 32756
rect 32364 32716 32370 32728
rect 32493 32725 32505 32728
rect 32539 32725 32551 32759
rect 38194 32756 38200 32768
rect 38155 32728 38200 32756
rect 32493 32719 32551 32725
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 10796 32524 12020 32552
rect 9858 32484 9864 32496
rect 9819 32456 9864 32484
rect 9858 32444 9864 32456
rect 9916 32444 9922 32496
rect 10796 32493 10824 32524
rect 10781 32487 10839 32493
rect 10781 32453 10793 32487
rect 10827 32453 10839 32487
rect 11885 32487 11943 32493
rect 11885 32484 11897 32487
rect 10781 32447 10839 32453
rect 10888 32456 11897 32484
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 5902 32416 5908 32428
rect 1627 32388 5908 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 5902 32376 5908 32388
rect 5960 32376 5966 32428
rect 9214 32416 9220 32428
rect 9175 32388 9220 32416
rect 9214 32376 9220 32388
rect 9272 32376 9278 32428
rect 9766 32348 9772 32360
rect 9727 32320 9772 32348
rect 9766 32308 9772 32320
rect 9824 32308 9830 32360
rect 9033 32283 9091 32289
rect 9033 32249 9045 32283
rect 9079 32280 9091 32283
rect 10888 32280 10916 32456
rect 11885 32453 11897 32456
rect 11931 32453 11943 32487
rect 11992 32484 12020 32524
rect 12526 32512 12532 32564
rect 12584 32552 12590 32564
rect 15013 32555 15071 32561
rect 12584 32524 14964 32552
rect 12584 32512 12590 32524
rect 13354 32484 13360 32496
rect 11992 32456 13360 32484
rect 11885 32447 11943 32453
rect 13354 32444 13360 32456
rect 13412 32444 13418 32496
rect 14936 32484 14964 32524
rect 15013 32521 15025 32555
rect 15059 32552 15071 32555
rect 16114 32552 16120 32564
rect 15059 32524 16120 32552
rect 15059 32521 15071 32524
rect 15013 32515 15071 32521
rect 16114 32512 16120 32524
rect 16172 32512 16178 32564
rect 17862 32512 17868 32564
rect 17920 32552 17926 32564
rect 17920 32524 18828 32552
rect 17920 32512 17926 32524
rect 13832 32456 14136 32484
rect 14936 32456 15056 32484
rect 12897 32419 12955 32425
rect 12897 32385 12909 32419
rect 12943 32416 12955 32419
rect 13538 32416 13544 32428
rect 12943 32388 13544 32416
rect 12943 32385 12955 32388
rect 12897 32379 12955 32385
rect 13538 32376 13544 32388
rect 13596 32376 13602 32428
rect 11790 32348 11796 32360
rect 11751 32320 11796 32348
rect 11790 32308 11796 32320
rect 11848 32308 11854 32360
rect 13832 32348 13860 32456
rect 13998 32416 14004 32428
rect 13959 32388 14004 32416
rect 13998 32376 14004 32388
rect 14056 32376 14062 32428
rect 14108 32416 14136 32456
rect 14918 32416 14924 32428
rect 14108 32388 14924 32416
rect 14918 32376 14924 32388
rect 14976 32376 14982 32428
rect 15028 32416 15056 32456
rect 15470 32444 15476 32496
rect 15528 32484 15534 32496
rect 15749 32487 15807 32493
rect 15749 32484 15761 32487
rect 15528 32456 15761 32484
rect 15528 32444 15534 32456
rect 15749 32453 15761 32456
rect 15795 32453 15807 32487
rect 15749 32447 15807 32453
rect 16022 32444 16028 32496
rect 16080 32484 16086 32496
rect 17402 32484 17408 32496
rect 16080 32456 17408 32484
rect 16080 32444 16086 32456
rect 17402 32444 17408 32456
rect 17460 32444 17466 32496
rect 18800 32484 18828 32524
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 19610 32552 19616 32564
rect 19392 32524 19616 32552
rect 19392 32512 19398 32524
rect 19610 32512 19616 32524
rect 19668 32512 19674 32564
rect 22646 32552 22652 32564
rect 19904 32524 22652 32552
rect 18800 32456 19090 32484
rect 15028 32388 15516 32416
rect 11992 32320 13860 32348
rect 14093 32351 14151 32357
rect 9079 32252 10916 32280
rect 9079 32249 9091 32252
rect 9033 32243 9091 32249
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 8662 32172 8668 32224
rect 8720 32212 8726 32224
rect 11992 32212 12020 32320
rect 14093 32317 14105 32351
rect 14139 32317 14151 32351
rect 15488 32348 15516 32388
rect 15657 32351 15715 32357
rect 15657 32348 15669 32351
rect 15488 32320 15669 32348
rect 14093 32311 14151 32317
rect 15657 32317 15669 32320
rect 15703 32317 15715 32351
rect 15657 32311 15715 32317
rect 12342 32280 12348 32292
rect 12303 32252 12348 32280
rect 12342 32240 12348 32252
rect 12400 32240 12406 32292
rect 14108 32280 14136 32311
rect 15838 32308 15844 32360
rect 15896 32348 15902 32360
rect 15933 32351 15991 32357
rect 15933 32348 15945 32351
rect 15896 32320 15945 32348
rect 15896 32308 15902 32320
rect 15933 32317 15945 32320
rect 15979 32317 15991 32351
rect 17954 32348 17960 32360
rect 15933 32311 15991 32317
rect 16132 32320 17960 32348
rect 16132 32280 16160 32320
rect 17954 32308 17960 32320
rect 18012 32308 18018 32360
rect 18230 32308 18236 32360
rect 18288 32348 18294 32360
rect 18325 32351 18383 32357
rect 18325 32348 18337 32351
rect 18288 32320 18337 32348
rect 18288 32308 18294 32320
rect 18325 32317 18337 32320
rect 18371 32317 18383 32351
rect 18325 32311 18383 32317
rect 18601 32351 18659 32357
rect 18601 32317 18613 32351
rect 18647 32348 18659 32351
rect 18690 32348 18696 32360
rect 18647 32320 18696 32348
rect 18647 32317 18659 32320
rect 18601 32311 18659 32317
rect 18690 32308 18696 32320
rect 18748 32308 18754 32360
rect 12636 32252 13124 32280
rect 14108 32252 16160 32280
rect 8720 32184 12020 32212
rect 8720 32172 8726 32184
rect 12250 32172 12256 32224
rect 12308 32212 12314 32224
rect 12636 32212 12664 32252
rect 12308 32184 12664 32212
rect 12308 32172 12314 32184
rect 12710 32172 12716 32224
rect 12768 32212 12774 32224
rect 12989 32215 13047 32221
rect 12989 32212 13001 32215
rect 12768 32184 13001 32212
rect 12768 32172 12774 32184
rect 12989 32181 13001 32184
rect 13035 32181 13047 32215
rect 13096 32212 13124 32252
rect 19904 32212 19932 32524
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 22833 32555 22891 32561
rect 22833 32521 22845 32555
rect 22879 32552 22891 32555
rect 24118 32552 24124 32564
rect 22879 32524 24124 32552
rect 22879 32521 22891 32524
rect 22833 32515 22891 32521
rect 24118 32512 24124 32524
rect 24176 32512 24182 32564
rect 29362 32552 29368 32564
rect 24412 32524 29368 32552
rect 20254 32444 20260 32496
rect 20312 32484 20318 32496
rect 23934 32484 23940 32496
rect 20312 32456 23940 32484
rect 20312 32444 20318 32456
rect 23934 32444 23940 32456
rect 23992 32444 23998 32496
rect 24029 32487 24087 32493
rect 24029 32453 24041 32487
rect 24075 32484 24087 32487
rect 24302 32484 24308 32496
rect 24075 32456 24308 32484
rect 24075 32453 24087 32456
rect 24029 32447 24087 32453
rect 24302 32444 24308 32456
rect 24360 32484 24366 32496
rect 24412 32484 24440 32524
rect 29362 32512 29368 32524
rect 29420 32512 29426 32564
rect 32769 32555 32827 32561
rect 32769 32521 32781 32555
rect 32815 32552 32827 32555
rect 33410 32552 33416 32564
rect 32815 32524 33416 32552
rect 32815 32521 32827 32524
rect 32769 32515 32827 32521
rect 33410 32512 33416 32524
rect 33468 32512 33474 32564
rect 36722 32552 36728 32564
rect 35176 32524 36728 32552
rect 24360 32456 24453 32484
rect 24360 32444 24366 32456
rect 24486 32444 24492 32496
rect 24544 32444 24550 32496
rect 34238 32444 34244 32496
rect 34296 32484 34302 32496
rect 35176 32493 35204 32524
rect 36722 32512 36728 32524
rect 36780 32512 36786 32564
rect 35161 32487 35219 32493
rect 35161 32484 35173 32487
rect 34296 32456 35173 32484
rect 34296 32444 34302 32456
rect 35161 32453 35173 32456
rect 35207 32453 35219 32487
rect 35161 32447 35219 32453
rect 20346 32416 20352 32428
rect 20259 32388 20352 32416
rect 20346 32376 20352 32388
rect 20404 32416 20410 32428
rect 22278 32416 22284 32428
rect 20404 32388 22284 32416
rect 20404 32376 20410 32388
rect 22278 32376 22284 32388
rect 22336 32376 22342 32428
rect 22738 32416 22744 32428
rect 22699 32388 22744 32416
rect 22738 32376 22744 32388
rect 22796 32376 22802 32428
rect 23750 32416 23756 32428
rect 23711 32388 23756 32416
rect 23750 32376 23756 32388
rect 23808 32376 23814 32428
rect 27525 32419 27583 32425
rect 27525 32416 27537 32419
rect 25240 32388 27537 32416
rect 20438 32308 20444 32360
rect 20496 32348 20502 32360
rect 25240 32348 25268 32388
rect 27525 32385 27537 32388
rect 27571 32385 27583 32419
rect 27525 32379 27583 32385
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 32677 32419 32735 32425
rect 32677 32416 32689 32419
rect 31812 32388 32689 32416
rect 31812 32376 31818 32388
rect 32677 32385 32689 32388
rect 32723 32385 32735 32419
rect 32677 32379 32735 32385
rect 34790 32376 34796 32428
rect 34848 32416 34854 32428
rect 34885 32419 34943 32425
rect 34885 32416 34897 32419
rect 34848 32388 34897 32416
rect 34848 32376 34854 32388
rect 34885 32385 34897 32388
rect 34931 32385 34943 32419
rect 34885 32379 34943 32385
rect 36262 32376 36268 32428
rect 36320 32376 36326 32428
rect 36814 32376 36820 32428
rect 36872 32416 36878 32428
rect 37645 32419 37703 32425
rect 37645 32416 37657 32419
rect 36872 32388 37657 32416
rect 36872 32376 36878 32388
rect 37645 32385 37657 32388
rect 37691 32385 37703 32419
rect 37645 32379 37703 32385
rect 25774 32348 25780 32360
rect 20496 32320 25268 32348
rect 25735 32320 25780 32348
rect 20496 32308 20502 32320
rect 25774 32308 25780 32320
rect 25832 32308 25838 32360
rect 35894 32308 35900 32360
rect 35952 32348 35958 32360
rect 35952 32320 36216 32348
rect 35952 32308 35958 32320
rect 21266 32240 21272 32292
rect 21324 32280 21330 32292
rect 23658 32280 23664 32292
rect 21324 32252 23664 32280
rect 21324 32240 21330 32252
rect 23658 32240 23664 32252
rect 23716 32240 23722 32292
rect 36188 32280 36216 32320
rect 36446 32308 36452 32360
rect 36504 32348 36510 32360
rect 36909 32351 36967 32357
rect 36909 32348 36921 32351
rect 36504 32320 36921 32348
rect 36504 32308 36510 32320
rect 36909 32317 36921 32320
rect 36955 32317 36967 32351
rect 36909 32311 36967 32317
rect 37461 32351 37519 32357
rect 37461 32317 37473 32351
rect 37507 32317 37519 32351
rect 37461 32311 37519 32317
rect 37476 32280 37504 32311
rect 36188 32252 37504 32280
rect 13096 32184 19932 32212
rect 12989 32175 13047 32181
rect 19978 32172 19984 32224
rect 20036 32212 20042 32224
rect 21910 32212 21916 32224
rect 20036 32184 21916 32212
rect 20036 32172 20042 32184
rect 21910 32172 21916 32184
rect 21968 32172 21974 32224
rect 23750 32172 23756 32224
rect 23808 32212 23814 32224
rect 24394 32212 24400 32224
rect 23808 32184 24400 32212
rect 23808 32172 23814 32184
rect 24394 32172 24400 32184
rect 24452 32172 24458 32224
rect 24578 32172 24584 32224
rect 24636 32212 24642 32224
rect 25314 32212 25320 32224
rect 24636 32184 25320 32212
rect 24636 32172 24642 32184
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 27338 32212 27344 32224
rect 27299 32184 27344 32212
rect 27338 32172 27344 32184
rect 27396 32172 27402 32224
rect 37826 32212 37832 32224
rect 37787 32184 37832 32212
rect 37826 32172 37832 32184
rect 37884 32172 37890 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 9401 32011 9459 32017
rect 9401 31977 9413 32011
rect 9447 32008 9459 32011
rect 9766 32008 9772 32020
rect 9447 31980 9772 32008
rect 9447 31977 9459 31980
rect 9401 31971 9459 31977
rect 9766 31968 9772 31980
rect 9824 31968 9830 32020
rect 11330 31968 11336 32020
rect 11388 32008 11394 32020
rect 15105 32011 15163 32017
rect 11388 31980 15056 32008
rect 11388 31968 11394 31980
rect 6549 31943 6607 31949
rect 6549 31909 6561 31943
rect 6595 31909 6607 31943
rect 6549 31903 6607 31909
rect 7745 31943 7803 31949
rect 7745 31909 7757 31943
rect 7791 31940 7803 31943
rect 8938 31940 8944 31952
rect 7791 31912 8944 31940
rect 7791 31909 7803 31912
rect 7745 31903 7803 31909
rect 6564 31872 6592 31903
rect 8938 31900 8944 31912
rect 8996 31900 9002 31952
rect 12250 31940 12256 31952
rect 9968 31912 12256 31940
rect 6564 31844 8524 31872
rect 6733 31807 6791 31813
rect 6733 31773 6745 31807
rect 6779 31804 6791 31807
rect 6822 31804 6828 31816
rect 6779 31776 6828 31804
rect 6779 31773 6791 31776
rect 6733 31767 6791 31773
rect 6822 31764 6828 31776
rect 6880 31764 6886 31816
rect 6914 31764 6920 31816
rect 6972 31804 6978 31816
rect 8496 31813 8524 31844
rect 7653 31807 7711 31813
rect 7653 31804 7665 31807
rect 6972 31776 7665 31804
rect 6972 31764 6978 31776
rect 7653 31773 7665 31776
rect 7699 31773 7711 31807
rect 7653 31767 7711 31773
rect 8481 31807 8539 31813
rect 8481 31773 8493 31807
rect 8527 31773 8539 31807
rect 8481 31767 8539 31773
rect 9122 31764 9128 31816
rect 9180 31804 9186 31816
rect 9968 31813 9996 31912
rect 12250 31900 12256 31912
rect 12308 31900 12314 31952
rect 13633 31943 13691 31949
rect 13633 31909 13645 31943
rect 13679 31940 13691 31943
rect 14918 31940 14924 31952
rect 13679 31912 14924 31940
rect 13679 31909 13691 31912
rect 13633 31903 13691 31909
rect 14918 31900 14924 31912
rect 14976 31900 14982 31952
rect 15028 31940 15056 31980
rect 15105 31977 15117 32011
rect 15151 32008 15163 32011
rect 15378 32008 15384 32020
rect 15151 31980 15384 32008
rect 15151 31977 15163 31980
rect 15105 31971 15163 31977
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 15746 32008 15752 32020
rect 15488 31980 15752 32008
rect 15488 31940 15516 31980
rect 15746 31968 15752 31980
rect 15804 31968 15810 32020
rect 15838 31968 15844 32020
rect 15896 32008 15902 32020
rect 16390 32008 16396 32020
rect 15896 31980 16396 32008
rect 15896 31968 15902 31980
rect 16390 31968 16396 31980
rect 16448 31968 16454 32020
rect 16942 31968 16948 32020
rect 17000 32008 17006 32020
rect 17037 32011 17095 32017
rect 17037 32008 17049 32011
rect 17000 31980 17049 32008
rect 17000 31968 17006 31980
rect 17037 31977 17049 31980
rect 17083 32008 17095 32011
rect 17586 32008 17592 32020
rect 17083 31980 17592 32008
rect 17083 31977 17095 31980
rect 17037 31971 17095 31977
rect 17586 31968 17592 31980
rect 17644 31968 17650 32020
rect 19426 31968 19432 32020
rect 19484 32008 19490 32020
rect 23569 32011 23627 32017
rect 23569 32008 23581 32011
rect 19484 31980 23581 32008
rect 19484 31968 19490 31980
rect 23569 31977 23581 31980
rect 23615 31977 23627 32011
rect 23569 31971 23627 31977
rect 23658 31968 23664 32020
rect 23716 32008 23722 32020
rect 23716 31980 24440 32008
rect 23716 31968 23722 31980
rect 23750 31940 23756 31952
rect 15028 31912 15516 31940
rect 15580 31912 19564 31940
rect 11698 31872 11704 31884
rect 10704 31844 11704 31872
rect 10704 31813 10732 31844
rect 11698 31832 11704 31844
rect 11756 31832 11762 31884
rect 12066 31872 12072 31884
rect 12027 31844 12072 31872
rect 12066 31832 12072 31844
rect 12124 31832 12130 31884
rect 12713 31875 12771 31881
rect 12713 31841 12725 31875
rect 12759 31872 12771 31875
rect 12802 31872 12808 31884
rect 12759 31844 12808 31872
rect 12759 31841 12771 31844
rect 12713 31835 12771 31841
rect 12802 31832 12808 31844
rect 12860 31832 12866 31884
rect 9309 31807 9367 31813
rect 9309 31804 9321 31807
rect 9180 31776 9321 31804
rect 9180 31764 9186 31776
rect 9309 31773 9321 31776
rect 9355 31773 9367 31807
rect 9309 31767 9367 31773
rect 9953 31807 10011 31813
rect 9953 31773 9965 31807
rect 9999 31773 10011 31807
rect 9953 31767 10011 31773
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 11054 31764 11060 31816
rect 11112 31804 11118 31816
rect 11333 31807 11391 31813
rect 11333 31804 11345 31807
rect 11112 31776 11345 31804
rect 11112 31764 11118 31776
rect 11333 31773 11345 31776
rect 11379 31773 11391 31807
rect 11333 31767 11391 31773
rect 13170 31764 13176 31816
rect 13228 31804 13234 31816
rect 13541 31807 13599 31813
rect 13541 31804 13553 31807
rect 13228 31776 13553 31804
rect 13228 31764 13234 31776
rect 13541 31773 13553 31776
rect 13587 31773 13599 31807
rect 13541 31767 13599 31773
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31773 14335 31807
rect 14277 31767 14335 31773
rect 11425 31739 11483 31745
rect 11425 31705 11437 31739
rect 11471 31736 11483 31739
rect 12161 31739 12219 31745
rect 12161 31736 12173 31739
rect 11471 31708 12173 31736
rect 11471 31705 11483 31708
rect 11425 31699 11483 31705
rect 12161 31705 12173 31708
rect 12207 31705 12219 31739
rect 12161 31699 12219 31705
rect 13262 31696 13268 31748
rect 13320 31736 13326 31748
rect 14292 31736 14320 31767
rect 14366 31764 14372 31816
rect 14424 31804 14430 31816
rect 15013 31807 15071 31813
rect 14424 31776 14469 31804
rect 14424 31764 14430 31776
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 15059 31776 15148 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 13320 31708 14320 31736
rect 15120 31736 15148 31776
rect 15580 31736 15608 31912
rect 15749 31875 15807 31881
rect 15749 31841 15761 31875
rect 15795 31872 15807 31875
rect 19536 31872 19564 31912
rect 23308 31912 23756 31940
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 15795 31844 16574 31872
rect 19536 31844 21189 31872
rect 15795 31841 15807 31844
rect 15749 31835 15807 31841
rect 16390 31764 16396 31816
rect 16448 31804 16454 31816
rect 16448 31776 16493 31804
rect 16448 31764 16454 31776
rect 16546 31748 16574 31844
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 21177 31835 21235 31841
rect 21821 31875 21879 31881
rect 21821 31841 21833 31875
rect 21867 31872 21879 31875
rect 23308 31872 23336 31912
rect 23750 31900 23756 31912
rect 23808 31900 23814 31952
rect 24118 31900 24124 31952
rect 24176 31940 24182 31952
rect 24302 31940 24308 31952
rect 24176 31912 24308 31940
rect 24176 31900 24182 31912
rect 24302 31900 24308 31912
rect 24360 31900 24366 31952
rect 24412 31940 24440 31980
rect 24578 31968 24584 32020
rect 24636 32008 24642 32020
rect 24636 31980 26464 32008
rect 24636 31968 24642 31980
rect 24412 31912 24716 31940
rect 24578 31872 24584 31884
rect 21867 31844 23336 31872
rect 23400 31844 23612 31872
rect 24539 31844 24584 31872
rect 21867 31841 21879 31844
rect 21821 31835 21879 31841
rect 16850 31764 16856 31816
rect 16908 31804 16914 31816
rect 16945 31807 17003 31813
rect 16945 31804 16957 31807
rect 16908 31776 16957 31804
rect 16908 31764 16914 31776
rect 16945 31773 16957 31776
rect 16991 31773 17003 31807
rect 16945 31767 17003 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 21192 31804 21220 31835
rect 21192 31776 21864 31804
rect 19429 31767 19487 31773
rect 15838 31736 15844 31748
rect 15120 31708 15608 31736
rect 15799 31708 15844 31736
rect 13320 31696 13326 31708
rect 15838 31696 15844 31708
rect 15896 31696 15902 31748
rect 16546 31708 16580 31748
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 19058 31736 19064 31748
rect 16684 31708 19064 31736
rect 8294 31668 8300 31680
rect 8255 31640 8300 31668
rect 8294 31628 8300 31640
rect 8352 31628 8358 31680
rect 10042 31668 10048 31680
rect 10003 31640 10048 31668
rect 10042 31628 10048 31640
rect 10100 31628 10106 31680
rect 10781 31671 10839 31677
rect 10781 31637 10793 31671
rect 10827 31668 10839 31671
rect 10870 31668 10876 31680
rect 10827 31640 10876 31668
rect 10827 31637 10839 31640
rect 10781 31631 10839 31637
rect 10870 31628 10876 31640
rect 10928 31628 10934 31680
rect 10962 31628 10968 31680
rect 11020 31668 11026 31680
rect 13906 31668 13912 31680
rect 11020 31640 13912 31668
rect 11020 31628 11026 31640
rect 13906 31628 13912 31640
rect 13964 31668 13970 31680
rect 15010 31668 15016 31680
rect 13964 31640 15016 31668
rect 13964 31628 13970 31640
rect 15010 31628 15016 31640
rect 15068 31668 15074 31680
rect 16684 31668 16712 31708
rect 19058 31696 19064 31708
rect 19116 31696 19122 31748
rect 15068 31640 16712 31668
rect 15068 31628 15074 31640
rect 18230 31628 18236 31680
rect 18288 31668 18294 31680
rect 19444 31668 19472 31767
rect 19610 31696 19616 31748
rect 19668 31736 19674 31748
rect 19705 31739 19763 31745
rect 19705 31736 19717 31739
rect 19668 31708 19717 31736
rect 19668 31696 19674 31708
rect 19705 31705 19717 31708
rect 19751 31705 19763 31739
rect 19705 31699 19763 31705
rect 20162 31696 20168 31748
rect 20220 31696 20226 31748
rect 20990 31668 20996 31680
rect 18288 31640 20996 31668
rect 18288 31628 18294 31640
rect 20990 31628 20996 31640
rect 21048 31628 21054 31680
rect 21836 31668 21864 31776
rect 22094 31736 22100 31748
rect 22055 31708 22100 31736
rect 22094 31696 22100 31708
rect 22152 31696 22158 31748
rect 22554 31696 22560 31748
rect 22612 31696 22618 31748
rect 23400 31668 23428 31844
rect 23584 31804 23612 31844
rect 24578 31832 24584 31844
rect 24636 31832 24642 31884
rect 24688 31872 24716 31912
rect 24857 31875 24915 31881
rect 24857 31872 24869 31875
rect 24688 31844 24869 31872
rect 24857 31841 24869 31844
rect 24903 31841 24915 31875
rect 24857 31835 24915 31841
rect 24946 31832 24952 31884
rect 25004 31872 25010 31884
rect 26329 31875 26387 31881
rect 26329 31872 26341 31875
rect 25004 31844 26341 31872
rect 25004 31832 25010 31844
rect 26329 31841 26341 31844
rect 26375 31841 26387 31875
rect 26436 31872 26464 31980
rect 27338 31968 27344 32020
rect 27396 32008 27402 32020
rect 36998 32008 37004 32020
rect 27396 31980 37004 32008
rect 27396 31968 27402 31980
rect 36998 31968 37004 31980
rect 37056 31968 37062 32020
rect 27617 31875 27675 31881
rect 27617 31872 27629 31875
rect 26436 31844 27629 31872
rect 26329 31835 26387 31841
rect 27617 31841 27629 31844
rect 27663 31841 27675 31875
rect 27617 31835 27675 31841
rect 36449 31875 36507 31881
rect 36449 31841 36461 31875
rect 36495 31872 36507 31875
rect 36906 31872 36912 31884
rect 36495 31844 36912 31872
rect 36495 31841 36507 31844
rect 36449 31835 36507 31841
rect 36906 31832 36912 31844
rect 36964 31832 36970 31884
rect 23584 31776 24624 31804
rect 24596 31736 24624 31776
rect 36170 31764 36176 31816
rect 36228 31804 36234 31816
rect 38286 31804 38292 31816
rect 36228 31776 36492 31804
rect 38199 31776 38292 31804
rect 36228 31764 36234 31776
rect 24596 31708 24900 31736
rect 21836 31640 23428 31668
rect 24872 31668 24900 31708
rect 25314 31696 25320 31748
rect 25372 31696 25378 31748
rect 26786 31696 26792 31748
rect 26844 31736 26850 31748
rect 26881 31739 26939 31745
rect 26881 31736 26893 31739
rect 26844 31708 26893 31736
rect 26844 31696 26850 31708
rect 26881 31705 26893 31708
rect 26927 31705 26939 31739
rect 36464 31736 36492 31776
rect 38286 31764 38292 31776
rect 38344 31804 38350 31816
rect 39390 31804 39396 31816
rect 38344 31776 39396 31804
rect 38344 31764 38350 31776
rect 39390 31764 39396 31776
rect 39448 31764 39454 31816
rect 36633 31739 36691 31745
rect 36633 31736 36645 31739
rect 36464 31708 36645 31736
rect 26881 31699 26939 31705
rect 36633 31705 36645 31708
rect 36679 31705 36691 31739
rect 36633 31699 36691 31705
rect 25498 31668 25504 31680
rect 24872 31640 25504 31668
rect 25498 31628 25504 31640
rect 25556 31628 25562 31680
rect 31294 31628 31300 31680
rect 31352 31668 31358 31680
rect 36906 31668 36912 31680
rect 31352 31640 36912 31668
rect 31352 31628 31358 31640
rect 36906 31628 36912 31640
rect 36964 31628 36970 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 9033 31467 9091 31473
rect 9033 31433 9045 31467
rect 9079 31464 9091 31467
rect 9214 31464 9220 31476
rect 9079 31436 9220 31464
rect 9079 31433 9091 31436
rect 9033 31427 9091 31433
rect 9214 31424 9220 31436
rect 9272 31424 9278 31476
rect 10410 31464 10416 31476
rect 10371 31436 10416 31464
rect 10410 31424 10416 31436
rect 10468 31424 10474 31476
rect 14826 31464 14832 31476
rect 11072 31436 14832 31464
rect 9769 31399 9827 31405
rect 9769 31365 9781 31399
rect 9815 31396 9827 31399
rect 11072 31396 11100 31436
rect 14826 31424 14832 31436
rect 14884 31424 14890 31476
rect 15470 31424 15476 31476
rect 15528 31464 15534 31476
rect 15841 31467 15899 31473
rect 15841 31464 15853 31467
rect 15528 31436 15853 31464
rect 15528 31424 15534 31436
rect 15841 31433 15853 31436
rect 15887 31433 15899 31467
rect 19426 31464 19432 31476
rect 15841 31427 15899 31433
rect 18892 31436 19432 31464
rect 9815 31368 11100 31396
rect 11793 31399 11851 31405
rect 9815 31365 9827 31368
rect 9769 31359 9827 31365
rect 11793 31365 11805 31399
rect 11839 31396 11851 31399
rect 14369 31399 14427 31405
rect 14369 31396 14381 31399
rect 11839 31368 14381 31396
rect 11839 31365 11851 31368
rect 11793 31359 11851 31365
rect 14369 31365 14381 31368
rect 14415 31365 14427 31399
rect 15286 31396 15292 31408
rect 15247 31368 15292 31396
rect 14369 31359 14427 31365
rect 15286 31356 15292 31368
rect 15344 31356 15350 31408
rect 18892 31396 18920 31436
rect 19426 31424 19432 31436
rect 19484 31424 19490 31476
rect 25222 31464 25228 31476
rect 20640 31436 25228 31464
rect 15764 31368 18920 31396
rect 3878 31288 3884 31340
rect 3936 31328 3942 31340
rect 8389 31331 8447 31337
rect 8389 31328 8401 31331
rect 3936 31300 8401 31328
rect 3936 31288 3942 31300
rect 8389 31297 8401 31300
rect 8435 31297 8447 31331
rect 8389 31291 8447 31297
rect 9030 31288 9036 31340
rect 9088 31328 9094 31340
rect 9217 31331 9275 31337
rect 9217 31328 9229 31331
rect 9088 31300 9229 31328
rect 9088 31288 9094 31300
rect 9217 31297 9229 31300
rect 9263 31297 9275 31331
rect 9217 31291 9275 31297
rect 8478 31124 8484 31136
rect 8439 31096 8484 31124
rect 8478 31084 8484 31096
rect 8536 31084 8542 31136
rect 9232 31124 9260 31291
rect 9306 31288 9312 31340
rect 9364 31328 9370 31340
rect 9677 31331 9735 31337
rect 9677 31328 9689 31331
rect 9364 31300 9689 31328
rect 9364 31288 9370 31300
rect 9677 31297 9689 31300
rect 9723 31297 9735 31331
rect 9677 31291 9735 31297
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10962 31328 10968 31340
rect 10923 31300 10968 31328
rect 10321 31291 10379 31297
rect 10336 31260 10364 31291
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11698 31328 11704 31340
rect 11659 31300 11704 31328
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 12897 31331 12955 31337
rect 12897 31297 12909 31331
rect 12943 31328 12955 31331
rect 13170 31328 13176 31340
rect 12943 31300 13176 31328
rect 12943 31297 12955 31300
rect 12897 31291 12955 31297
rect 13170 31288 13176 31300
rect 13228 31288 13234 31340
rect 13541 31331 13599 31337
rect 13541 31297 13553 31331
rect 13587 31328 13599 31331
rect 13906 31328 13912 31340
rect 13587 31300 13912 31328
rect 13587 31297 13599 31300
rect 13541 31291 13599 31297
rect 13906 31288 13912 31300
rect 13964 31288 13970 31340
rect 15764 31337 15792 31368
rect 18966 31356 18972 31408
rect 19024 31356 19030 31408
rect 20530 31396 20536 31408
rect 20491 31368 20536 31396
rect 20530 31356 20536 31368
rect 20588 31356 20594 31408
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 18230 31328 18236 31340
rect 18191 31300 18236 31328
rect 15749 31291 15807 31297
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 13998 31260 14004 31272
rect 10336 31232 14004 31260
rect 13998 31220 14004 31232
rect 14056 31220 14062 31272
rect 14277 31263 14335 31269
rect 14277 31229 14289 31263
rect 14323 31260 14335 31263
rect 15194 31260 15200 31272
rect 14323 31232 15200 31260
rect 14323 31229 14335 31232
rect 14277 31223 14335 31229
rect 15194 31220 15200 31232
rect 15252 31220 15258 31272
rect 18506 31260 18512 31272
rect 18467 31232 18512 31260
rect 18506 31220 18512 31232
rect 18564 31260 18570 31272
rect 20640 31260 20668 31436
rect 25222 31424 25228 31436
rect 25280 31424 25286 31476
rect 36814 31464 36820 31476
rect 36775 31436 36820 31464
rect 36814 31424 36820 31436
rect 36872 31424 36878 31476
rect 27430 31396 27436 31408
rect 27264 31368 27436 31396
rect 21082 31288 21088 31340
rect 21140 31328 21146 31340
rect 22462 31328 22468 31340
rect 21140 31300 22468 31328
rect 21140 31288 21146 31300
rect 22462 31288 22468 31300
rect 22520 31288 22526 31340
rect 24578 31288 24584 31340
rect 24636 31288 24642 31340
rect 27264 31337 27292 31368
rect 27430 31356 27436 31368
rect 27488 31356 27494 31408
rect 30558 31356 30564 31408
rect 30616 31356 30622 31408
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 28626 31288 28632 31340
rect 28684 31288 28690 31340
rect 33778 31288 33784 31340
rect 33836 31288 33842 31340
rect 36722 31328 36728 31340
rect 36683 31300 36728 31328
rect 36722 31288 36728 31300
rect 36780 31288 36786 31340
rect 18564 31232 20668 31260
rect 18564 31220 18570 31232
rect 20990 31220 20996 31272
rect 21048 31260 21054 31272
rect 21361 31263 21419 31269
rect 21361 31260 21373 31263
rect 21048 31232 21373 31260
rect 21048 31220 21054 31232
rect 21361 31229 21373 31232
rect 21407 31260 21419 31263
rect 23201 31263 23259 31269
rect 23201 31260 23213 31263
rect 21407 31232 23213 31260
rect 21407 31229 21419 31232
rect 21361 31223 21419 31229
rect 23201 31229 23213 31232
rect 23247 31229 23259 31263
rect 23474 31260 23480 31272
rect 23435 31232 23480 31260
rect 23201 31223 23259 31229
rect 23474 31220 23480 31232
rect 23532 31220 23538 31272
rect 25406 31260 25412 31272
rect 25367 31232 25412 31260
rect 25406 31220 25412 31232
rect 25464 31220 25470 31272
rect 25498 31220 25504 31272
rect 25556 31260 25562 31272
rect 27525 31263 27583 31269
rect 27525 31260 27537 31263
rect 25556 31232 27537 31260
rect 25556 31220 25562 31232
rect 27525 31229 27537 31232
rect 27571 31229 27583 31263
rect 29822 31260 29828 31272
rect 29783 31232 29828 31260
rect 27525 31223 27583 31229
rect 29822 31220 29828 31232
rect 29880 31220 29886 31272
rect 30101 31263 30159 31269
rect 30101 31229 30113 31263
rect 30147 31260 30159 31263
rect 32122 31260 32128 31272
rect 30147 31232 32128 31260
rect 30147 31229 30159 31232
rect 30101 31223 30159 31229
rect 32122 31220 32128 31232
rect 32180 31220 32186 31272
rect 32398 31260 32404 31272
rect 32359 31232 32404 31260
rect 32398 31220 32404 31232
rect 32456 31220 32462 31272
rect 32677 31263 32735 31269
rect 32677 31229 32689 31263
rect 32723 31260 32735 31263
rect 32766 31260 32772 31272
rect 32723 31232 32772 31260
rect 32723 31229 32735 31232
rect 32677 31223 32735 31229
rect 32766 31220 32772 31232
rect 32824 31260 32830 31272
rect 34330 31260 34336 31272
rect 32824 31232 34336 31260
rect 32824 31220 32830 31232
rect 34330 31220 34336 31232
rect 34388 31220 34394 31272
rect 37458 31220 37464 31272
rect 37516 31260 37522 31272
rect 37553 31263 37611 31269
rect 37553 31260 37565 31263
rect 37516 31232 37565 31260
rect 37516 31220 37522 31232
rect 37553 31229 37565 31232
rect 37599 31229 37611 31263
rect 37553 31223 37611 31229
rect 11054 31192 11060 31204
rect 11015 31164 11060 31192
rect 11054 31152 11060 31164
rect 11112 31152 11118 31204
rect 12989 31195 13047 31201
rect 12989 31161 13001 31195
rect 13035 31192 13047 31195
rect 17310 31192 17316 31204
rect 13035 31164 17316 31192
rect 13035 31161 13047 31164
rect 12989 31155 13047 31161
rect 17310 31152 17316 31164
rect 17368 31152 17374 31204
rect 17494 31152 17500 31204
rect 17552 31192 17558 31204
rect 21634 31192 21640 31204
rect 17552 31164 18368 31192
rect 17552 31152 17558 31164
rect 13538 31124 13544 31136
rect 9232 31096 13544 31124
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 13633 31127 13691 31133
rect 13633 31093 13645 31127
rect 13679 31124 13691 31127
rect 17862 31124 17868 31136
rect 13679 31096 17868 31124
rect 13679 31093 13691 31096
rect 13633 31087 13691 31093
rect 17862 31084 17868 31096
rect 17920 31084 17926 31136
rect 18340 31124 18368 31164
rect 19904 31164 21640 31192
rect 19904 31124 19932 31164
rect 21634 31152 21640 31164
rect 21692 31152 21698 31204
rect 24872 31164 27384 31192
rect 18340 31096 19932 31124
rect 19978 31084 19984 31136
rect 20036 31124 20042 31136
rect 20036 31096 20081 31124
rect 20036 31084 20042 31096
rect 22646 31084 22652 31136
rect 22704 31124 22710 31136
rect 24872 31124 24900 31164
rect 22704 31096 24900 31124
rect 24949 31127 25007 31133
rect 22704 31084 22710 31096
rect 24949 31093 24961 31127
rect 24995 31124 25007 31127
rect 25222 31124 25228 31136
rect 24995 31096 25228 31124
rect 24995 31093 25007 31096
rect 24949 31087 25007 31093
rect 25222 31084 25228 31096
rect 25280 31084 25286 31136
rect 27356 31124 27384 31164
rect 28997 31127 29055 31133
rect 28997 31124 29009 31127
rect 27356 31096 29009 31124
rect 28997 31093 29009 31096
rect 29043 31124 29055 31127
rect 30466 31124 30472 31136
rect 29043 31096 30472 31124
rect 29043 31093 29055 31096
rect 28997 31087 29055 31093
rect 30466 31084 30472 31096
rect 30524 31084 30530 31136
rect 31202 31084 31208 31136
rect 31260 31124 31266 31136
rect 31570 31124 31576 31136
rect 31260 31096 31576 31124
rect 31260 31084 31266 31096
rect 31570 31084 31576 31096
rect 31628 31084 31634 31136
rect 34149 31127 34207 31133
rect 34149 31093 34161 31127
rect 34195 31124 34207 31127
rect 34238 31124 34244 31136
rect 34195 31096 34244 31124
rect 34195 31093 34207 31096
rect 34149 31087 34207 31093
rect 34238 31084 34244 31096
rect 34296 31084 34302 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 10410 30880 10416 30932
rect 10468 30920 10474 30932
rect 16850 30920 16856 30932
rect 10468 30892 11284 30920
rect 16763 30892 16856 30920
rect 10468 30880 10474 30892
rect 11146 30852 11152 30864
rect 7944 30824 11152 30852
rect 7944 30793 7972 30824
rect 11146 30812 11152 30824
rect 11204 30812 11210 30864
rect 11256 30852 11284 30892
rect 16850 30880 16856 30892
rect 16908 30920 16914 30932
rect 17392 30923 17450 30929
rect 17392 30920 17404 30923
rect 16908 30892 17404 30920
rect 16908 30880 16914 30892
rect 17392 30889 17404 30892
rect 17438 30920 17450 30923
rect 18874 30920 18880 30932
rect 17438 30892 18460 30920
rect 18835 30892 18880 30920
rect 17438 30889 17450 30892
rect 17392 30883 17450 30889
rect 15562 30852 15568 30864
rect 11256 30824 15568 30852
rect 15562 30812 15568 30824
rect 15620 30812 15626 30864
rect 18432 30852 18460 30892
rect 18874 30880 18880 30892
rect 18932 30880 18938 30932
rect 19150 30880 19156 30932
rect 19208 30920 19214 30932
rect 34606 30920 34612 30932
rect 19208 30892 34612 30920
rect 19208 30880 19214 30892
rect 26326 30852 26332 30864
rect 18432 30824 21128 30852
rect 7929 30787 7987 30793
rect 7929 30753 7941 30787
rect 7975 30753 7987 30787
rect 7929 30747 7987 30753
rect 8113 30787 8171 30793
rect 8113 30753 8125 30787
rect 8159 30784 8171 30787
rect 8294 30784 8300 30796
rect 8159 30756 8300 30784
rect 8159 30753 8171 30756
rect 8113 30747 8171 30753
rect 8294 30744 8300 30756
rect 8352 30744 8358 30796
rect 8478 30744 8484 30796
rect 8536 30784 8542 30796
rect 9217 30787 9275 30793
rect 9217 30784 9229 30787
rect 8536 30756 9229 30784
rect 8536 30744 8542 30756
rect 9217 30753 9229 30756
rect 9263 30753 9275 30787
rect 9217 30747 9275 30753
rect 10134 30744 10140 30796
rect 10192 30784 10198 30796
rect 10781 30787 10839 30793
rect 10781 30784 10793 30787
rect 10192 30756 10793 30784
rect 10192 30744 10198 30756
rect 10781 30753 10793 30756
rect 10827 30753 10839 30787
rect 11238 30784 11244 30796
rect 11199 30756 11244 30784
rect 10781 30747 10839 30753
rect 11238 30744 11244 30756
rect 11296 30744 11302 30796
rect 11422 30744 11428 30796
rect 11480 30784 11486 30796
rect 12621 30787 12679 30793
rect 12621 30784 12633 30787
rect 11480 30756 12633 30784
rect 11480 30744 11486 30756
rect 12621 30753 12633 30756
rect 12667 30784 12679 30787
rect 15746 30784 15752 30796
rect 12667 30756 15752 30784
rect 12667 30753 12679 30756
rect 12621 30747 12679 30753
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 17129 30787 17187 30793
rect 17129 30753 17141 30787
rect 17175 30784 17187 30787
rect 18138 30784 18144 30796
rect 17175 30756 18144 30784
rect 17175 30753 17187 30756
rect 17129 30747 17187 30753
rect 18138 30744 18144 30756
rect 18196 30744 18202 30796
rect 18414 30744 18420 30796
rect 18472 30784 18478 30796
rect 18690 30784 18696 30796
rect 18472 30756 18696 30784
rect 18472 30744 18478 30756
rect 18690 30744 18696 30756
rect 18748 30784 18754 30796
rect 19978 30784 19984 30796
rect 18748 30756 19984 30784
rect 18748 30744 18754 30756
rect 19978 30744 19984 30756
rect 20036 30744 20042 30796
rect 20990 30784 20996 30796
rect 20951 30756 20996 30784
rect 20990 30744 20996 30756
rect 21048 30744 21054 30796
rect 21100 30784 21128 30824
rect 24504 30824 26332 30852
rect 24504 30784 24532 30824
rect 26326 30812 26332 30824
rect 26384 30812 26390 30864
rect 21100 30756 24532 30784
rect 24581 30787 24639 30793
rect 24581 30753 24593 30787
rect 24627 30784 24639 30787
rect 25406 30784 25412 30796
rect 24627 30756 25412 30784
rect 24627 30753 24639 30756
rect 24581 30747 24639 30753
rect 25406 30744 25412 30756
rect 25464 30744 25470 30796
rect 26421 30787 26479 30793
rect 26421 30753 26433 30787
rect 26467 30784 26479 30787
rect 26804 30784 26832 30892
rect 34606 30880 34612 30892
rect 34664 30880 34670 30932
rect 37826 30920 37832 30932
rect 37787 30892 37832 30920
rect 37826 30880 37832 30892
rect 37884 30880 37890 30932
rect 38378 30852 38384 30864
rect 36188 30824 38384 30852
rect 26467 30756 26832 30784
rect 26467 30753 26479 30756
rect 26421 30747 26479 30753
rect 27246 30744 27252 30796
rect 27304 30784 27310 30796
rect 29181 30787 29239 30793
rect 29181 30784 29193 30787
rect 27304 30756 29193 30784
rect 27304 30744 27310 30756
rect 29181 30753 29193 30756
rect 29227 30753 29239 30787
rect 29181 30747 29239 30753
rect 30466 30744 30472 30796
rect 30524 30784 30530 30796
rect 31021 30787 31079 30793
rect 31021 30784 31033 30787
rect 30524 30756 31033 30784
rect 30524 30744 30530 30756
rect 31021 30753 31033 30756
rect 31067 30753 31079 30787
rect 31021 30747 31079 30753
rect 34238 30744 34244 30796
rect 34296 30784 34302 30796
rect 35161 30787 35219 30793
rect 35161 30784 35173 30787
rect 34296 30756 35173 30784
rect 34296 30744 34302 30756
rect 35161 30753 35173 30756
rect 35207 30784 35219 30787
rect 36188 30784 36216 30824
rect 38378 30812 38384 30824
rect 38436 30812 38442 30864
rect 37458 30784 37464 30796
rect 35207 30756 36216 30784
rect 37419 30756 37464 30784
rect 35207 30753 35219 30756
rect 35161 30747 35219 30753
rect 37458 30744 37464 30756
rect 37516 30744 37522 30796
rect 1581 30719 1639 30725
rect 1581 30685 1593 30719
rect 1627 30716 1639 30719
rect 1627 30688 2774 30716
rect 1627 30685 1639 30688
rect 1581 30679 1639 30685
rect 2746 30648 2774 30688
rect 3142 30676 3148 30728
rect 3200 30716 3206 30728
rect 11885 30719 11943 30725
rect 3200 30688 8708 30716
rect 3200 30676 3206 30688
rect 8386 30648 8392 30660
rect 2746 30620 8392 30648
rect 8386 30608 8392 30620
rect 8444 30608 8450 30660
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 8202 30540 8208 30592
rect 8260 30580 8266 30592
rect 8573 30583 8631 30589
rect 8573 30580 8585 30583
rect 8260 30552 8585 30580
rect 8260 30540 8266 30552
rect 8573 30549 8585 30552
rect 8619 30549 8631 30583
rect 8680 30580 8708 30688
rect 11885 30685 11897 30719
rect 11931 30685 11943 30719
rect 27430 30716 27436 30728
rect 27391 30688 27436 30716
rect 11885 30679 11943 30685
rect 9309 30651 9367 30657
rect 9309 30617 9321 30651
rect 9355 30648 9367 30651
rect 10042 30648 10048 30660
rect 9355 30620 10048 30648
rect 9355 30617 9367 30620
rect 9309 30611 9367 30617
rect 10042 30608 10048 30620
rect 10100 30608 10106 30660
rect 10229 30651 10287 30657
rect 10229 30617 10241 30651
rect 10275 30648 10287 30651
rect 10410 30648 10416 30660
rect 10275 30620 10416 30648
rect 10275 30617 10287 30620
rect 10229 30611 10287 30617
rect 10410 30608 10416 30620
rect 10468 30608 10474 30660
rect 10870 30608 10876 30660
rect 10928 30648 10934 30660
rect 11900 30648 11928 30679
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 29914 30676 29920 30728
rect 29972 30716 29978 30728
rect 30745 30719 30803 30725
rect 30745 30716 30757 30719
rect 29972 30688 30757 30716
rect 29972 30676 29978 30688
rect 30745 30685 30757 30688
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 32398 30676 32404 30728
rect 32456 30716 32462 30728
rect 34149 30719 34207 30725
rect 34149 30716 34161 30719
rect 32456 30688 34161 30716
rect 32456 30676 32462 30688
rect 34149 30685 34161 30688
rect 34195 30716 34207 30719
rect 34698 30716 34704 30728
rect 34195 30688 34704 30716
rect 34195 30685 34207 30688
rect 34149 30679 34207 30685
rect 34698 30676 34704 30688
rect 34756 30716 34762 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34756 30688 34897 30716
rect 34756 30676 34762 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 37550 30676 37556 30728
rect 37608 30716 37614 30728
rect 37645 30719 37703 30725
rect 37645 30716 37657 30719
rect 37608 30688 37657 30716
rect 37608 30676 37614 30688
rect 37645 30685 37657 30688
rect 37691 30685 37703 30719
rect 37645 30679 37703 30685
rect 10928 30620 10973 30648
rect 11072 30620 11928 30648
rect 10928 30608 10934 30620
rect 11072 30580 11100 30620
rect 12710 30608 12716 30660
rect 12768 30648 12774 30660
rect 13262 30648 13268 30660
rect 12768 30620 12813 30648
rect 13223 30620 13268 30648
rect 12768 30608 12774 30620
rect 13262 30608 13268 30620
rect 13320 30608 13326 30660
rect 13354 30608 13360 30660
rect 13412 30648 13418 30660
rect 13906 30648 13912 30660
rect 13412 30620 13912 30648
rect 13412 30608 13418 30620
rect 13906 30608 13912 30620
rect 13964 30648 13970 30660
rect 15194 30648 15200 30660
rect 13964 30620 15200 30648
rect 13964 30608 13970 30620
rect 15194 30608 15200 30620
rect 15252 30608 15258 30660
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 15473 30651 15531 30657
rect 15473 30648 15485 30651
rect 15344 30620 15485 30648
rect 15344 30608 15350 30620
rect 15473 30617 15485 30620
rect 15519 30617 15531 30651
rect 15473 30611 15531 30617
rect 15565 30651 15623 30657
rect 15565 30617 15577 30651
rect 15611 30617 15623 30651
rect 15565 30611 15623 30617
rect 16485 30651 16543 30657
rect 16485 30617 16497 30651
rect 16531 30648 16543 30651
rect 17494 30648 17500 30660
rect 16531 30620 17500 30648
rect 16531 30617 16543 30620
rect 16485 30611 16543 30617
rect 8680 30552 11100 30580
rect 8573 30543 8631 30549
rect 11882 30540 11888 30592
rect 11940 30580 11946 30592
rect 11977 30583 12035 30589
rect 11977 30580 11989 30583
rect 11940 30552 11989 30580
rect 11940 30540 11946 30552
rect 11977 30549 11989 30552
rect 12023 30549 12035 30583
rect 11977 30543 12035 30549
rect 13078 30540 13084 30592
rect 13136 30580 13142 30592
rect 14277 30583 14335 30589
rect 14277 30580 14289 30583
rect 13136 30552 14289 30580
rect 13136 30540 13142 30552
rect 14277 30549 14289 30552
rect 14323 30549 14335 30583
rect 15580 30580 15608 30611
rect 17494 30608 17500 30620
rect 17552 30608 17558 30660
rect 17954 30608 17960 30660
rect 18012 30608 18018 30660
rect 21266 30648 21272 30660
rect 21227 30620 21272 30648
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 21376 30620 21758 30648
rect 16666 30580 16672 30592
rect 15580 30552 16672 30580
rect 14277 30543 14335 30549
rect 16666 30540 16672 30552
rect 16724 30540 16730 30592
rect 17310 30540 17316 30592
rect 17368 30580 17374 30592
rect 21376 30580 21404 30620
rect 22922 30608 22928 30660
rect 22980 30648 22986 30660
rect 23017 30651 23075 30657
rect 23017 30648 23029 30651
rect 22980 30620 23029 30648
rect 22980 30608 22986 30620
rect 23017 30617 23029 30620
rect 23063 30617 23075 30651
rect 23017 30611 23075 30617
rect 24302 30608 24308 30660
rect 24360 30648 24366 30660
rect 24765 30651 24823 30657
rect 24765 30648 24777 30651
rect 24360 30620 24777 30648
rect 24360 30608 24366 30620
rect 24765 30617 24777 30620
rect 24811 30617 24823 30651
rect 24765 30611 24823 30617
rect 27709 30651 27767 30657
rect 27709 30617 27721 30651
rect 27755 30617 27767 30651
rect 27709 30611 27767 30617
rect 17368 30552 21404 30580
rect 27724 30580 27752 30611
rect 27798 30608 27804 30660
rect 27856 30648 27862 30660
rect 27856 30620 28198 30648
rect 27856 30608 27862 30620
rect 32030 30608 32036 30660
rect 32088 30608 32094 30660
rect 33410 30648 33416 30660
rect 33371 30620 33416 30648
rect 33410 30608 33416 30620
rect 33468 30608 33474 30660
rect 39206 30648 39212 30660
rect 36386 30620 39212 30648
rect 39206 30608 39212 30620
rect 39264 30608 39270 30660
rect 29822 30580 29828 30592
rect 27724 30552 29828 30580
rect 17368 30540 17374 30552
rect 29822 30540 29828 30552
rect 29880 30540 29886 30592
rect 30190 30540 30196 30592
rect 30248 30580 30254 30592
rect 32493 30583 32551 30589
rect 32493 30580 32505 30583
rect 30248 30552 32505 30580
rect 30248 30540 30254 30552
rect 32493 30549 32505 30552
rect 32539 30549 32551 30583
rect 36630 30580 36636 30592
rect 36591 30552 36636 30580
rect 32493 30543 32551 30549
rect 36630 30540 36636 30552
rect 36688 30540 36694 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 10594 30336 10600 30388
rect 10652 30376 10658 30388
rect 16850 30376 16856 30388
rect 10652 30348 16856 30376
rect 10652 30336 10658 30348
rect 16850 30336 16856 30348
rect 16908 30336 16914 30388
rect 17034 30336 17040 30388
rect 17092 30376 17098 30388
rect 21266 30376 21272 30388
rect 17092 30348 21272 30376
rect 17092 30336 17098 30348
rect 21266 30336 21272 30348
rect 21324 30336 21330 30388
rect 29546 30336 29552 30388
rect 29604 30376 29610 30388
rect 38194 30376 38200 30388
rect 29604 30348 36768 30376
rect 38155 30348 38200 30376
rect 29604 30336 29610 30348
rect 14182 30308 14188 30320
rect 14143 30280 14188 30308
rect 14182 30268 14188 30280
rect 14240 30268 14246 30320
rect 14734 30308 14740 30320
rect 14695 30280 14740 30308
rect 14734 30268 14740 30280
rect 14792 30268 14798 30320
rect 15286 30308 15292 30320
rect 15247 30280 15292 30308
rect 15286 30268 15292 30280
rect 15344 30268 15350 30320
rect 15378 30268 15384 30320
rect 15436 30308 15442 30320
rect 15436 30280 15481 30308
rect 15436 30268 15442 30280
rect 16666 30268 16672 30320
rect 16724 30308 16730 30320
rect 16945 30311 17003 30317
rect 16945 30308 16957 30311
rect 16724 30280 16957 30308
rect 16724 30268 16730 30280
rect 16945 30277 16957 30280
rect 16991 30277 17003 30311
rect 16945 30271 17003 30277
rect 17052 30280 18998 30308
rect 10226 30200 10232 30252
rect 10284 30240 10290 30252
rect 10321 30243 10379 30249
rect 10321 30240 10333 30243
rect 10284 30212 10333 30240
rect 10284 30200 10290 30212
rect 10321 30209 10333 30212
rect 10367 30209 10379 30243
rect 10321 30203 10379 30209
rect 10965 30243 11023 30249
rect 10965 30209 10977 30243
rect 11011 30209 11023 30243
rect 10965 30203 11023 30209
rect 9677 30175 9735 30181
rect 9677 30141 9689 30175
rect 9723 30172 9735 30175
rect 9950 30172 9956 30184
rect 9723 30144 9956 30172
rect 9723 30141 9735 30144
rect 9677 30135 9735 30141
rect 9950 30132 9956 30144
rect 10008 30132 10014 30184
rect 10980 30172 11008 30203
rect 11330 30200 11336 30252
rect 11388 30240 11394 30252
rect 11793 30243 11851 30249
rect 11793 30240 11805 30243
rect 11388 30212 11805 30240
rect 11388 30200 11394 30212
rect 11793 30209 11805 30212
rect 11839 30240 11851 30243
rect 11974 30240 11980 30252
rect 11839 30212 11980 30240
rect 11839 30209 11851 30212
rect 11793 30203 11851 30209
rect 11974 30200 11980 30212
rect 12032 30200 12038 30252
rect 12437 30243 12495 30249
rect 12437 30209 12449 30243
rect 12483 30240 12495 30243
rect 12802 30240 12808 30252
rect 12483 30212 12808 30240
rect 12483 30209 12495 30212
rect 12437 30203 12495 30209
rect 12802 30200 12808 30212
rect 12860 30200 12866 30252
rect 13170 30240 13176 30252
rect 13131 30212 13176 30240
rect 13170 30200 13176 30212
rect 13228 30200 13234 30252
rect 16850 30240 16856 30252
rect 16811 30212 16856 30240
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 13262 30172 13268 30184
rect 10980 30144 13268 30172
rect 13262 30132 13268 30144
rect 13320 30132 13326 30184
rect 14093 30175 14151 30181
rect 14093 30141 14105 30175
rect 14139 30172 14151 30175
rect 14458 30172 14464 30184
rect 14139 30144 14464 30172
rect 14139 30141 14151 30144
rect 14093 30135 14151 30141
rect 14458 30132 14464 30144
rect 14516 30132 14522 30184
rect 14918 30132 14924 30184
rect 14976 30172 14982 30184
rect 15562 30172 15568 30184
rect 14976 30144 15240 30172
rect 15523 30144 15568 30172
rect 14976 30132 14982 30144
rect 10413 30107 10471 30113
rect 10413 30073 10425 30107
rect 10459 30104 10471 30107
rect 11238 30104 11244 30116
rect 10459 30076 11244 30104
rect 10459 30073 10471 30076
rect 10413 30067 10471 30073
rect 11238 30064 11244 30076
rect 11296 30064 11302 30116
rect 11885 30107 11943 30113
rect 11885 30073 11897 30107
rect 11931 30104 11943 30107
rect 13170 30104 13176 30116
rect 11931 30076 13176 30104
rect 11931 30073 11943 30076
rect 11885 30067 11943 30073
rect 13170 30064 13176 30076
rect 13228 30064 13234 30116
rect 15010 30104 15016 30116
rect 13280 30076 15016 30104
rect 9490 29996 9496 30048
rect 9548 30036 9554 30048
rect 11057 30039 11115 30045
rect 11057 30036 11069 30039
rect 9548 30008 11069 30036
rect 9548 29996 9554 30008
rect 11057 30005 11069 30008
rect 11103 30005 11115 30039
rect 11057 29999 11115 30005
rect 11974 29996 11980 30048
rect 12032 30036 12038 30048
rect 13280 30045 13308 30076
rect 15010 30064 15016 30076
rect 15068 30064 15074 30116
rect 15212 30104 15240 30144
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 17052 30104 17080 30280
rect 19794 30268 19800 30320
rect 19852 30308 19858 30320
rect 21174 30308 21180 30320
rect 19852 30280 21180 30308
rect 19852 30268 19858 30280
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 23382 30268 23388 30320
rect 23440 30308 23446 30320
rect 27522 30308 27528 30320
rect 23440 30280 24978 30308
rect 27172 30280 27528 30308
rect 23440 30268 23446 30280
rect 18230 30240 18236 30252
rect 18191 30212 18236 30240
rect 18230 30200 18236 30212
rect 18288 30200 18294 30252
rect 23474 30240 23480 30252
rect 20088 30212 23480 30240
rect 18509 30175 18567 30181
rect 18509 30172 18521 30175
rect 18248 30144 18521 30172
rect 18248 30116 18276 30144
rect 18509 30141 18521 30144
rect 18555 30141 18567 30175
rect 18509 30135 18567 30141
rect 18598 30132 18604 30184
rect 18656 30172 18662 30184
rect 19981 30175 20039 30181
rect 19981 30172 19993 30175
rect 18656 30144 19993 30172
rect 18656 30132 18662 30144
rect 19981 30141 19993 30144
rect 20027 30141 20039 30175
rect 19981 30135 20039 30141
rect 15212 30076 17080 30104
rect 18230 30064 18236 30116
rect 18288 30064 18294 30116
rect 12529 30039 12587 30045
rect 12529 30036 12541 30039
rect 12032 30008 12541 30036
rect 12032 29996 12038 30008
rect 12529 30005 12541 30008
rect 12575 30005 12587 30039
rect 12529 29999 12587 30005
rect 13265 30039 13323 30045
rect 13265 30005 13277 30039
rect 13311 30005 13323 30039
rect 13265 29999 13323 30005
rect 13538 29996 13544 30048
rect 13596 30036 13602 30048
rect 20088 30036 20116 30212
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 24210 30240 24216 30252
rect 24171 30212 24216 30240
rect 24210 30200 24216 30212
rect 24268 30200 24274 30252
rect 27172 30249 27200 30280
rect 27522 30268 27528 30280
rect 27580 30268 27586 30320
rect 29270 30268 29276 30320
rect 29328 30308 29334 30320
rect 30190 30308 30196 30320
rect 29328 30280 30196 30308
rect 29328 30268 29334 30280
rect 30190 30268 30196 30280
rect 30248 30268 30254 30320
rect 31478 30268 31484 30320
rect 31536 30308 31542 30320
rect 33413 30311 33471 30317
rect 33413 30308 33425 30311
rect 31536 30280 33425 30308
rect 31536 30268 31542 30280
rect 33413 30277 33425 30280
rect 33459 30277 33471 30311
rect 35066 30308 35072 30320
rect 33413 30271 33471 30277
rect 34532 30280 35072 30308
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 28534 30200 28540 30252
rect 28592 30200 28598 30252
rect 31294 30200 31300 30252
rect 31352 30200 31358 30252
rect 33321 30243 33379 30249
rect 33321 30209 33333 30243
rect 33367 30240 33379 30243
rect 34532 30240 34560 30280
rect 35066 30268 35072 30280
rect 35124 30268 35130 30320
rect 36740 30317 36768 30348
rect 38194 30336 38200 30348
rect 38252 30336 38258 30388
rect 36725 30311 36783 30317
rect 36725 30277 36737 30311
rect 36771 30277 36783 30311
rect 36725 30271 36783 30277
rect 34698 30240 34704 30252
rect 33367 30212 34560 30240
rect 34659 30212 34704 30240
rect 33367 30209 33379 30212
rect 33321 30203 33379 30209
rect 34698 30200 34704 30212
rect 34756 30200 34762 30252
rect 36078 30200 36084 30252
rect 36136 30200 36142 30252
rect 36998 30200 37004 30252
rect 37056 30240 37062 30252
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 37056 30212 38025 30240
rect 37056 30200 37062 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 20162 30132 20168 30184
rect 20220 30172 20226 30184
rect 26237 30175 26295 30181
rect 26237 30172 26249 30175
rect 20220 30144 26249 30172
rect 20220 30132 20226 30144
rect 26237 30141 26249 30144
rect 26283 30141 26295 30175
rect 27433 30175 27491 30181
rect 27433 30172 27445 30175
rect 26237 30135 26295 30141
rect 26344 30144 27445 30172
rect 24210 30104 24216 30116
rect 22066 30076 24216 30104
rect 13596 30008 20116 30036
rect 13596 29996 13602 30008
rect 20622 29996 20628 30048
rect 20680 30036 20686 30048
rect 22066 30036 22094 30076
rect 24210 30064 24216 30076
rect 24268 30064 24274 30116
rect 26344 30104 26372 30144
rect 25884 30076 26372 30104
rect 20680 30008 22094 30036
rect 20680 29996 20686 30008
rect 23934 29996 23940 30048
rect 23992 30036 23998 30048
rect 24470 30039 24528 30045
rect 24470 30036 24482 30039
rect 23992 30008 24482 30036
rect 23992 29996 23998 30008
rect 24470 30005 24482 30008
rect 24516 30036 24528 30039
rect 24670 30036 24676 30048
rect 24516 30008 24676 30036
rect 24516 30005 24528 30008
rect 24470 29999 24528 30005
rect 24670 29996 24676 30008
rect 24728 29996 24734 30048
rect 24854 29996 24860 30048
rect 24912 30036 24918 30048
rect 25884 30036 25912 30076
rect 24912 30008 25912 30036
rect 27264 30036 27292 30144
rect 27433 30141 27445 30144
rect 27479 30141 27491 30175
rect 27433 30135 27491 30141
rect 27522 30132 27528 30184
rect 27580 30172 27586 30184
rect 29914 30172 29920 30184
rect 27580 30144 29920 30172
rect 27580 30132 27586 30144
rect 29914 30132 29920 30144
rect 29972 30132 29978 30184
rect 34606 30132 34612 30184
rect 34664 30172 34670 30184
rect 34977 30175 35035 30181
rect 34977 30172 34989 30175
rect 34664 30144 34989 30172
rect 34664 30132 34670 30144
rect 34977 30141 34989 30144
rect 35023 30141 35035 30175
rect 34977 30135 35035 30141
rect 35066 30132 35072 30184
rect 35124 30172 35130 30184
rect 36354 30172 36360 30184
rect 35124 30144 36360 30172
rect 35124 30132 35130 30144
rect 36354 30132 36360 30144
rect 36412 30132 36418 30184
rect 28074 30036 28080 30048
rect 27264 30008 28080 30036
rect 24912 29996 24918 30008
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28902 30036 28908 30048
rect 28863 30008 28908 30036
rect 28902 29996 28908 30008
rect 28960 29996 28966 30048
rect 31386 29996 31392 30048
rect 31444 30036 31450 30048
rect 31662 30036 31668 30048
rect 31444 30008 31668 30036
rect 31444 29996 31450 30008
rect 31662 29996 31668 30008
rect 31720 29996 31726 30048
rect 32122 29996 32128 30048
rect 32180 30036 32186 30048
rect 33042 30036 33048 30048
rect 32180 30008 33048 30036
rect 32180 29996 32186 30008
rect 33042 29996 33048 30008
rect 33100 29996 33106 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 8202 29832 8208 29844
rect 8163 29804 8208 29832
rect 8202 29792 8208 29804
rect 8260 29792 8266 29844
rect 10597 29835 10655 29841
rect 10597 29801 10609 29835
rect 10643 29832 10655 29835
rect 11790 29832 11796 29844
rect 10643 29804 11796 29832
rect 10643 29801 10655 29804
rect 10597 29795 10655 29801
rect 11790 29792 11796 29804
rect 11848 29792 11854 29844
rect 13170 29792 13176 29844
rect 13228 29832 13234 29844
rect 14734 29832 14740 29844
rect 13228 29804 14740 29832
rect 13228 29792 13234 29804
rect 14734 29792 14740 29804
rect 14792 29792 14798 29844
rect 14829 29835 14887 29841
rect 14829 29801 14841 29835
rect 14875 29832 14887 29835
rect 15838 29832 15844 29844
rect 14875 29804 15844 29832
rect 14875 29801 14887 29804
rect 14829 29795 14887 29801
rect 15838 29792 15844 29804
rect 15896 29792 15902 29844
rect 16850 29792 16856 29844
rect 16908 29832 16914 29844
rect 19058 29832 19064 29844
rect 16908 29804 19064 29832
rect 16908 29792 16914 29804
rect 19058 29792 19064 29804
rect 19116 29792 19122 29844
rect 19686 29835 19744 29841
rect 19686 29832 19698 29835
rect 19536 29804 19698 29832
rect 1581 29767 1639 29773
rect 1581 29733 1593 29767
rect 1627 29764 1639 29767
rect 9306 29764 9312 29776
rect 1627 29736 9312 29764
rect 1627 29733 1639 29736
rect 1581 29727 1639 29733
rect 9306 29724 9312 29736
rect 9364 29724 9370 29776
rect 13262 29724 13268 29776
rect 13320 29764 13326 29776
rect 13633 29767 13691 29773
rect 13633 29764 13645 29767
rect 13320 29736 13645 29764
rect 13320 29724 13326 29736
rect 13633 29733 13645 29736
rect 13679 29764 13691 29767
rect 16025 29767 16083 29773
rect 16025 29764 16037 29767
rect 13679 29736 16037 29764
rect 13679 29733 13691 29736
rect 13633 29727 13691 29733
rect 16025 29733 16037 29736
rect 16071 29733 16083 29767
rect 16025 29727 16083 29733
rect 18966 29724 18972 29776
rect 19024 29764 19030 29776
rect 19536 29764 19564 29804
rect 19686 29801 19698 29804
rect 19732 29801 19744 29835
rect 19686 29795 19744 29801
rect 19794 29792 19800 29844
rect 19852 29832 19858 29844
rect 26878 29832 26884 29844
rect 19852 29804 26884 29832
rect 19852 29792 19858 29804
rect 26878 29792 26884 29804
rect 26936 29792 26942 29844
rect 35342 29832 35348 29844
rect 26988 29804 35348 29832
rect 19024 29736 19564 29764
rect 19024 29724 19030 29736
rect 20898 29724 20904 29776
rect 20956 29764 20962 29776
rect 23566 29764 23572 29776
rect 20956 29736 23572 29764
rect 20956 29724 20962 29736
rect 23566 29724 23572 29736
rect 23624 29724 23630 29776
rect 9950 29696 9956 29708
rect 9911 29668 9956 29696
rect 9950 29656 9956 29668
rect 10008 29656 10014 29708
rect 11514 29696 11520 29708
rect 11475 29668 11520 29696
rect 11514 29656 11520 29668
rect 11572 29656 11578 29708
rect 13078 29696 13084 29708
rect 13039 29668 13084 29696
rect 13078 29656 13084 29668
rect 13136 29656 13142 29708
rect 21177 29699 21235 29705
rect 21177 29696 21189 29699
rect 14752 29668 21189 29696
rect 1762 29628 1768 29640
rect 1723 29600 1768 29628
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 7282 29588 7288 29640
rect 7340 29628 7346 29640
rect 7558 29628 7564 29640
rect 7340 29600 7564 29628
rect 7340 29588 7346 29600
rect 7558 29588 7564 29600
rect 7616 29588 7622 29640
rect 7742 29628 7748 29640
rect 7703 29600 7748 29628
rect 7742 29588 7748 29600
rect 7800 29588 7806 29640
rect 9490 29628 9496 29640
rect 9451 29600 9496 29628
rect 9490 29588 9496 29600
rect 9548 29588 9554 29640
rect 9674 29588 9680 29640
rect 9732 29628 9738 29640
rect 14752 29637 14780 29668
rect 21177 29665 21189 29668
rect 21223 29696 21235 29699
rect 22094 29696 22100 29708
rect 21223 29668 22100 29696
rect 21223 29665 21235 29668
rect 21177 29659 21235 29665
rect 22094 29656 22100 29668
rect 22152 29656 22158 29708
rect 24581 29699 24639 29705
rect 24581 29665 24593 29699
rect 24627 29696 24639 29699
rect 24854 29696 24860 29708
rect 24627 29668 24860 29696
rect 24627 29665 24639 29668
rect 24581 29659 24639 29665
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 25590 29656 25596 29708
rect 25648 29696 25654 29708
rect 25648 29668 26740 29696
rect 25648 29656 25654 29668
rect 10137 29631 10195 29637
rect 10137 29628 10149 29631
rect 9732 29600 10149 29628
rect 9732 29588 9738 29600
rect 10137 29597 10149 29600
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29597 14795 29631
rect 14737 29591 14795 29597
rect 18138 29588 18144 29640
rect 18196 29628 18202 29640
rect 18984 29628 19334 29638
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18196 29610 19441 29628
rect 18196 29600 19012 29610
rect 19306 29600 19441 29610
rect 18196 29588 18202 29600
rect 11146 29560 11152 29572
rect 11107 29532 11152 29560
rect 11146 29520 11152 29532
rect 11204 29520 11210 29572
rect 11238 29520 11244 29572
rect 11296 29560 11302 29572
rect 11296 29532 11341 29560
rect 11296 29520 11302 29532
rect 13170 29520 13176 29572
rect 13228 29560 13234 29572
rect 15470 29560 15476 29572
rect 13228 29532 13273 29560
rect 15431 29532 15476 29560
rect 13228 29520 13234 29532
rect 15470 29520 15476 29532
rect 15528 29520 15534 29572
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 15620 29532 15665 29560
rect 15620 29520 15626 29532
rect 19306 29504 19334 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 24486 29628 24492 29640
rect 19429 29591 19487 29597
rect 22066 29600 24492 29628
rect 20162 29520 20168 29572
rect 20220 29520 20226 29572
rect 5902 29452 5908 29504
rect 5960 29492 5966 29504
rect 9309 29495 9367 29501
rect 9309 29492 9321 29495
rect 5960 29464 9321 29492
rect 5960 29452 5966 29464
rect 9309 29461 9321 29464
rect 9355 29461 9367 29495
rect 9309 29455 9367 29461
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 12894 29492 12900 29504
rect 9456 29464 12900 29492
rect 9456 29452 9462 29464
rect 12894 29452 12900 29464
rect 12952 29452 12958 29504
rect 19306 29464 19340 29504
rect 19334 29452 19340 29464
rect 19392 29452 19398 29504
rect 21266 29452 21272 29504
rect 21324 29492 21330 29504
rect 22066 29492 22094 29600
rect 24486 29588 24492 29600
rect 24544 29588 24550 29640
rect 22922 29520 22928 29572
rect 22980 29560 22986 29572
rect 24857 29563 24915 29569
rect 24857 29560 24869 29563
rect 22980 29532 24869 29560
rect 22980 29520 22986 29532
rect 24857 29529 24869 29532
rect 24903 29529 24915 29563
rect 26602 29560 26608 29572
rect 26082 29532 26608 29560
rect 24857 29523 24915 29529
rect 26602 29520 26608 29532
rect 26660 29520 26666 29572
rect 26712 29560 26740 29668
rect 26988 29637 27016 29804
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 33042 29724 33048 29776
rect 33100 29764 33106 29776
rect 33100 29736 35020 29764
rect 33100 29724 33106 29736
rect 29914 29656 29920 29708
rect 29972 29696 29978 29708
rect 30469 29699 30527 29705
rect 30469 29696 30481 29699
rect 29972 29668 30481 29696
rect 29972 29656 29978 29668
rect 30469 29665 30481 29668
rect 30515 29665 30527 29699
rect 30469 29659 30527 29665
rect 31389 29699 31447 29705
rect 31389 29665 31401 29699
rect 31435 29696 31447 29699
rect 32398 29696 32404 29708
rect 31435 29668 32404 29696
rect 31435 29665 31447 29668
rect 31389 29659 31447 29665
rect 32398 29656 32404 29668
rect 32456 29656 32462 29708
rect 34698 29656 34704 29708
rect 34756 29696 34762 29708
rect 34885 29699 34943 29705
rect 34885 29696 34897 29699
rect 34756 29668 34897 29696
rect 34756 29656 34762 29668
rect 34885 29665 34897 29668
rect 34931 29665 34943 29699
rect 34992 29696 35020 29736
rect 36633 29699 36691 29705
rect 36633 29696 36645 29699
rect 34992 29668 36645 29696
rect 34885 29659 34943 29665
rect 36633 29665 36645 29668
rect 36679 29665 36691 29699
rect 36633 29659 36691 29665
rect 26973 29631 27031 29637
rect 26973 29597 26985 29631
rect 27019 29597 27031 29631
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 26973 29591 27031 29597
rect 29656 29600 29745 29628
rect 29546 29560 29552 29572
rect 26712 29532 29552 29560
rect 29546 29520 29552 29532
rect 29604 29520 29610 29572
rect 29656 29504 29684 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 36722 29588 36728 29640
rect 36780 29628 36786 29640
rect 37277 29631 37335 29637
rect 37277 29628 37289 29631
rect 36780 29600 37289 29628
rect 36780 29588 36786 29600
rect 37277 29597 37289 29600
rect 37323 29597 37335 29631
rect 37277 29591 37335 29597
rect 37826 29588 37832 29640
rect 37884 29628 37890 29640
rect 38013 29631 38071 29637
rect 38013 29628 38025 29631
rect 37884 29600 38025 29628
rect 37884 29588 37890 29600
rect 38013 29597 38025 29600
rect 38059 29597 38071 29631
rect 38013 29591 38071 29597
rect 31662 29560 31668 29572
rect 31623 29532 31668 29560
rect 31662 29520 31668 29532
rect 31720 29520 31726 29572
rect 32214 29520 32220 29572
rect 32272 29520 32278 29572
rect 35161 29563 35219 29569
rect 35161 29529 35173 29563
rect 35207 29529 35219 29563
rect 37918 29560 37924 29572
rect 36386 29532 37924 29560
rect 35161 29523 35219 29529
rect 21324 29464 22094 29492
rect 21324 29452 21330 29464
rect 23566 29452 23572 29504
rect 23624 29492 23630 29504
rect 25130 29492 25136 29504
rect 23624 29464 25136 29492
rect 23624 29452 23630 29464
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 26329 29495 26387 29501
rect 26329 29461 26341 29495
rect 26375 29492 26387 29495
rect 27430 29492 27436 29504
rect 26375 29464 27436 29492
rect 26375 29461 26387 29464
rect 26329 29455 26387 29461
rect 27430 29452 27436 29464
rect 27488 29452 27494 29504
rect 28074 29452 28080 29504
rect 28132 29492 28138 29504
rect 28261 29495 28319 29501
rect 28261 29492 28273 29495
rect 28132 29464 28273 29492
rect 28132 29452 28138 29464
rect 28261 29461 28273 29464
rect 28307 29492 28319 29495
rect 29638 29492 29644 29504
rect 28307 29464 29644 29492
rect 28307 29461 28319 29464
rect 28261 29455 28319 29461
rect 29638 29452 29644 29464
rect 29696 29452 29702 29504
rect 33134 29492 33140 29504
rect 33095 29464 33140 29492
rect 33134 29452 33140 29464
rect 33192 29452 33198 29504
rect 34146 29452 34152 29504
rect 34204 29492 34210 29504
rect 35176 29492 35204 29523
rect 37918 29520 37924 29532
rect 37976 29520 37982 29572
rect 34204 29464 35204 29492
rect 37093 29495 37151 29501
rect 34204 29452 34210 29464
rect 37093 29461 37105 29495
rect 37139 29492 37151 29495
rect 37642 29492 37648 29504
rect 37139 29464 37648 29492
rect 37139 29461 37151 29464
rect 37093 29455 37151 29461
rect 37642 29452 37648 29464
rect 37700 29452 37706 29504
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9769 29291 9827 29297
rect 9769 29257 9781 29291
rect 9815 29288 9827 29291
rect 9815 29260 12434 29288
rect 9815 29257 9827 29260
rect 9769 29251 9827 29257
rect 6638 29180 6644 29232
rect 6696 29220 6702 29232
rect 11057 29223 11115 29229
rect 6696 29192 10364 29220
rect 6696 29180 6702 29192
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 1854 29152 1860 29164
rect 1627 29124 1860 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 1854 29112 1860 29124
rect 1912 29112 1918 29164
rect 7650 29112 7656 29164
rect 7708 29152 7714 29164
rect 9677 29155 9735 29161
rect 9677 29152 9689 29155
rect 7708 29124 9689 29152
rect 7708 29112 7714 29124
rect 9677 29121 9689 29124
rect 9723 29152 9735 29155
rect 10042 29152 10048 29164
rect 9723 29124 10048 29152
rect 9723 29121 9735 29124
rect 9677 29115 9735 29121
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 10336 29161 10364 29192
rect 11057 29189 11069 29223
rect 11103 29220 11115 29223
rect 11885 29223 11943 29229
rect 11885 29220 11897 29223
rect 11103 29192 11897 29220
rect 11103 29189 11115 29192
rect 11057 29183 11115 29189
rect 11885 29189 11897 29192
rect 11931 29189 11943 29223
rect 12406 29220 12434 29260
rect 13170 29248 13176 29300
rect 13228 29288 13234 29300
rect 13633 29291 13691 29297
rect 13633 29288 13645 29291
rect 13228 29260 13645 29288
rect 13228 29248 13234 29260
rect 13633 29257 13645 29260
rect 13679 29257 13691 29291
rect 21266 29288 21272 29300
rect 13633 29251 13691 29257
rect 16868 29260 21272 29288
rect 12406 29192 13676 29220
rect 11885 29183 11943 29189
rect 10321 29155 10379 29161
rect 10321 29121 10333 29155
rect 10367 29121 10379 29155
rect 10962 29152 10968 29164
rect 10923 29124 10968 29152
rect 10321 29115 10379 29121
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 12894 29152 12900 29164
rect 12807 29124 12900 29152
rect 12894 29112 12900 29124
rect 12952 29152 12958 29164
rect 13538 29152 13544 29164
rect 12952 29124 13400 29152
rect 13499 29124 13544 29152
rect 12952 29112 12958 29124
rect 10413 29087 10471 29093
rect 10413 29053 10425 29087
rect 10459 29084 10471 29087
rect 11422 29084 11428 29096
rect 10459 29056 11428 29084
rect 10459 29053 10471 29056
rect 10413 29047 10471 29053
rect 11422 29044 11428 29056
rect 11480 29044 11486 29096
rect 11793 29087 11851 29093
rect 11793 29053 11805 29087
rect 11839 29053 11851 29087
rect 12158 29084 12164 29096
rect 12119 29056 12164 29084
rect 11793 29047 11851 29053
rect 1762 29016 1768 29028
rect 1723 28988 1768 29016
rect 1762 28976 1768 28988
rect 1820 28976 1826 29028
rect 7558 28976 7564 29028
rect 7616 29016 7622 29028
rect 7616 28988 8340 29016
rect 7616 28976 7622 28988
rect 8312 28948 8340 28988
rect 9766 28976 9772 29028
rect 9824 29016 9830 29028
rect 11808 29016 11836 29047
rect 12158 29044 12164 29056
rect 12216 29044 12222 29096
rect 9824 28988 11836 29016
rect 9824 28976 9830 28988
rect 11238 28948 11244 28960
rect 8312 28920 11244 28948
rect 11238 28908 11244 28920
rect 11296 28948 11302 28960
rect 12066 28948 12072 28960
rect 11296 28920 12072 28948
rect 11296 28908 11302 28920
rect 12066 28908 12072 28920
rect 12124 28908 12130 28960
rect 12986 28948 12992 28960
rect 12947 28920 12992 28948
rect 12986 28908 12992 28920
rect 13044 28908 13050 28960
rect 13372 28948 13400 29124
rect 13538 29112 13544 29124
rect 13596 29112 13602 29164
rect 13648 29016 13676 29192
rect 13722 29180 13728 29232
rect 13780 29220 13786 29232
rect 15654 29229 15660 29232
rect 14461 29223 14519 29229
rect 14461 29220 14473 29223
rect 13780 29192 14473 29220
rect 13780 29180 13786 29192
rect 14461 29189 14473 29192
rect 14507 29189 14519 29223
rect 14461 29183 14519 29189
rect 15650 29183 15660 29229
rect 15712 29220 15718 29232
rect 15712 29192 15750 29220
rect 15654 29180 15660 29183
rect 15712 29180 15718 29192
rect 16868 29161 16896 29260
rect 21266 29248 21272 29260
rect 21324 29248 21330 29300
rect 26786 29288 26792 29300
rect 22112 29260 26792 29288
rect 22112 29232 22140 29260
rect 17954 29180 17960 29232
rect 18012 29220 18018 29232
rect 20530 29220 20536 29232
rect 18012 29192 18998 29220
rect 20491 29192 20536 29220
rect 18012 29180 18018 29192
rect 20530 29180 20536 29192
rect 20588 29220 20594 29232
rect 22094 29220 22100 29232
rect 20588 29192 22100 29220
rect 20588 29180 20594 29192
rect 22094 29180 22100 29192
rect 22152 29180 22158 29232
rect 23290 29220 23296 29232
rect 23251 29192 23296 29220
rect 23290 29180 23296 29192
rect 23348 29180 23354 29232
rect 23842 29180 23848 29232
rect 23900 29180 23906 29232
rect 25332 29229 25360 29260
rect 26786 29248 26792 29260
rect 26844 29288 26850 29300
rect 28074 29288 28080 29300
rect 26844 29260 28080 29288
rect 26844 29248 26850 29260
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 33594 29248 33600 29300
rect 33652 29288 33658 29300
rect 34241 29291 34299 29297
rect 34241 29288 34253 29291
rect 33652 29260 34253 29288
rect 33652 29248 33658 29260
rect 34241 29257 34253 29260
rect 34287 29257 34299 29291
rect 34241 29251 34299 29257
rect 25317 29223 25375 29229
rect 25317 29189 25329 29223
rect 25363 29189 25375 29223
rect 25317 29183 25375 29189
rect 33226 29180 33232 29232
rect 33284 29180 33290 29232
rect 16853 29155 16911 29161
rect 16853 29121 16865 29155
rect 16899 29121 16911 29155
rect 16853 29115 16911 29121
rect 19720 29124 21404 29152
rect 13814 29044 13820 29096
rect 13872 29084 13878 29096
rect 14369 29087 14427 29093
rect 14369 29084 14381 29087
rect 13872 29056 14381 29084
rect 13872 29044 13878 29056
rect 14369 29053 14381 29056
rect 14415 29053 14427 29087
rect 14369 29047 14427 29053
rect 14550 29044 14556 29096
rect 14608 29084 14614 29096
rect 14645 29087 14703 29093
rect 14645 29084 14657 29087
rect 14608 29056 14657 29084
rect 14608 29044 14614 29056
rect 14645 29053 14657 29056
rect 14691 29053 14703 29087
rect 14645 29047 14703 29053
rect 14826 29044 14832 29096
rect 14884 29084 14890 29096
rect 15565 29087 15623 29093
rect 15565 29084 15577 29087
rect 14884 29072 15424 29084
rect 15488 29072 15577 29084
rect 14884 29056 15577 29072
rect 14884 29044 14890 29056
rect 15396 29044 15516 29056
rect 15565 29053 15577 29056
rect 15611 29053 15623 29087
rect 15565 29047 15623 29053
rect 15930 29044 15936 29096
rect 15988 29084 15994 29096
rect 16209 29087 16267 29093
rect 16209 29084 16221 29087
rect 15988 29056 16221 29084
rect 15988 29044 15994 29056
rect 16209 29053 16221 29056
rect 16255 29084 16267 29087
rect 16298 29084 16304 29096
rect 16255 29056 16304 29084
rect 16255 29053 16267 29056
rect 16209 29047 16267 29053
rect 16298 29044 16304 29056
rect 16356 29044 16362 29096
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 18233 29087 18291 29093
rect 18233 29084 18245 29087
rect 18196 29056 18245 29084
rect 18196 29044 18202 29056
rect 18233 29053 18245 29056
rect 18279 29053 18291 29087
rect 18233 29047 18291 29053
rect 15286 29016 15292 29028
rect 13648 28988 15292 29016
rect 15286 28976 15292 28988
rect 15344 28976 15350 29028
rect 19720 29016 19748 29124
rect 20714 29044 20720 29096
rect 20772 29084 20778 29096
rect 21269 29087 21327 29093
rect 21269 29084 21281 29087
rect 20772 29056 21281 29084
rect 20772 29044 20778 29056
rect 21269 29053 21281 29056
rect 21315 29053 21327 29087
rect 21376 29084 21404 29124
rect 21542 29112 21548 29164
rect 21600 29152 21606 29164
rect 22922 29152 22928 29164
rect 21600 29124 22928 29152
rect 21600 29112 21606 29124
rect 22922 29112 22928 29124
rect 22980 29112 22986 29164
rect 24578 29112 24584 29164
rect 24636 29152 24642 29164
rect 31570 29152 31576 29164
rect 24636 29124 31576 29152
rect 24636 29112 24642 29124
rect 31570 29112 31576 29124
rect 31628 29112 31634 29164
rect 32398 29112 32404 29164
rect 32456 29152 32462 29164
rect 32493 29155 32551 29161
rect 32493 29152 32505 29155
rect 32456 29124 32505 29152
rect 32456 29112 32462 29124
rect 32493 29121 32505 29124
rect 32539 29121 32551 29155
rect 32493 29115 32551 29121
rect 38013 29155 38071 29161
rect 38013 29121 38025 29155
rect 38059 29152 38071 29155
rect 39114 29152 39120 29164
rect 38059 29124 39120 29152
rect 38059 29121 38071 29124
rect 38013 29115 38071 29121
rect 39114 29112 39120 29124
rect 39172 29112 39178 29164
rect 22554 29084 22560 29096
rect 21376 29056 22560 29084
rect 21269 29047 21327 29053
rect 22554 29044 22560 29056
rect 22612 29044 22618 29096
rect 23014 29084 23020 29096
rect 22975 29056 23020 29084
rect 23014 29044 23020 29056
rect 23072 29044 23078 29096
rect 24765 29087 24823 29093
rect 24765 29084 24777 29087
rect 23124 29056 24777 29084
rect 19978 29016 19984 29028
rect 16776 28988 17080 29016
rect 16776 28948 16804 28988
rect 16942 28948 16948 28960
rect 13372 28920 16804 28948
rect 16903 28920 16948 28948
rect 16942 28908 16948 28920
rect 17000 28908 17006 28960
rect 17052 28948 17080 28988
rect 19536 28988 19748 29016
rect 19939 28988 19984 29016
rect 17770 28948 17776 28960
rect 17052 28920 17776 28948
rect 17770 28908 17776 28920
rect 17828 28908 17834 28960
rect 18496 28951 18554 28957
rect 18496 28917 18508 28951
rect 18542 28948 18554 28951
rect 18966 28948 18972 28960
rect 18542 28920 18972 28948
rect 18542 28917 18554 28920
rect 18496 28911 18554 28917
rect 18966 28908 18972 28920
rect 19024 28908 19030 28960
rect 19242 28908 19248 28960
rect 19300 28948 19306 28960
rect 19536 28948 19564 28988
rect 19978 28976 19984 28988
rect 20036 29016 20042 29028
rect 20990 29016 20996 29028
rect 20036 28988 20996 29016
rect 20036 28976 20042 28988
rect 20990 28976 20996 28988
rect 21048 28976 21054 29028
rect 21082 28976 21088 29028
rect 21140 29016 21146 29028
rect 23124 29016 23152 29056
rect 24765 29053 24777 29056
rect 24811 29053 24823 29087
rect 24765 29047 24823 29053
rect 24854 29044 24860 29096
rect 24912 29084 24918 29096
rect 26053 29087 26111 29093
rect 26053 29084 26065 29087
rect 24912 29056 26065 29084
rect 24912 29044 24918 29056
rect 26053 29053 26065 29056
rect 26099 29053 26111 29087
rect 26053 29047 26111 29053
rect 26878 29044 26884 29096
rect 26936 29084 26942 29096
rect 32306 29084 32312 29096
rect 26936 29056 32312 29084
rect 26936 29044 26942 29056
rect 32306 29044 32312 29056
rect 32364 29044 32370 29096
rect 21140 28988 23152 29016
rect 21140 28976 21146 28988
rect 24946 28976 24952 29028
rect 25004 29016 25010 29028
rect 25590 29016 25596 29028
rect 25004 28988 25596 29016
rect 25004 28976 25010 28988
rect 25590 28976 25596 28988
rect 25648 28976 25654 29028
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 19300 28920 19564 28948
rect 19300 28908 19306 28920
rect 20070 28908 20076 28960
rect 20128 28948 20134 28960
rect 26878 28948 26884 28960
rect 20128 28920 26884 28948
rect 20128 28908 20134 28920
rect 26878 28908 26884 28920
rect 26936 28908 26942 28960
rect 32582 28908 32588 28960
rect 32640 28948 32646 28960
rect 32750 28951 32808 28957
rect 32750 28948 32762 28951
rect 32640 28920 32762 28948
rect 32640 28908 32646 28920
rect 32750 28917 32762 28920
rect 32796 28948 32808 28951
rect 36630 28948 36636 28960
rect 32796 28920 36636 28948
rect 32796 28917 32808 28920
rect 32750 28911 32808 28917
rect 36630 28908 36636 28920
rect 36688 28908 36694 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1578 28704 1584 28756
rect 1636 28744 1642 28756
rect 6641 28747 6699 28753
rect 6641 28744 6653 28747
rect 1636 28716 6653 28744
rect 1636 28704 1642 28716
rect 6641 28713 6653 28716
rect 6687 28713 6699 28747
rect 10502 28744 10508 28756
rect 10463 28716 10508 28744
rect 6641 28707 6699 28713
rect 10502 28704 10508 28716
rect 10560 28704 10566 28756
rect 11701 28747 11759 28753
rect 11701 28713 11713 28747
rect 11747 28744 11759 28747
rect 11790 28744 11796 28756
rect 11747 28716 11796 28744
rect 11747 28713 11759 28716
rect 11701 28707 11759 28713
rect 11790 28704 11796 28716
rect 11848 28704 11854 28756
rect 13633 28747 13691 28753
rect 13633 28713 13645 28747
rect 13679 28744 13691 28747
rect 13722 28744 13728 28756
rect 13679 28716 13728 28744
rect 13679 28713 13691 28716
rect 13633 28707 13691 28713
rect 13722 28704 13728 28716
rect 13780 28704 13786 28756
rect 14182 28704 14188 28756
rect 14240 28744 14246 28756
rect 14369 28747 14427 28753
rect 14369 28744 14381 28747
rect 14240 28716 14381 28744
rect 14240 28704 14246 28716
rect 14369 28713 14381 28716
rect 14415 28713 14427 28747
rect 14369 28707 14427 28713
rect 15013 28747 15071 28753
rect 15013 28713 15025 28747
rect 15059 28744 15071 28747
rect 15378 28744 15384 28756
rect 15059 28716 15384 28744
rect 15059 28713 15071 28716
rect 15013 28707 15071 28713
rect 15378 28704 15384 28716
rect 15436 28704 15442 28756
rect 15488 28716 17724 28744
rect 5442 28636 5448 28688
rect 5500 28676 5506 28688
rect 11330 28676 11336 28688
rect 5500 28648 9168 28676
rect 5500 28636 5506 28648
rect 7745 28611 7803 28617
rect 7745 28577 7757 28611
rect 7791 28608 7803 28611
rect 8202 28608 8208 28620
rect 7791 28580 8208 28608
rect 7791 28577 7803 28580
rect 7745 28571 7803 28577
rect 8202 28568 8208 28580
rect 8260 28568 8266 28620
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28509 6883 28543
rect 7926 28540 7932 28552
rect 7887 28512 7932 28540
rect 6825 28503 6883 28509
rect 6840 28472 6868 28503
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 9140 28549 9168 28648
rect 10980 28648 11336 28676
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28540 10471 28543
rect 10980 28540 11008 28648
rect 11330 28636 11336 28648
rect 11388 28636 11394 28688
rect 15488 28676 15516 28716
rect 14200 28648 15516 28676
rect 17696 28676 17724 28716
rect 17862 28704 17868 28756
rect 17920 28744 17926 28756
rect 20070 28744 20076 28756
rect 17920 28716 20076 28744
rect 17920 28704 17926 28716
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 20346 28704 20352 28756
rect 20404 28744 20410 28756
rect 20806 28744 20812 28756
rect 20404 28716 20812 28744
rect 20404 28704 20410 28716
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 20990 28704 20996 28756
rect 21048 28744 21054 28756
rect 21048 28716 22048 28744
rect 21048 28704 21054 28716
rect 17696 28648 20852 28676
rect 11241 28611 11299 28617
rect 11241 28577 11253 28611
rect 11287 28608 11299 28611
rect 12986 28608 12992 28620
rect 11287 28580 12992 28608
rect 11287 28577 11299 28580
rect 11241 28571 11299 28577
rect 12986 28568 12992 28580
rect 13044 28568 13050 28620
rect 10459 28512 11008 28540
rect 11057 28543 11115 28549
rect 10459 28509 10471 28512
rect 10413 28503 10471 28509
rect 11057 28509 11069 28543
rect 11103 28540 11115 28543
rect 11606 28540 11612 28552
rect 11103 28512 11612 28540
rect 11103 28509 11115 28512
rect 11057 28503 11115 28509
rect 11606 28500 11612 28512
rect 11664 28500 11670 28552
rect 12161 28543 12219 28549
rect 12161 28509 12173 28543
rect 12207 28540 12219 28543
rect 12250 28540 12256 28552
rect 12207 28512 12256 28540
rect 12207 28509 12219 28512
rect 12161 28503 12219 28509
rect 12250 28500 12256 28512
rect 12308 28500 12314 28552
rect 12802 28540 12808 28552
rect 12763 28512 12808 28540
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13722 28540 13728 28552
rect 13587 28512 13728 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 13722 28500 13728 28512
rect 13780 28540 13786 28552
rect 14200 28540 14228 28648
rect 15930 28608 15936 28620
rect 14292 28580 15936 28608
rect 14292 28549 14320 28580
rect 15930 28568 15936 28580
rect 15988 28568 15994 28620
rect 16209 28611 16267 28617
rect 16209 28577 16221 28611
rect 16255 28608 16267 28611
rect 16942 28608 16948 28620
rect 16255 28580 16948 28608
rect 16255 28577 16267 28580
rect 16209 28571 16267 28577
rect 16942 28568 16948 28580
rect 17000 28568 17006 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28577 17463 28611
rect 20346 28608 20352 28620
rect 17405 28571 17463 28577
rect 17604 28580 20352 28608
rect 13780 28512 14228 28540
rect 14277 28543 14335 28549
rect 13780 28500 13786 28512
rect 14277 28509 14289 28543
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 14918 28500 14924 28552
rect 14976 28540 14982 28552
rect 16022 28540 16028 28552
rect 14976 28512 15021 28540
rect 15983 28512 16028 28540
rect 14976 28500 14982 28512
rect 16022 28500 16028 28512
rect 16080 28500 16086 28552
rect 17420 28540 17448 28571
rect 17494 28540 17500 28552
rect 17420 28512 17500 28540
rect 17494 28500 17500 28512
rect 17552 28500 17558 28552
rect 8202 28472 8208 28484
rect 6840 28444 8208 28472
rect 8202 28432 8208 28444
rect 8260 28432 8266 28484
rect 15930 28432 15936 28484
rect 15988 28472 15994 28484
rect 17604 28472 17632 28580
rect 20346 28568 20352 28580
rect 20404 28568 20410 28620
rect 20714 28608 20720 28620
rect 20675 28580 20720 28608
rect 20714 28568 20720 28580
rect 20772 28568 20778 28620
rect 20824 28608 20852 28648
rect 21726 28608 21732 28620
rect 20824 28580 21732 28608
rect 21726 28568 21732 28580
rect 21784 28568 21790 28620
rect 22020 28608 22048 28716
rect 26878 28704 26884 28756
rect 26936 28744 26942 28756
rect 37461 28747 37519 28753
rect 26936 28716 35020 28744
rect 26936 28704 26942 28716
rect 24854 28608 24860 28620
rect 22020 28580 22968 28608
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 20438 28540 20444 28552
rect 17828 28512 20444 28540
rect 17828 28500 17834 28512
rect 20438 28500 20444 28512
rect 20496 28500 20502 28552
rect 15988 28444 17632 28472
rect 15988 28432 15994 28444
rect 17678 28432 17684 28484
rect 17736 28472 17742 28484
rect 19978 28472 19984 28484
rect 17736 28444 19984 28472
rect 17736 28432 17742 28444
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 20990 28472 20996 28484
rect 20951 28444 20996 28472
rect 20990 28432 20996 28444
rect 21048 28432 21054 28484
rect 21100 28444 21482 28472
rect 8386 28404 8392 28416
rect 8347 28376 8392 28404
rect 8386 28364 8392 28376
rect 8444 28364 8450 28416
rect 9217 28407 9275 28413
rect 9217 28373 9229 28407
rect 9263 28404 9275 28407
rect 11146 28404 11152 28416
rect 9263 28376 11152 28404
rect 9263 28373 9275 28376
rect 9217 28367 9275 28373
rect 11146 28364 11152 28376
rect 11204 28364 11210 28416
rect 12253 28407 12311 28413
rect 12253 28373 12265 28407
rect 12299 28404 12311 28407
rect 12342 28404 12348 28416
rect 12299 28376 12348 28404
rect 12299 28373 12311 28376
rect 12253 28367 12311 28373
rect 12342 28364 12348 28376
rect 12400 28364 12406 28416
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 21100 28404 21128 28444
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 22741 28475 22799 28481
rect 22741 28472 22753 28475
rect 22612 28444 22753 28472
rect 22612 28432 22618 28444
rect 22741 28441 22753 28444
rect 22787 28441 22799 28475
rect 22940 28472 22968 28580
rect 24596 28580 24860 28608
rect 23014 28500 23020 28552
rect 23072 28540 23078 28552
rect 24596 28549 24624 28580
rect 24854 28568 24860 28580
rect 24912 28568 24918 28620
rect 26142 28568 26148 28620
rect 26200 28608 26206 28620
rect 26329 28611 26387 28617
rect 26329 28608 26341 28611
rect 26200 28580 26341 28608
rect 26200 28568 26206 28580
rect 26329 28577 26341 28580
rect 26375 28577 26387 28611
rect 26329 28571 26387 28577
rect 26694 28568 26700 28620
rect 26752 28608 26758 28620
rect 31389 28611 31447 28617
rect 31389 28608 31401 28611
rect 26752 28580 31401 28608
rect 26752 28568 26758 28580
rect 31389 28577 31401 28580
rect 31435 28577 31447 28611
rect 34992 28608 35020 28716
rect 37461 28713 37473 28747
rect 37507 28744 37519 28747
rect 37550 28744 37556 28756
rect 37507 28716 37556 28744
rect 37507 28713 37519 28716
rect 37461 28707 37519 28713
rect 37550 28704 37556 28716
rect 37608 28704 37614 28756
rect 34992 28580 38332 28608
rect 31389 28571 31447 28577
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 23072 28512 24593 28540
rect 23072 28500 23078 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 27614 28500 27620 28552
rect 27672 28540 27678 28552
rect 28813 28543 28871 28549
rect 28813 28540 28825 28543
rect 27672 28512 28825 28540
rect 27672 28500 27678 28512
rect 28813 28509 28825 28512
rect 28859 28509 28871 28543
rect 31110 28540 31116 28552
rect 31071 28512 31116 28540
rect 28813 28503 28871 28509
rect 31110 28500 31116 28512
rect 31168 28500 31174 28552
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34848 28512 34897 28540
rect 34848 28500 34854 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 37642 28540 37648 28552
rect 37603 28512 37648 28540
rect 34885 28503 34943 28509
rect 37642 28500 37648 28512
rect 37700 28500 37706 28552
rect 38304 28549 38332 28580
rect 38289 28543 38347 28549
rect 38289 28509 38301 28543
rect 38335 28509 38347 28543
rect 38289 28503 38347 28509
rect 24857 28475 24915 28481
rect 24857 28472 24869 28475
rect 22940 28444 24869 28472
rect 22741 28435 22799 28441
rect 24857 28441 24869 28444
rect 24903 28441 24915 28475
rect 24857 28435 24915 28441
rect 25314 28432 25320 28484
rect 25372 28432 25378 28484
rect 28074 28472 28080 28484
rect 28035 28444 28080 28472
rect 28074 28432 28080 28444
rect 28132 28432 28138 28484
rect 32030 28432 32036 28484
rect 32088 28432 32094 28484
rect 32784 28444 33088 28472
rect 15252 28376 21128 28404
rect 15252 28364 15258 28376
rect 21726 28364 21732 28416
rect 21784 28404 21790 28416
rect 31662 28404 31668 28416
rect 21784 28376 31668 28404
rect 21784 28364 21790 28376
rect 31662 28364 31668 28376
rect 31720 28404 31726 28416
rect 32784 28404 32812 28444
rect 31720 28376 32812 28404
rect 31720 28364 31726 28376
rect 32858 28364 32864 28416
rect 32916 28404 32922 28416
rect 33060 28404 33088 28444
rect 34054 28432 34060 28484
rect 34112 28472 34118 28484
rect 35161 28475 35219 28481
rect 35161 28472 35173 28475
rect 34112 28444 35173 28472
rect 34112 28432 34118 28444
rect 35161 28441 35173 28444
rect 35207 28441 35219 28475
rect 38654 28472 38660 28484
rect 36386 28444 38660 28472
rect 35161 28435 35219 28441
rect 38654 28432 38660 28444
rect 38712 28432 38718 28484
rect 36633 28407 36691 28413
rect 36633 28404 36645 28407
rect 32916 28376 32961 28404
rect 33060 28376 36645 28404
rect 32916 28364 32922 28376
rect 36633 28373 36645 28376
rect 36679 28373 36691 28407
rect 36633 28367 36691 28373
rect 38010 28364 38016 28416
rect 38068 28404 38074 28416
rect 38105 28407 38163 28413
rect 38105 28404 38117 28407
rect 38068 28376 38117 28404
rect 38068 28364 38074 28376
rect 38105 28373 38117 28376
rect 38151 28373 38163 28407
rect 38105 28367 38163 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 7561 28203 7619 28209
rect 7561 28169 7573 28203
rect 7607 28200 7619 28203
rect 7926 28200 7932 28212
rect 7607 28172 7932 28200
rect 7607 28169 7619 28172
rect 7561 28163 7619 28169
rect 7926 28160 7932 28172
rect 7984 28160 7990 28212
rect 8202 28200 8208 28212
rect 8163 28172 8208 28200
rect 8202 28160 8208 28172
rect 8260 28160 8266 28212
rect 23934 28200 23940 28212
rect 8312 28172 23940 28200
rect 6917 28135 6975 28141
rect 6917 28101 6929 28135
rect 6963 28132 6975 28135
rect 7742 28132 7748 28144
rect 6963 28104 7748 28132
rect 6963 28101 6975 28104
rect 6917 28095 6975 28101
rect 7742 28092 7748 28104
rect 7800 28092 7806 28144
rect 8312 28132 8340 28172
rect 23934 28160 23940 28172
rect 23992 28160 23998 28212
rect 24026 28160 24032 28212
rect 24084 28200 24090 28212
rect 36446 28200 36452 28212
rect 24084 28172 36452 28200
rect 24084 28160 24090 28172
rect 36446 28160 36452 28172
rect 36504 28160 36510 28212
rect 8036 28104 8340 28132
rect 6822 28064 6828 28076
rect 6783 28036 6828 28064
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 7098 28024 7104 28076
rect 7156 28064 7162 28076
rect 7469 28067 7527 28073
rect 7469 28064 7481 28067
rect 7156 28036 7481 28064
rect 7156 28024 7162 28036
rect 7469 28033 7481 28036
rect 7515 28064 7527 28067
rect 8036 28064 8064 28104
rect 10042 28092 10048 28144
rect 10100 28132 10106 28144
rect 10137 28135 10195 28141
rect 10137 28132 10149 28135
rect 10100 28104 10149 28132
rect 10100 28092 10106 28104
rect 10137 28101 10149 28104
rect 10183 28101 10195 28135
rect 10137 28095 10195 28101
rect 11057 28135 11115 28141
rect 11057 28101 11069 28135
rect 11103 28132 11115 28135
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 11103 28104 11897 28132
rect 11103 28101 11115 28104
rect 11057 28095 11115 28101
rect 11885 28101 11897 28104
rect 11931 28101 11943 28135
rect 13906 28132 13912 28144
rect 11885 28095 11943 28101
rect 13280 28104 13912 28132
rect 7515 28036 8064 28064
rect 8113 28067 8171 28073
rect 7515 28033 7527 28036
rect 7469 28027 7527 28033
rect 8113 28033 8125 28067
rect 8159 28064 8171 28067
rect 9766 28064 9772 28076
rect 8159 28036 9772 28064
rect 8159 28033 8171 28036
rect 8113 28027 8171 28033
rect 9766 28024 9772 28036
rect 9824 28024 9830 28076
rect 10778 28024 10784 28076
rect 10836 28064 10842 28076
rect 10965 28067 11023 28073
rect 10965 28064 10977 28067
rect 10836 28036 10977 28064
rect 10836 28024 10842 28036
rect 10965 28033 10977 28036
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 10502 27956 10508 28008
rect 10560 27996 10566 28008
rect 11793 27999 11851 28005
rect 11793 27996 11805 27999
rect 10560 27968 11805 27996
rect 10560 27956 10566 27968
rect 11793 27965 11805 27968
rect 11839 27965 11851 27999
rect 11793 27959 11851 27965
rect 12434 27956 12440 28008
rect 12492 27996 12498 28008
rect 13280 27996 13308 28104
rect 13906 28092 13912 28104
rect 13964 28092 13970 28144
rect 14182 28132 14188 28144
rect 14143 28104 14188 28132
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 15378 28132 15384 28144
rect 15339 28104 15384 28132
rect 15378 28092 15384 28104
rect 15436 28092 15442 28144
rect 19518 28092 19524 28144
rect 19576 28092 19582 28144
rect 20257 28135 20315 28141
rect 20257 28101 20269 28135
rect 20303 28132 20315 28135
rect 20438 28132 20444 28144
rect 20303 28104 20444 28132
rect 20303 28101 20315 28104
rect 20257 28095 20315 28101
rect 20438 28092 20444 28104
rect 20496 28092 20502 28144
rect 26050 28132 26056 28144
rect 24334 28104 26056 28132
rect 26050 28092 26056 28104
rect 26108 28092 26114 28144
rect 29730 28092 29736 28144
rect 29788 28132 29794 28144
rect 33321 28135 33379 28141
rect 33321 28132 33333 28135
rect 29788 28104 33333 28132
rect 29788 28092 29794 28104
rect 33321 28101 33333 28104
rect 33367 28132 33379 28135
rect 33410 28132 33416 28144
rect 33367 28104 33416 28132
rect 33367 28101 33379 28104
rect 33321 28095 33379 28101
rect 33410 28092 33416 28104
rect 33468 28092 33474 28144
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 12492 27968 13308 27996
rect 12492 27956 12498 27968
rect 10318 27928 10324 27940
rect 10279 27900 10324 27928
rect 10318 27888 10324 27900
rect 10376 27888 10382 27940
rect 10870 27888 10876 27940
rect 10928 27928 10934 27940
rect 13372 27928 13400 28027
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 22833 28067 22891 28073
rect 22833 28064 22845 28067
rect 20772 28036 22845 28064
rect 20772 28024 20778 28036
rect 22833 28033 22845 28036
rect 22879 28033 22891 28067
rect 31294 28064 31300 28076
rect 29026 28036 31300 28064
rect 22833 28027 22891 28033
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 36170 28024 36176 28076
rect 36228 28064 36234 28076
rect 37737 28067 37795 28073
rect 37737 28064 37749 28067
rect 36228 28036 37749 28064
rect 36228 28024 36234 28036
rect 37737 28033 37749 28036
rect 37783 28033 37795 28067
rect 37737 28027 37795 28033
rect 14093 27999 14151 28005
rect 14093 27965 14105 27999
rect 14139 27996 14151 27999
rect 14366 27996 14372 28008
rect 14139 27968 14372 27996
rect 14139 27965 14151 27968
rect 14093 27959 14151 27965
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 14550 27996 14556 28008
rect 14511 27968 14556 27996
rect 14550 27956 14556 27968
rect 14608 27956 14614 28008
rect 15289 27999 15347 28005
rect 15289 27965 15301 27999
rect 15335 27996 15347 27999
rect 15746 27996 15752 28008
rect 15335 27968 15752 27996
rect 15335 27965 15347 27968
rect 15289 27959 15347 27965
rect 15746 27956 15752 27968
rect 15804 27956 15810 28008
rect 16206 27996 16212 28008
rect 16167 27968 16212 27996
rect 16206 27956 16212 27968
rect 16264 27956 16270 28008
rect 18138 27956 18144 28008
rect 18196 27996 18202 28008
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 18196 27968 18245 27996
rect 18196 27956 18202 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 18509 27999 18567 28005
rect 18509 27996 18521 27999
rect 18233 27959 18291 27965
rect 18340 27968 18521 27996
rect 10928 27900 13400 27928
rect 13449 27931 13507 27937
rect 10928 27888 10934 27900
rect 13449 27897 13461 27931
rect 13495 27928 13507 27931
rect 15654 27928 15660 27940
rect 13495 27900 15660 27928
rect 13495 27897 13507 27900
rect 13449 27891 13507 27897
rect 15654 27888 15660 27900
rect 15712 27888 15718 27940
rect 15838 27888 15844 27940
rect 15896 27928 15902 27940
rect 18340 27928 18368 27968
rect 18509 27965 18521 27968
rect 18555 27996 18567 27999
rect 21082 27996 21088 28008
rect 18555 27968 21088 27996
rect 18555 27965 18567 27968
rect 18509 27959 18567 27965
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 23109 27999 23167 28005
rect 23109 27996 23121 27999
rect 22848 27968 23121 27996
rect 22848 27940 22876 27968
rect 23109 27965 23121 27968
rect 23155 27965 23167 27999
rect 27614 27996 27620 28008
rect 27575 27968 27620 27996
rect 23109 27959 23167 27965
rect 27614 27956 27620 27968
rect 27672 27956 27678 28008
rect 27893 27999 27951 28005
rect 27893 27965 27905 27999
rect 27939 27996 27951 27999
rect 28902 27996 28908 28008
rect 27939 27968 28908 27996
rect 27939 27965 27951 27968
rect 27893 27959 27951 27965
rect 28902 27956 28908 27968
rect 28960 27996 28966 28008
rect 29638 27996 29644 28008
rect 28960 27968 29644 27996
rect 28960 27956 28966 27968
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 31110 27956 31116 28008
rect 31168 27996 31174 28008
rect 31662 27996 31668 28008
rect 31168 27968 31668 27996
rect 31168 27956 31174 27968
rect 31662 27956 31668 27968
rect 31720 27996 31726 28008
rect 34057 27999 34115 28005
rect 34057 27996 34069 27999
rect 31720 27968 34069 27996
rect 31720 27956 31726 27968
rect 34057 27965 34069 27968
rect 34103 27996 34115 27999
rect 34790 27996 34796 28008
rect 34103 27968 34796 27996
rect 34103 27965 34115 27968
rect 34057 27959 34115 27965
rect 34790 27956 34796 27968
rect 34848 27956 34854 28008
rect 15896 27900 18368 27928
rect 15896 27888 15902 27900
rect 22830 27888 22836 27940
rect 22888 27888 22894 27940
rect 26234 27928 26240 27940
rect 24136 27900 26240 27928
rect 12894 27820 12900 27872
rect 12952 27860 12958 27872
rect 24136 27860 24164 27900
rect 26234 27888 26240 27900
rect 26292 27888 26298 27940
rect 12952 27832 24164 27860
rect 24581 27863 24639 27869
rect 12952 27820 12958 27832
rect 24581 27829 24593 27863
rect 24627 27860 24639 27863
rect 24946 27860 24952 27872
rect 24627 27832 24952 27860
rect 24627 27829 24639 27832
rect 24581 27823 24639 27829
rect 24946 27820 24952 27832
rect 25004 27820 25010 27872
rect 25038 27820 25044 27872
rect 25096 27860 25102 27872
rect 26970 27860 26976 27872
rect 25096 27832 26976 27860
rect 25096 27820 25102 27832
rect 26970 27820 26976 27832
rect 27028 27820 27034 27872
rect 29362 27860 29368 27872
rect 29323 27832 29368 27860
rect 29362 27820 29368 27832
rect 29420 27820 29426 27872
rect 33410 27820 33416 27872
rect 33468 27860 33474 27872
rect 37829 27863 37887 27869
rect 37829 27860 37841 27863
rect 33468 27832 37841 27860
rect 33468 27820 33474 27832
rect 37829 27829 37841 27832
rect 37875 27829 37887 27863
rect 37829 27823 37887 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 10410 27616 10416 27668
rect 10468 27656 10474 27668
rect 10870 27656 10876 27668
rect 10468 27628 10876 27656
rect 10468 27616 10474 27628
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 14200 27628 14412 27656
rect 9674 27588 9680 27600
rect 9635 27560 9680 27588
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 13633 27591 13691 27597
rect 13633 27557 13645 27591
rect 13679 27588 13691 27591
rect 14200 27588 14228 27628
rect 13679 27560 14228 27588
rect 14277 27591 14335 27597
rect 13679 27557 13691 27560
rect 13633 27551 13691 27557
rect 14277 27557 14289 27591
rect 14323 27557 14335 27591
rect 14384 27588 14412 27628
rect 14734 27616 14740 27668
rect 14792 27656 14798 27668
rect 25314 27656 25320 27668
rect 14792 27628 25320 27656
rect 14792 27616 14798 27628
rect 25314 27616 25320 27628
rect 25372 27616 25378 27668
rect 27706 27616 27712 27668
rect 27764 27656 27770 27668
rect 28350 27656 28356 27668
rect 27764 27628 28356 27656
rect 27764 27616 27770 27628
rect 28350 27616 28356 27628
rect 28408 27616 28414 27668
rect 31386 27616 31392 27668
rect 31444 27656 31450 27668
rect 32198 27659 32256 27665
rect 32198 27656 32210 27659
rect 31444 27628 32210 27656
rect 31444 27616 31450 27628
rect 32198 27625 32210 27628
rect 32244 27625 32256 27659
rect 32198 27619 32256 27625
rect 32858 27616 32864 27668
rect 32916 27656 32922 27668
rect 35142 27659 35200 27665
rect 35142 27656 35154 27659
rect 32916 27628 35154 27656
rect 32916 27616 32922 27628
rect 35142 27625 35154 27628
rect 35188 27625 35200 27659
rect 35142 27619 35200 27625
rect 23382 27588 23388 27600
rect 14384 27560 23388 27588
rect 14277 27551 14335 27557
rect 11146 27480 11152 27532
rect 11204 27520 11210 27532
rect 11885 27523 11943 27529
rect 11885 27520 11897 27523
rect 11204 27492 11897 27520
rect 11204 27480 11210 27492
rect 11885 27489 11897 27492
rect 11931 27489 11943 27523
rect 14292 27520 14320 27551
rect 23382 27548 23388 27560
rect 23440 27548 23446 27600
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 26421 27591 26479 27597
rect 26421 27588 26433 27591
rect 26384 27560 26433 27588
rect 26384 27548 26390 27560
rect 26421 27557 26433 27560
rect 26467 27557 26479 27591
rect 26421 27551 26479 27557
rect 31036 27560 32076 27588
rect 24394 27520 24400 27532
rect 14292 27492 24400 27520
rect 11885 27483 11943 27489
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 27341 27523 27399 27529
rect 27341 27489 27353 27523
rect 27387 27520 27399 27523
rect 27614 27520 27620 27532
rect 27387 27492 27620 27520
rect 27387 27489 27399 27492
rect 27341 27483 27399 27489
rect 27614 27480 27620 27492
rect 27672 27480 27678 27532
rect 30006 27480 30012 27532
rect 30064 27520 30070 27532
rect 31036 27520 31064 27560
rect 30064 27492 31064 27520
rect 31481 27523 31539 27529
rect 30064 27480 30070 27492
rect 31481 27489 31493 27523
rect 31527 27489 31539 27523
rect 31481 27483 31539 27489
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 9214 27412 9220 27464
rect 9272 27452 9278 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 9272 27424 9873 27452
rect 9272 27412 9278 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 10321 27455 10379 27461
rect 10321 27421 10333 27455
rect 10367 27452 10379 27455
rect 10594 27452 10600 27464
rect 10367 27424 10600 27452
rect 10367 27421 10379 27424
rect 10321 27415 10379 27421
rect 10594 27412 10600 27424
rect 10652 27412 10658 27464
rect 12802 27412 12808 27464
rect 12860 27452 12866 27464
rect 13541 27455 13599 27461
rect 13541 27452 13553 27455
rect 12860 27424 13553 27452
rect 12860 27412 12866 27424
rect 13541 27421 13553 27424
rect 13587 27452 13599 27455
rect 13998 27452 14004 27464
rect 13587 27424 14004 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 13998 27412 14004 27424
rect 14056 27412 14062 27464
rect 14274 27412 14280 27464
rect 14332 27452 14338 27464
rect 14461 27455 14519 27461
rect 14461 27452 14473 27455
rect 14332 27424 14473 27452
rect 14332 27412 14338 27424
rect 14461 27421 14473 27424
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 15105 27455 15163 27461
rect 15105 27421 15117 27455
rect 15151 27421 15163 27455
rect 15105 27415 15163 27421
rect 11974 27344 11980 27396
rect 12032 27384 12038 27396
rect 12526 27384 12532 27396
rect 12032 27356 12077 27384
rect 12487 27356 12532 27384
rect 12032 27344 12038 27356
rect 12526 27344 12532 27356
rect 12584 27344 12590 27396
rect 14016 27384 14044 27412
rect 15120 27384 15148 27415
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 15252 27424 15297 27452
rect 15252 27412 15258 27424
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 24636 27424 24685 27452
rect 24636 27412 24642 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 28902 27412 28908 27464
rect 28960 27452 28966 27464
rect 29733 27455 29791 27461
rect 29733 27452 29745 27455
rect 28960 27424 29745 27452
rect 28960 27412 28966 27424
rect 29733 27421 29745 27424
rect 29779 27421 29791 27455
rect 31496 27452 31524 27483
rect 31662 27480 31668 27532
rect 31720 27520 31726 27532
rect 31941 27523 31999 27529
rect 31941 27520 31953 27523
rect 31720 27492 31953 27520
rect 31720 27480 31726 27492
rect 31941 27489 31953 27492
rect 31987 27489 31999 27523
rect 32048 27520 32076 27560
rect 33689 27523 33747 27529
rect 33689 27520 33701 27523
rect 32048 27492 33701 27520
rect 31941 27483 31999 27489
rect 33689 27489 33701 27492
rect 33735 27489 33747 27523
rect 33689 27483 33747 27489
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 34885 27523 34943 27529
rect 34885 27520 34897 27523
rect 34848 27492 34897 27520
rect 34848 27480 34854 27492
rect 34885 27489 34897 27492
rect 34931 27489 34943 27523
rect 34885 27483 34943 27489
rect 31754 27452 31760 27464
rect 31496 27424 31760 27452
rect 29733 27415 29791 27421
rect 31754 27412 31760 27424
rect 31812 27412 31818 27464
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 37660 27424 38025 27452
rect 14016 27356 15148 27384
rect 15841 27387 15899 27393
rect 15841 27353 15853 27387
rect 15887 27353 15899 27387
rect 15841 27347 15899 27353
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 6822 27316 6828 27328
rect 1627 27288 6828 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 10410 27316 10416 27328
rect 10371 27288 10416 27316
rect 10410 27276 10416 27288
rect 10468 27276 10474 27328
rect 12158 27276 12164 27328
rect 12216 27316 12222 27328
rect 15856 27316 15884 27347
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 16850 27384 16856 27396
rect 15988 27356 16033 27384
rect 16811 27356 16856 27384
rect 15988 27344 15994 27356
rect 16850 27344 16856 27356
rect 16908 27344 16914 27396
rect 20070 27344 20076 27396
rect 20128 27384 20134 27396
rect 23290 27384 23296 27396
rect 20128 27356 23296 27384
rect 20128 27344 20134 27356
rect 23290 27344 23296 27356
rect 23348 27344 23354 27396
rect 24949 27387 25007 27393
rect 24949 27353 24961 27387
rect 24995 27384 25007 27387
rect 25038 27384 25044 27396
rect 24995 27356 25044 27384
rect 24995 27353 25007 27356
rect 24949 27347 25007 27353
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 25682 27344 25688 27396
rect 25740 27344 25746 27396
rect 27617 27387 27675 27393
rect 27617 27353 27629 27387
rect 27663 27384 27675 27387
rect 27706 27384 27712 27396
rect 27663 27356 27712 27384
rect 27663 27353 27675 27356
rect 27617 27347 27675 27353
rect 27706 27344 27712 27356
rect 27764 27344 27770 27396
rect 28842 27356 29960 27384
rect 16758 27316 16764 27328
rect 12216 27288 16764 27316
rect 12216 27276 12222 27288
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 20622 27276 20628 27328
rect 20680 27316 20686 27328
rect 29086 27316 29092 27328
rect 20680 27288 29092 27316
rect 20680 27276 20686 27288
rect 29086 27276 29092 27288
rect 29144 27276 29150 27328
rect 29932 27316 29960 27356
rect 30006 27344 30012 27396
rect 30064 27384 30070 27396
rect 31478 27384 31484 27396
rect 30064 27356 30109 27384
rect 31234 27356 31484 27384
rect 30064 27344 30070 27356
rect 31478 27344 31484 27356
rect 31536 27344 31542 27396
rect 37550 27384 37556 27396
rect 33442 27356 34100 27384
rect 36386 27356 37556 27384
rect 33226 27316 33232 27328
rect 29932 27288 33232 27316
rect 33226 27276 33232 27288
rect 33284 27276 33290 27328
rect 34072 27316 34100 27356
rect 37550 27344 37556 27356
rect 37608 27344 37614 27396
rect 37660 27328 37688 27424
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 35894 27316 35900 27328
rect 34072 27288 35900 27316
rect 35894 27276 35900 27288
rect 35952 27276 35958 27328
rect 36630 27316 36636 27328
rect 36591 27288 36636 27316
rect 36630 27276 36636 27288
rect 36688 27276 36694 27328
rect 37642 27316 37648 27328
rect 37603 27288 37648 27316
rect 37642 27276 37648 27288
rect 37700 27276 37706 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 9214 27112 9220 27124
rect 9175 27084 9220 27112
rect 9214 27072 9220 27084
rect 9272 27072 9278 27124
rect 13633 27115 13691 27121
rect 13633 27081 13645 27115
rect 13679 27112 13691 27115
rect 14182 27112 14188 27124
rect 13679 27084 14188 27112
rect 13679 27081 13691 27084
rect 13633 27075 13691 27081
rect 14182 27072 14188 27084
rect 14240 27072 14246 27124
rect 23014 27112 23020 27124
rect 22020 27084 23020 27112
rect 15194 27004 15200 27056
rect 15252 27044 15258 27056
rect 15252 27016 18906 27044
rect 15252 27004 15258 27016
rect 9398 26976 9404 26988
rect 9359 26948 9404 26976
rect 9398 26936 9404 26948
rect 9456 26936 9462 26988
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26976 11023 26979
rect 11146 26976 11152 26988
rect 11011 26948 11152 26976
rect 11011 26945 11023 26948
rect 10965 26939 11023 26945
rect 11146 26936 11152 26948
rect 11204 26936 11210 26988
rect 11974 26976 11980 26988
rect 11935 26948 11980 26976
rect 11974 26936 11980 26948
rect 12032 26936 12038 26988
rect 12621 26979 12679 26985
rect 12621 26945 12633 26979
rect 12667 26976 12679 26979
rect 12710 26976 12716 26988
rect 12667 26948 12716 26976
rect 12667 26945 12679 26948
rect 12621 26939 12679 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 13538 26936 13544 26988
rect 13596 26976 13602 26988
rect 13817 26979 13875 26985
rect 13817 26976 13829 26979
rect 13596 26948 13829 26976
rect 13596 26936 13602 26948
rect 13817 26945 13829 26948
rect 13863 26945 13875 26979
rect 18138 26976 18144 26988
rect 18099 26948 18144 26976
rect 13817 26939 13875 26945
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 22020 26985 22048 27084
rect 23014 27072 23020 27084
rect 23072 27112 23078 27124
rect 23072 27084 24256 27112
rect 23072 27072 23078 27084
rect 23658 27044 23664 27056
rect 23506 27016 23664 27044
rect 23658 27004 23664 27016
rect 23716 27004 23722 27056
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26945 22063 26979
rect 24228 26976 24256 27084
rect 24578 27072 24584 27124
rect 24636 27112 24642 27124
rect 27614 27112 27620 27124
rect 24636 27084 27620 27112
rect 24636 27072 24642 27084
rect 25130 27044 25136 27056
rect 25091 27016 25136 27044
rect 25130 27004 25136 27016
rect 25188 27004 25194 27056
rect 26510 27044 26516 27056
rect 26358 27016 26516 27044
rect 26510 27004 26516 27016
rect 26568 27004 26574 27056
rect 27172 26985 27200 27084
rect 27614 27072 27620 27084
rect 27672 27112 27678 27124
rect 28902 27112 28908 27124
rect 27672 27084 28908 27112
rect 27672 27072 27678 27084
rect 28902 27072 28908 27084
rect 28960 27112 28966 27124
rect 28960 27084 29500 27112
rect 28960 27072 28966 27084
rect 27890 27004 27896 27056
rect 27948 27004 27954 27056
rect 29472 26985 29500 27084
rect 30650 27072 30656 27124
rect 30708 27112 30714 27124
rect 36630 27112 36636 27124
rect 30708 27084 36636 27112
rect 30708 27072 30714 27084
rect 36630 27072 36636 27084
rect 36688 27072 36694 27124
rect 31018 27044 31024 27056
rect 30958 27016 31024 27044
rect 31018 27004 31024 27016
rect 31076 27004 31082 27056
rect 34422 27044 34428 27056
rect 34362 27016 34428 27044
rect 34422 27004 34428 27016
rect 34480 27004 34486 27056
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24228 26948 24869 26976
rect 22005 26939 22063 26945
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26945 29515 26979
rect 29457 26939 29515 26945
rect 31662 26936 31668 26988
rect 31720 26976 31726 26988
rect 32861 26979 32919 26985
rect 32861 26976 32873 26979
rect 31720 26948 32873 26976
rect 31720 26936 31726 26948
rect 32861 26945 32873 26948
rect 32907 26945 32919 26979
rect 32861 26939 32919 26945
rect 15102 26868 15108 26920
rect 15160 26908 15166 26920
rect 18417 26911 18475 26917
rect 18417 26908 18429 26911
rect 15160 26880 18429 26908
rect 15160 26868 15166 26880
rect 18417 26877 18429 26880
rect 18463 26908 18475 26911
rect 19150 26908 19156 26920
rect 18463 26880 19156 26908
rect 18463 26877 18475 26880
rect 18417 26871 18475 26877
rect 19150 26868 19156 26880
rect 19208 26868 19214 26920
rect 19426 26868 19432 26920
rect 19484 26908 19490 26920
rect 20165 26911 20223 26917
rect 20165 26908 20177 26911
rect 19484 26880 20177 26908
rect 19484 26868 19490 26880
rect 20165 26877 20177 26880
rect 20211 26908 20223 26911
rect 20990 26908 20996 26920
rect 20211 26880 20996 26908
rect 20211 26877 20223 26880
rect 20165 26871 20223 26877
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 22281 26911 22339 26917
rect 22281 26877 22293 26911
rect 22327 26908 22339 26911
rect 22370 26908 22376 26920
rect 22327 26880 22376 26908
rect 22327 26877 22339 26880
rect 22281 26871 22339 26877
rect 22370 26868 22376 26880
rect 22428 26868 22434 26920
rect 23290 26868 23296 26920
rect 23348 26908 23354 26920
rect 24029 26911 24087 26917
rect 24029 26908 24041 26911
rect 23348 26880 24041 26908
rect 23348 26868 23354 26880
rect 24029 26877 24041 26880
rect 24075 26877 24087 26911
rect 25866 26908 25872 26920
rect 24029 26871 24087 26877
rect 24320 26880 25872 26908
rect 11057 26843 11115 26849
rect 11057 26809 11069 26843
rect 11103 26840 11115 26843
rect 11103 26812 17264 26840
rect 11103 26809 11115 26812
rect 11057 26803 11115 26809
rect 12066 26772 12072 26784
rect 12027 26744 12072 26772
rect 12066 26732 12072 26744
rect 12124 26732 12130 26784
rect 12710 26772 12716 26784
rect 12671 26744 12716 26772
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 17236 26772 17264 26812
rect 24320 26772 24348 26880
rect 25866 26868 25872 26880
rect 25924 26868 25930 26920
rect 26326 26868 26332 26920
rect 26384 26908 26390 26920
rect 27433 26911 27491 26917
rect 27433 26908 27445 26911
rect 26384 26880 27445 26908
rect 26384 26868 26390 26880
rect 27433 26877 27445 26880
rect 27479 26877 27491 26911
rect 27433 26871 27491 26877
rect 28994 26868 29000 26920
rect 29052 26908 29058 26920
rect 29362 26908 29368 26920
rect 29052 26880 29368 26908
rect 29052 26868 29058 26880
rect 29362 26868 29368 26880
rect 29420 26908 29426 26920
rect 29733 26911 29791 26917
rect 29733 26908 29745 26911
rect 29420 26880 29745 26908
rect 29420 26868 29426 26880
rect 29733 26877 29745 26880
rect 29779 26877 29791 26911
rect 29733 26871 29791 26877
rect 29822 26868 29828 26920
rect 29880 26908 29886 26920
rect 31754 26908 31760 26920
rect 29880 26880 31760 26908
rect 29880 26868 29886 26880
rect 31754 26868 31760 26880
rect 31812 26868 31818 26920
rect 33137 26911 33195 26917
rect 33137 26877 33149 26911
rect 33183 26908 33195 26911
rect 33594 26908 33600 26920
rect 33183 26880 33600 26908
rect 33183 26877 33195 26880
rect 33137 26871 33195 26877
rect 33594 26868 33600 26880
rect 33652 26868 33658 26920
rect 27062 26840 27068 26852
rect 26160 26812 27068 26840
rect 17236 26744 24348 26772
rect 24394 26732 24400 26784
rect 24452 26772 24458 26784
rect 26160 26772 26188 26812
rect 27062 26800 27068 26812
rect 27120 26800 27126 26852
rect 24452 26744 26188 26772
rect 26605 26775 26663 26781
rect 24452 26732 24458 26744
rect 26605 26741 26617 26775
rect 26651 26772 26663 26775
rect 26694 26772 26700 26784
rect 26651 26744 26700 26772
rect 26651 26741 26663 26744
rect 26605 26735 26663 26741
rect 26694 26732 26700 26744
rect 26752 26732 26758 26784
rect 28902 26772 28908 26784
rect 28863 26744 28908 26772
rect 28902 26732 28908 26744
rect 28960 26732 28966 26784
rect 31202 26772 31208 26784
rect 31163 26744 31208 26772
rect 31202 26732 31208 26744
rect 31260 26732 31266 26784
rect 34609 26775 34667 26781
rect 34609 26741 34621 26775
rect 34655 26772 34667 26775
rect 34698 26772 34704 26784
rect 34655 26744 34704 26772
rect 34655 26741 34667 26744
rect 34609 26735 34667 26741
rect 34698 26732 34704 26744
rect 34756 26732 34762 26784
rect 35434 26732 35440 26784
rect 35492 26772 35498 26784
rect 38194 26772 38200 26784
rect 35492 26744 38200 26772
rect 35492 26732 35498 26744
rect 38194 26732 38200 26744
rect 38252 26732 38258 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 9766 26568 9772 26580
rect 9727 26540 9772 26568
rect 9766 26528 9772 26540
rect 9824 26528 9830 26580
rect 13538 26568 13544 26580
rect 13499 26540 13544 26568
rect 13538 26528 13544 26540
rect 13596 26528 13602 26580
rect 15562 26568 15568 26580
rect 15523 26540 15568 26568
rect 15562 26528 15568 26540
rect 15620 26528 15626 26580
rect 17954 26528 17960 26580
rect 18012 26568 18018 26580
rect 21453 26571 21511 26577
rect 21453 26568 21465 26571
rect 18012 26540 21465 26568
rect 18012 26528 18018 26540
rect 21453 26537 21465 26540
rect 21499 26537 21511 26571
rect 24854 26568 24860 26580
rect 21453 26531 21511 26537
rect 22066 26540 24860 26568
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 6730 26500 6736 26512
rect 1627 26472 6736 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 6730 26460 6736 26472
rect 6788 26460 6794 26512
rect 11974 26460 11980 26512
rect 12032 26500 12038 26512
rect 19334 26500 19340 26512
rect 12032 26472 19340 26500
rect 12032 26460 12038 26472
rect 19334 26460 19340 26472
rect 19392 26460 19398 26512
rect 22066 26500 22094 26540
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 25314 26528 25320 26580
rect 25372 26568 25378 26580
rect 28994 26568 29000 26580
rect 25372 26540 29000 26568
rect 25372 26528 25378 26540
rect 28994 26528 29000 26540
rect 29052 26528 29058 26580
rect 29178 26528 29184 26580
rect 29236 26568 29242 26580
rect 36633 26571 36691 26577
rect 36633 26568 36645 26571
rect 29236 26540 36645 26568
rect 29236 26528 29242 26540
rect 36633 26537 36645 26540
rect 36679 26537 36691 26571
rect 36633 26531 36691 26537
rect 21008 26472 22094 26500
rect 10318 26392 10324 26444
rect 10376 26432 10382 26444
rect 14366 26432 14372 26444
rect 10376 26404 13676 26432
rect 14327 26404 14372 26432
rect 10376 26392 10382 26404
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8435 26336 9137 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9306 26364 9312 26376
rect 9267 26336 9312 26364
rect 9125 26327 9183 26333
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 10318 26296 10324 26308
rect 10279 26268 10324 26296
rect 10318 26256 10324 26268
rect 10376 26256 10382 26308
rect 10410 26256 10416 26308
rect 10468 26296 10474 26308
rect 11333 26299 11391 26305
rect 10468 26268 10513 26296
rect 10468 26256 10474 26268
rect 11333 26265 11345 26299
rect 11379 26296 11391 26299
rect 12434 26296 12440 26308
rect 11379 26268 12440 26296
rect 11379 26265 11391 26268
rect 11333 26259 11391 26265
rect 12434 26256 12440 26268
rect 12492 26256 12498 26308
rect 13648 26228 13676 26404
rect 14366 26392 14372 26404
rect 14424 26392 14430 26444
rect 14458 26392 14464 26444
rect 14516 26432 14522 26444
rect 14645 26435 14703 26441
rect 14645 26432 14657 26435
rect 14516 26404 14657 26432
rect 14516 26392 14522 26404
rect 14645 26401 14657 26404
rect 14691 26401 14703 26435
rect 21008 26432 21036 26472
rect 25866 26460 25872 26512
rect 25924 26500 25930 26512
rect 30374 26500 30380 26512
rect 25924 26472 30380 26500
rect 25924 26460 25930 26472
rect 30374 26460 30380 26472
rect 30432 26460 30438 26512
rect 38930 26500 38936 26512
rect 34716 26472 35020 26500
rect 23014 26432 23020 26444
rect 14645 26395 14703 26401
rect 15488 26404 21036 26432
rect 21100 26404 23020 26432
rect 13722 26324 13728 26376
rect 13780 26364 13786 26376
rect 15488 26373 15516 26404
rect 15473 26367 15531 26373
rect 13780 26336 13825 26364
rect 13780 26324 13786 26336
rect 15473 26333 15485 26367
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19705 26367 19763 26373
rect 19705 26364 19717 26367
rect 19392 26336 19717 26364
rect 19392 26324 19398 26336
rect 19705 26333 19717 26336
rect 19751 26333 19763 26367
rect 21100 26350 21128 26404
rect 23014 26392 23020 26404
rect 23072 26392 23078 26444
rect 24578 26432 24584 26444
rect 24539 26404 24584 26432
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 24857 26435 24915 26441
rect 24857 26401 24869 26435
rect 24903 26432 24915 26435
rect 25590 26432 25596 26444
rect 24903 26404 25596 26432
rect 24903 26401 24915 26404
rect 24857 26395 24915 26401
rect 25590 26392 25596 26404
rect 25648 26392 25654 26444
rect 29086 26392 29092 26444
rect 29144 26432 29150 26444
rect 30837 26435 30895 26441
rect 30837 26432 30849 26435
rect 29144 26404 30849 26432
rect 29144 26392 29150 26404
rect 30837 26401 30849 26404
rect 30883 26401 30895 26435
rect 30837 26395 30895 26401
rect 30926 26392 30932 26444
rect 30984 26432 30990 26444
rect 32309 26435 32367 26441
rect 32309 26432 32321 26435
rect 30984 26404 32321 26432
rect 30984 26392 30990 26404
rect 32309 26401 32321 26404
rect 32355 26401 32367 26435
rect 32309 26395 32367 26401
rect 19705 26327 19763 26333
rect 21266 26324 21272 26376
rect 21324 26364 21330 26376
rect 22005 26367 22063 26373
rect 22005 26364 22017 26367
rect 21324 26336 22017 26364
rect 21324 26324 21330 26336
rect 22005 26333 22017 26336
rect 22051 26333 22063 26367
rect 30558 26364 30564 26376
rect 30519 26336 30564 26364
rect 22005 26327 22063 26333
rect 30558 26324 30564 26336
rect 30616 26324 30622 26376
rect 34716 26364 34744 26472
rect 34790 26392 34796 26444
rect 34848 26432 34854 26444
rect 34885 26435 34943 26441
rect 34885 26432 34897 26435
rect 34848 26404 34897 26432
rect 34848 26392 34854 26404
rect 34885 26401 34897 26404
rect 34931 26401 34943 26435
rect 34992 26432 35020 26472
rect 37108 26472 38936 26500
rect 37108 26432 37136 26472
rect 38930 26460 38936 26472
rect 38988 26460 38994 26512
rect 34992 26404 37136 26432
rect 37185 26435 37243 26441
rect 34885 26395 34943 26401
rect 37185 26401 37197 26435
rect 37231 26432 37243 26435
rect 38470 26432 38476 26444
rect 37231 26404 38476 26432
rect 37231 26401 37243 26404
rect 37185 26395 37243 26401
rect 38470 26392 38476 26404
rect 38528 26392 38534 26444
rect 31970 26336 34744 26364
rect 13906 26256 13912 26308
rect 13964 26296 13970 26308
rect 14461 26299 14519 26305
rect 14461 26296 14473 26299
rect 13964 26268 14473 26296
rect 13964 26256 13970 26268
rect 14461 26265 14473 26268
rect 14507 26265 14519 26299
rect 14461 26259 14519 26265
rect 19981 26299 20039 26305
rect 19981 26265 19993 26299
rect 20027 26296 20039 26299
rect 20254 26296 20260 26308
rect 20027 26268 20260 26296
rect 20027 26265 20039 26268
rect 19981 26259 20039 26265
rect 20254 26256 20260 26268
rect 20312 26256 20318 26308
rect 26234 26296 26240 26308
rect 21376 26268 22324 26296
rect 26082 26268 26240 26296
rect 21376 26228 21404 26268
rect 13648 26200 21404 26228
rect 22097 26231 22155 26237
rect 22097 26197 22109 26231
rect 22143 26228 22155 26231
rect 22186 26228 22192 26240
rect 22143 26200 22192 26228
rect 22143 26197 22155 26200
rect 22097 26191 22155 26197
rect 22186 26188 22192 26200
rect 22244 26188 22250 26240
rect 22296 26228 22324 26268
rect 26234 26256 26240 26268
rect 26292 26256 26298 26308
rect 26418 26256 26424 26308
rect 26476 26296 26482 26308
rect 26605 26299 26663 26305
rect 26605 26296 26617 26299
rect 26476 26268 26617 26296
rect 26476 26256 26482 26268
rect 26605 26265 26617 26268
rect 26651 26265 26663 26299
rect 26605 26259 26663 26265
rect 30098 26256 30104 26308
rect 30156 26296 30162 26308
rect 30926 26296 30932 26308
rect 30156 26268 30932 26296
rect 30156 26256 30162 26268
rect 30926 26256 30932 26268
rect 30984 26256 30990 26308
rect 32122 26256 32128 26308
rect 32180 26296 32186 26308
rect 35161 26299 35219 26305
rect 35161 26296 35173 26299
rect 32180 26268 35173 26296
rect 32180 26256 32186 26268
rect 35161 26265 35173 26268
rect 35207 26265 35219 26299
rect 36538 26296 36544 26308
rect 36386 26268 36544 26296
rect 35161 26259 35219 26265
rect 36538 26256 36544 26268
rect 36596 26256 36602 26308
rect 37277 26299 37335 26305
rect 37277 26265 37289 26299
rect 37323 26265 37335 26299
rect 38194 26296 38200 26308
rect 38155 26268 38200 26296
rect 37277 26259 37335 26265
rect 26878 26228 26884 26240
rect 22296 26200 26884 26228
rect 26878 26188 26884 26200
rect 26936 26188 26942 26240
rect 36998 26188 37004 26240
rect 37056 26228 37062 26240
rect 37292 26228 37320 26259
rect 38194 26256 38200 26268
rect 38252 26256 38258 26308
rect 37056 26200 37320 26228
rect 37056 26188 37062 26200
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 8297 26027 8355 26033
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 9306 26024 9312 26036
rect 8343 25996 9312 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 12250 25984 12256 26036
rect 12308 26024 12314 26036
rect 14458 26024 14464 26036
rect 12308 25996 14464 26024
rect 12308 25984 12314 25996
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 21726 26024 21732 26036
rect 19996 25996 21732 26024
rect 10597 25959 10655 25965
rect 10597 25925 10609 25959
rect 10643 25956 10655 25959
rect 12066 25956 12072 25968
rect 10643 25928 12072 25956
rect 10643 25925 10655 25928
rect 10597 25919 10655 25925
rect 12066 25916 12072 25928
rect 12124 25916 12130 25968
rect 12713 25959 12771 25965
rect 12713 25925 12725 25959
rect 12759 25956 12771 25959
rect 14182 25956 14188 25968
rect 12759 25928 14188 25956
rect 12759 25925 12771 25928
rect 12713 25919 12771 25925
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 15654 25916 15660 25968
rect 15712 25956 15718 25968
rect 17405 25959 17463 25965
rect 17405 25956 17417 25959
rect 15712 25928 17417 25956
rect 15712 25916 15718 25928
rect 5169 25891 5227 25897
rect 5169 25857 5181 25891
rect 5215 25888 5227 25891
rect 5442 25888 5448 25900
rect 5215 25860 5448 25888
rect 5215 25857 5227 25860
rect 5169 25851 5227 25857
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 7742 25848 7748 25900
rect 7800 25888 7806 25900
rect 8481 25891 8539 25897
rect 8481 25888 8493 25891
rect 7800 25860 8493 25888
rect 7800 25848 7806 25860
rect 8481 25857 8493 25860
rect 8527 25857 8539 25891
rect 8481 25851 8539 25857
rect 11146 25848 11152 25900
rect 11204 25888 11210 25900
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 11204 25860 11897 25888
rect 11204 25848 11210 25860
rect 11885 25857 11897 25860
rect 11931 25888 11943 25891
rect 11974 25888 11980 25900
rect 11931 25860 11980 25888
rect 11931 25857 11943 25860
rect 11885 25851 11943 25857
rect 11974 25848 11980 25860
rect 12032 25848 12038 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 14921 25891 14979 25897
rect 14921 25888 14933 25891
rect 13872 25860 14933 25888
rect 13872 25848 13878 25860
rect 14921 25857 14933 25860
rect 14967 25888 14979 25891
rect 15102 25888 15108 25900
rect 14967 25860 15108 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 10502 25820 10508 25832
rect 10463 25792 10508 25820
rect 10502 25780 10508 25792
rect 10560 25780 10566 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 10612 25792 12633 25820
rect 8938 25712 8944 25764
rect 8996 25752 9002 25764
rect 10612 25752 10640 25792
rect 12621 25789 12633 25792
rect 12667 25789 12679 25823
rect 13262 25820 13268 25832
rect 13223 25792 13268 25820
rect 12621 25783 12679 25789
rect 13262 25780 13268 25792
rect 13320 25780 13326 25832
rect 11054 25752 11060 25764
rect 8996 25724 10640 25752
rect 10967 25724 11060 25752
rect 8996 25712 9002 25724
rect 11054 25712 11060 25724
rect 11112 25752 11118 25764
rect 12158 25752 12164 25764
rect 11112 25724 12164 25752
rect 11112 25712 11118 25724
rect 12158 25712 12164 25724
rect 12216 25712 12222 25764
rect 16758 25752 16764 25764
rect 14568 25724 16764 25752
rect 4982 25684 4988 25696
rect 4943 25656 4988 25684
rect 4982 25644 4988 25656
rect 5040 25644 5046 25696
rect 11977 25687 12035 25693
rect 11977 25653 11989 25687
rect 12023 25684 12035 25687
rect 14568 25684 14596 25724
rect 16758 25712 16764 25724
rect 16816 25712 16822 25764
rect 12023 25656 14596 25684
rect 12023 25653 12035 25656
rect 11977 25647 12035 25653
rect 14642 25644 14648 25696
rect 14700 25684 14706 25696
rect 15013 25687 15071 25693
rect 15013 25684 15025 25687
rect 14700 25656 15025 25684
rect 14700 25644 14706 25656
rect 15013 25653 15025 25656
rect 15059 25653 15071 25687
rect 16960 25684 16988 25928
rect 17405 25925 17417 25928
rect 17451 25925 17463 25959
rect 19996 25956 20024 25996
rect 21726 25984 21732 25996
rect 21784 25984 21790 26036
rect 33870 26024 33876 26036
rect 32600 25996 33876 26024
rect 21174 25956 21180 25968
rect 18630 25928 20024 25956
rect 20838 25928 21180 25956
rect 17405 25919 17463 25925
rect 21174 25916 21180 25928
rect 21232 25916 21238 25968
rect 30006 25916 30012 25968
rect 30064 25916 30070 25968
rect 32600 25965 32628 25996
rect 33870 25984 33876 25996
rect 33928 25984 33934 26036
rect 32585 25959 32643 25965
rect 32585 25925 32597 25959
rect 32631 25925 32643 25959
rect 32585 25919 32643 25925
rect 34698 25916 34704 25968
rect 34756 25956 34762 25968
rect 34977 25959 35035 25965
rect 34977 25956 34989 25959
rect 34756 25928 34989 25956
rect 34756 25916 34762 25928
rect 34977 25925 34989 25928
rect 35023 25925 35035 25959
rect 37090 25956 37096 25968
rect 36202 25928 37096 25956
rect 34977 25919 35035 25925
rect 37090 25916 37096 25928
rect 37148 25916 37154 25968
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25888 22063 25891
rect 22094 25888 22100 25900
rect 22051 25860 22100 25888
rect 22051 25857 22063 25860
rect 22005 25851 22063 25857
rect 22094 25848 22100 25860
rect 22152 25888 22158 25900
rect 24394 25888 24400 25900
rect 22152 25860 24400 25888
rect 22152 25848 22158 25860
rect 24394 25848 24400 25860
rect 24452 25848 24458 25900
rect 30558 25848 30564 25900
rect 30616 25888 30622 25900
rect 31662 25888 31668 25900
rect 30616 25860 31668 25888
rect 30616 25848 30622 25860
rect 31662 25848 31668 25860
rect 31720 25888 31726 25900
rect 32309 25891 32367 25897
rect 32309 25888 32321 25891
rect 31720 25860 32321 25888
rect 31720 25848 31726 25860
rect 32309 25857 32321 25860
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 33686 25848 33692 25900
rect 33744 25848 33750 25900
rect 38286 25888 38292 25900
rect 38247 25860 38292 25888
rect 38286 25848 38292 25860
rect 38344 25848 38350 25900
rect 17126 25820 17132 25832
rect 17087 25792 17132 25820
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 18877 25823 18935 25829
rect 18877 25789 18889 25823
rect 18923 25820 18935 25823
rect 19058 25820 19064 25832
rect 18923 25792 19064 25820
rect 18923 25789 18935 25792
rect 18877 25783 18935 25789
rect 19058 25780 19064 25792
rect 19116 25780 19122 25832
rect 19334 25820 19340 25832
rect 19295 25792 19340 25820
rect 19334 25780 19340 25792
rect 19392 25780 19398 25832
rect 19613 25823 19671 25829
rect 19613 25789 19625 25823
rect 19659 25820 19671 25823
rect 20162 25820 20168 25832
rect 19659 25792 20168 25820
rect 19659 25789 19671 25792
rect 19613 25783 19671 25789
rect 20162 25780 20168 25792
rect 20220 25820 20226 25832
rect 20220 25792 22232 25820
rect 20220 25780 20226 25792
rect 22204 25752 22232 25792
rect 22278 25780 22284 25832
rect 22336 25820 22342 25832
rect 22741 25823 22799 25829
rect 22741 25820 22753 25823
rect 22336 25792 22753 25820
rect 22336 25780 22342 25792
rect 22741 25789 22753 25792
rect 22787 25789 22799 25823
rect 22741 25783 22799 25789
rect 28721 25823 28779 25829
rect 28721 25789 28733 25823
rect 28767 25789 28779 25823
rect 28721 25783 28779 25789
rect 28997 25823 29055 25829
rect 28997 25789 29009 25823
rect 29043 25820 29055 25823
rect 29086 25820 29092 25832
rect 29043 25792 29092 25820
rect 29043 25789 29055 25792
rect 28997 25783 29055 25789
rect 24026 25752 24032 25764
rect 18432 25724 19012 25752
rect 22204 25724 24032 25752
rect 18432 25684 18460 25724
rect 16960 25656 18460 25684
rect 18984 25684 19012 25724
rect 24026 25712 24032 25724
rect 24084 25712 24090 25764
rect 21085 25687 21143 25693
rect 21085 25684 21097 25687
rect 18984 25656 21097 25684
rect 15013 25647 15071 25653
rect 21085 25653 21097 25656
rect 21131 25653 21143 25687
rect 28736 25684 28764 25783
rect 29086 25780 29092 25792
rect 29144 25780 29150 25832
rect 30742 25820 30748 25832
rect 30703 25792 30748 25820
rect 30742 25780 30748 25792
rect 30800 25780 30806 25832
rect 34701 25823 34759 25829
rect 34701 25820 34713 25823
rect 32324 25792 34713 25820
rect 32324 25696 32352 25792
rect 34701 25789 34713 25792
rect 34747 25789 34759 25823
rect 34701 25783 34759 25789
rect 34057 25755 34115 25761
rect 34057 25721 34069 25755
rect 34103 25752 34115 25755
rect 34606 25752 34612 25764
rect 34103 25724 34612 25752
rect 34103 25721 34115 25724
rect 34057 25715 34115 25721
rect 34606 25712 34612 25724
rect 34664 25712 34670 25764
rect 32306 25684 32312 25696
rect 28736 25656 32312 25684
rect 21085 25647 21143 25653
rect 32306 25644 32312 25656
rect 32364 25644 32370 25696
rect 33870 25644 33876 25696
rect 33928 25684 33934 25696
rect 36449 25687 36507 25693
rect 36449 25684 36461 25687
rect 33928 25656 36461 25684
rect 33928 25644 33934 25656
rect 36449 25653 36461 25656
rect 36495 25684 36507 25687
rect 36814 25684 36820 25696
rect 36495 25656 36820 25684
rect 36495 25653 36507 25656
rect 36449 25647 36507 25653
rect 36814 25644 36820 25656
rect 36872 25644 36878 25696
rect 38105 25687 38163 25693
rect 38105 25653 38117 25687
rect 38151 25684 38163 25687
rect 39298 25684 39304 25696
rect 38151 25656 39304 25684
rect 38151 25653 38163 25656
rect 38105 25647 38163 25653
rect 39298 25644 39304 25656
rect 39356 25644 39362 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 7742 25480 7748 25492
rect 7703 25452 7748 25480
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 9766 25480 9772 25492
rect 9727 25452 9772 25480
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 14366 25480 14372 25492
rect 14327 25452 14372 25480
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 15378 25440 15384 25492
rect 15436 25480 15442 25492
rect 16209 25483 16267 25489
rect 16209 25480 16221 25483
rect 15436 25452 16221 25480
rect 15436 25440 15442 25452
rect 16209 25449 16221 25452
rect 16255 25449 16267 25483
rect 16209 25443 16267 25449
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 20898 25480 20904 25492
rect 16816 25452 20904 25480
rect 16816 25440 16822 25452
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 24029 25483 24087 25489
rect 24029 25480 24041 25483
rect 22066 25452 24041 25480
rect 6917 25415 6975 25421
rect 6917 25381 6929 25415
rect 6963 25412 6975 25415
rect 8662 25412 8668 25424
rect 6963 25384 8668 25412
rect 6963 25381 6975 25384
rect 6917 25375 6975 25381
rect 8662 25372 8668 25384
rect 8720 25372 8726 25424
rect 10226 25412 10232 25424
rect 9508 25384 10232 25412
rect 8481 25347 8539 25353
rect 8481 25313 8493 25347
rect 8527 25344 8539 25347
rect 9309 25347 9367 25353
rect 9309 25344 9321 25347
rect 8527 25316 9321 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 9309 25313 9321 25316
rect 9355 25313 9367 25347
rect 9309 25307 9367 25313
rect 7098 25276 7104 25288
rect 7059 25248 7104 25276
rect 7098 25236 7104 25248
rect 7156 25236 7162 25288
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25276 7987 25279
rect 8389 25279 8447 25285
rect 8389 25276 8401 25279
rect 7975 25248 8401 25276
rect 7975 25245 7987 25248
rect 7929 25239 7987 25245
rect 8389 25245 8401 25248
rect 8435 25245 8447 25279
rect 8389 25239 8447 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9508 25276 9536 25384
rect 10226 25372 10232 25384
rect 10284 25372 10290 25424
rect 20714 25372 20720 25424
rect 20772 25412 20778 25424
rect 22066 25412 22094 25452
rect 24029 25449 24041 25452
rect 24075 25449 24087 25483
rect 36998 25480 37004 25492
rect 36959 25452 37004 25480
rect 24029 25443 24087 25449
rect 36998 25440 37004 25452
rect 37056 25440 37062 25492
rect 20772 25384 22094 25412
rect 20772 25372 20778 25384
rect 26878 25372 26884 25424
rect 26936 25412 26942 25424
rect 37645 25415 37703 25421
rect 37645 25412 37657 25415
rect 26936 25384 37657 25412
rect 26936 25372 26942 25384
rect 37645 25381 37657 25384
rect 37691 25381 37703 25415
rect 37645 25375 37703 25381
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 19429 25347 19487 25353
rect 19429 25344 19441 25347
rect 19392 25316 19441 25344
rect 19392 25304 19398 25316
rect 19429 25313 19441 25316
rect 19475 25344 19487 25347
rect 22278 25344 22284 25356
rect 19475 25316 22284 25344
rect 19475 25313 19487 25316
rect 19429 25307 19487 25313
rect 22278 25304 22284 25316
rect 22336 25304 22342 25356
rect 24581 25347 24639 25353
rect 24581 25313 24593 25347
rect 24627 25344 24639 25347
rect 25222 25344 25228 25356
rect 24627 25316 25228 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 25222 25304 25228 25316
rect 25280 25304 25286 25356
rect 14274 25276 14280 25288
rect 9171 25248 9536 25276
rect 14235 25248 14280 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 8404 25208 8432 25239
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 17862 25276 17868 25288
rect 16163 25248 17868 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 17862 25236 17868 25248
rect 17920 25236 17926 25288
rect 22186 25276 22192 25288
rect 20838 25248 22192 25276
rect 22186 25236 22192 25248
rect 22244 25236 22250 25288
rect 32306 25236 32312 25288
rect 32364 25276 32370 25288
rect 33597 25279 33655 25285
rect 33597 25276 33609 25279
rect 32364 25248 33609 25276
rect 32364 25236 32370 25248
rect 33597 25245 33609 25248
rect 33643 25245 33655 25279
rect 36906 25276 36912 25288
rect 36867 25248 36912 25276
rect 33597 25239 33655 25245
rect 36906 25236 36912 25248
rect 36964 25236 36970 25288
rect 37660 25276 37688 25375
rect 38013 25279 38071 25285
rect 38013 25276 38025 25279
rect 37660 25248 38025 25276
rect 38013 25245 38025 25248
rect 38059 25245 38071 25279
rect 38013 25239 38071 25245
rect 10410 25208 10416 25220
rect 8404 25180 10416 25208
rect 10410 25168 10416 25180
rect 10468 25168 10474 25220
rect 11606 25208 11612 25220
rect 11567 25180 11612 25208
rect 11606 25168 11612 25180
rect 11664 25168 11670 25220
rect 11698 25168 11704 25220
rect 11756 25208 11762 25220
rect 12250 25208 12256 25220
rect 11756 25180 11801 25208
rect 12211 25180 12256 25208
rect 11756 25168 11762 25180
rect 12250 25168 12256 25180
rect 12308 25168 12314 25220
rect 15013 25211 15071 25217
rect 15013 25177 15025 25211
rect 15059 25177 15071 25211
rect 15013 25171 15071 25177
rect 6638 25100 6644 25152
rect 6696 25140 6702 25152
rect 13630 25140 13636 25152
rect 6696 25112 13636 25140
rect 6696 25100 6702 25112
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 13722 25100 13728 25152
rect 13780 25140 13786 25152
rect 15028 25140 15056 25171
rect 15102 25168 15108 25220
rect 15160 25208 15166 25220
rect 15657 25211 15715 25217
rect 15160 25180 15205 25208
rect 15160 25168 15166 25180
rect 15657 25177 15669 25211
rect 15703 25208 15715 25211
rect 16390 25208 16396 25220
rect 15703 25180 16396 25208
rect 15703 25177 15715 25180
rect 15657 25171 15715 25177
rect 16390 25168 16396 25180
rect 16448 25168 16454 25220
rect 19702 25208 19708 25220
rect 19663 25180 19708 25208
rect 19702 25168 19708 25180
rect 19760 25168 19766 25220
rect 20990 25168 20996 25220
rect 21048 25208 21054 25220
rect 21450 25208 21456 25220
rect 21048 25180 21456 25208
rect 21048 25168 21054 25180
rect 21450 25168 21456 25180
rect 21508 25168 21514 25220
rect 21818 25168 21824 25220
rect 21876 25208 21882 25220
rect 22557 25211 22615 25217
rect 22557 25208 22569 25211
rect 21876 25180 22569 25208
rect 21876 25168 21882 25180
rect 22557 25177 22569 25180
rect 22603 25177 22615 25211
rect 24578 25208 24584 25220
rect 23782 25180 24584 25208
rect 22557 25171 22615 25177
rect 24578 25168 24584 25180
rect 24636 25168 24642 25220
rect 24857 25211 24915 25217
rect 24857 25177 24869 25211
rect 24903 25208 24915 25211
rect 24946 25208 24952 25220
rect 24903 25180 24952 25208
rect 24903 25177 24915 25180
rect 24857 25171 24915 25177
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 25866 25168 25872 25220
rect 25924 25168 25930 25220
rect 29730 25168 29736 25220
rect 29788 25208 29794 25220
rect 32861 25211 32919 25217
rect 32861 25208 32873 25211
rect 29788 25180 32873 25208
rect 29788 25168 29794 25180
rect 32861 25177 32873 25180
rect 32907 25177 32919 25211
rect 32861 25171 32919 25177
rect 16022 25140 16028 25152
rect 13780 25112 16028 25140
rect 13780 25100 13786 25112
rect 16022 25100 16028 25112
rect 16080 25100 16086 25152
rect 16482 25100 16488 25152
rect 16540 25140 16546 25152
rect 20530 25140 20536 25152
rect 16540 25112 20536 25140
rect 16540 25100 16546 25112
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 22186 25100 22192 25152
rect 22244 25140 22250 25152
rect 22646 25140 22652 25152
rect 22244 25112 22652 25140
rect 22244 25100 22250 25112
rect 22646 25100 22652 25112
rect 22704 25100 22710 25152
rect 24026 25100 24032 25152
rect 24084 25140 24090 25152
rect 26326 25140 26332 25152
rect 24084 25112 26332 25140
rect 24084 25100 24090 25112
rect 26326 25100 26332 25112
rect 26384 25100 26390 25152
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 10410 24896 10416 24948
rect 10468 24936 10474 24948
rect 22370 24936 22376 24948
rect 10468 24908 22376 24936
rect 10468 24896 10474 24908
rect 22370 24896 22376 24908
rect 22428 24936 22434 24948
rect 24581 24939 24639 24945
rect 24581 24936 24593 24939
rect 22428 24908 24593 24936
rect 22428 24896 22434 24908
rect 24581 24905 24593 24908
rect 24627 24905 24639 24939
rect 24581 24899 24639 24905
rect 10505 24871 10563 24877
rect 10505 24837 10517 24871
rect 10551 24868 10563 24871
rect 12342 24868 12348 24880
rect 10551 24840 11100 24868
rect 12303 24840 12348 24868
rect 10551 24837 10563 24840
rect 10505 24831 10563 24837
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 4982 24800 4988 24812
rect 1627 24772 4988 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 4982 24760 4988 24772
rect 5040 24760 5046 24812
rect 7837 24803 7895 24809
rect 7837 24769 7849 24803
rect 7883 24800 7895 24803
rect 8386 24800 8392 24812
rect 7883 24772 8392 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 8662 24800 8668 24812
rect 8623 24772 8668 24800
rect 8662 24760 8668 24772
rect 8720 24760 8726 24812
rect 10410 24732 10416 24744
rect 10371 24704 10416 24732
rect 10410 24692 10416 24704
rect 10468 24692 10474 24744
rect 10962 24664 10968 24676
rect 10923 24636 10968 24664
rect 10962 24624 10968 24636
rect 11020 24624 11026 24676
rect 11072 24664 11100 24840
rect 12342 24828 12348 24840
rect 12400 24828 12406 24880
rect 14642 24868 14648 24880
rect 14603 24840 14648 24868
rect 14642 24828 14648 24840
rect 14700 24828 14706 24880
rect 16482 24868 16488 24880
rect 15672 24840 16488 24868
rect 13814 24800 13820 24812
rect 13775 24772 13820 24800
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 15672 24809 15700 24840
rect 16482 24828 16488 24840
rect 16540 24828 16546 24880
rect 19334 24868 19340 24880
rect 19168 24840 19340 24868
rect 15657 24803 15715 24809
rect 13964 24772 14009 24800
rect 13964 24760 13970 24772
rect 15657 24769 15669 24803
rect 15703 24769 15715 24803
rect 15657 24763 15715 24769
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24800 15807 24803
rect 15930 24800 15936 24812
rect 15795 24772 15936 24800
rect 15795 24769 15807 24772
rect 15749 24763 15807 24769
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 19168 24809 19196 24840
rect 19334 24828 19340 24840
rect 19392 24868 19398 24880
rect 19702 24868 19708 24880
rect 19392 24840 19708 24868
rect 19392 24828 19398 24840
rect 19702 24828 19708 24840
rect 19760 24828 19766 24880
rect 23109 24871 23167 24877
rect 23109 24868 23121 24871
rect 22848 24840 23121 24868
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 17184 24772 19165 24800
rect 17184 24760 17190 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 22278 24800 22284 24812
rect 20562 24772 22284 24800
rect 19153 24763 19211 24769
rect 22278 24760 22284 24772
rect 22336 24760 22342 24812
rect 22848 24800 22876 24840
rect 23109 24837 23121 24840
rect 23155 24837 23167 24871
rect 23109 24831 23167 24837
rect 23198 24828 23204 24880
rect 23256 24868 23262 24880
rect 23256 24840 23598 24868
rect 23256 24828 23262 24840
rect 24394 24828 24400 24880
rect 24452 24868 24458 24880
rect 25041 24871 25099 24877
rect 25041 24868 25053 24871
rect 24452 24840 25053 24868
rect 24452 24828 24458 24840
rect 25041 24837 25053 24840
rect 25087 24837 25099 24871
rect 25041 24831 25099 24837
rect 28810 24800 28816 24812
rect 22572 24772 22876 24800
rect 28566 24772 28816 24800
rect 11882 24692 11888 24744
rect 11940 24732 11946 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 11940 24704 12265 24732
rect 11940 24692 11946 24704
rect 12253 24701 12265 24704
rect 12299 24732 12311 24735
rect 12342 24732 12348 24744
rect 12299 24704 12348 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12802 24732 12808 24744
rect 12763 24704 12808 24732
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 14826 24732 14832 24744
rect 14599 24704 14832 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 19429 24735 19487 24741
rect 19429 24701 19441 24735
rect 19475 24732 19487 24735
rect 19978 24732 19984 24744
rect 19475 24704 19984 24732
rect 19475 24701 19487 24704
rect 19429 24695 19487 24701
rect 19978 24692 19984 24704
rect 20036 24692 20042 24744
rect 12710 24664 12716 24676
rect 11072 24636 12716 24664
rect 12710 24624 12716 24636
rect 12768 24624 12774 24676
rect 15105 24667 15163 24673
rect 15105 24633 15117 24667
rect 15151 24664 15163 24667
rect 16574 24664 16580 24676
rect 15151 24636 16580 24664
rect 15151 24633 15163 24636
rect 15105 24627 15163 24633
rect 16574 24624 16580 24636
rect 16632 24624 16638 24676
rect 20806 24624 20812 24676
rect 20864 24664 20870 24676
rect 22572 24664 22600 24772
rect 28810 24760 28816 24772
rect 28868 24760 28874 24812
rect 30834 24760 30840 24812
rect 30892 24760 30898 24812
rect 32306 24800 32312 24812
rect 32267 24772 32312 24800
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 38286 24800 38292 24812
rect 33718 24772 38292 24800
rect 38286 24760 38292 24772
rect 38344 24760 38350 24812
rect 22833 24735 22891 24741
rect 22833 24701 22845 24735
rect 22879 24732 22891 24735
rect 23474 24732 23480 24744
rect 22879 24704 23480 24732
rect 22879 24701 22891 24704
rect 22833 24695 22891 24701
rect 23474 24692 23480 24704
rect 23532 24692 23538 24744
rect 25222 24692 25228 24744
rect 25280 24732 25286 24744
rect 25777 24735 25835 24741
rect 25777 24732 25789 24735
rect 25280 24704 25789 24732
rect 25280 24692 25286 24704
rect 25777 24701 25789 24704
rect 25823 24701 25835 24735
rect 27154 24732 27160 24744
rect 27115 24704 27160 24732
rect 25777 24695 25835 24701
rect 27154 24692 27160 24704
rect 27212 24692 27218 24744
rect 27430 24732 27436 24744
rect 27391 24704 27436 24732
rect 27430 24692 27436 24704
rect 27488 24692 27494 24744
rect 29454 24732 29460 24744
rect 28460 24704 29460 24732
rect 20864 24636 22600 24664
rect 20864 24624 20870 24636
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 7929 24599 7987 24605
rect 7929 24596 7941 24599
rect 7340 24568 7941 24596
rect 7340 24556 7346 24568
rect 7929 24565 7941 24568
rect 7975 24565 7987 24599
rect 7929 24559 7987 24565
rect 8481 24599 8539 24605
rect 8481 24565 8493 24599
rect 8527 24596 8539 24599
rect 9306 24596 9312 24608
rect 8527 24568 9312 24596
rect 8527 24565 8539 24568
rect 8481 24559 8539 24565
rect 9306 24556 9312 24568
rect 9364 24556 9370 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20901 24599 20959 24605
rect 20901 24596 20913 24599
rect 19484 24568 20913 24596
rect 19484 24556 19490 24568
rect 20901 24565 20913 24568
rect 20947 24565 20959 24599
rect 20901 24559 20959 24565
rect 22094 24556 22100 24608
rect 22152 24596 22158 24608
rect 26694 24596 26700 24608
rect 22152 24568 26700 24596
rect 22152 24556 22158 24568
rect 26694 24556 26700 24568
rect 26752 24556 26758 24608
rect 27154 24556 27160 24608
rect 27212 24596 27218 24608
rect 28460 24596 28488 24704
rect 29454 24692 29460 24704
rect 29512 24692 29518 24744
rect 29733 24735 29791 24741
rect 29733 24732 29745 24735
rect 29564 24704 29745 24732
rect 28534 24624 28540 24676
rect 28592 24624 28598 24676
rect 28718 24624 28724 24676
rect 28776 24664 28782 24676
rect 29564 24664 29592 24704
rect 29733 24701 29745 24704
rect 29779 24701 29791 24735
rect 29733 24695 29791 24701
rect 30190 24692 30196 24744
rect 30248 24732 30254 24744
rect 32585 24735 32643 24741
rect 30248 24704 31754 24732
rect 30248 24692 30254 24704
rect 28776 24636 29592 24664
rect 28776 24624 28782 24636
rect 27212 24568 28488 24596
rect 28552 24596 28580 24624
rect 28905 24599 28963 24605
rect 28905 24596 28917 24599
rect 28552 24568 28917 24596
rect 27212 24556 27218 24568
rect 28905 24565 28917 24568
rect 28951 24565 28963 24599
rect 28905 24559 28963 24565
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 31205 24599 31263 24605
rect 31205 24596 31217 24599
rect 29052 24568 31217 24596
rect 29052 24556 29058 24568
rect 31205 24565 31217 24568
rect 31251 24565 31263 24599
rect 31726 24596 31754 24704
rect 32585 24701 32597 24735
rect 32631 24732 32643 24735
rect 33870 24732 33876 24744
rect 32631 24704 33876 24732
rect 32631 24701 32643 24704
rect 32585 24695 32643 24701
rect 33870 24692 33876 24704
rect 33928 24692 33934 24744
rect 34054 24732 34060 24744
rect 34015 24704 34060 24732
rect 34054 24692 34060 24704
rect 34112 24692 34118 24744
rect 36446 24596 36452 24608
rect 31726 24568 36452 24596
rect 31205 24559 31263 24565
rect 36446 24556 36452 24568
rect 36504 24556 36510 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 8386 24352 8392 24404
rect 8444 24392 8450 24404
rect 9677 24395 9735 24401
rect 9677 24392 9689 24395
rect 8444 24364 9689 24392
rect 8444 24352 8450 24364
rect 9677 24361 9689 24364
rect 9723 24361 9735 24395
rect 9677 24355 9735 24361
rect 11149 24395 11207 24401
rect 11149 24361 11161 24395
rect 11195 24392 11207 24395
rect 11606 24392 11612 24404
rect 11195 24364 11612 24392
rect 11195 24361 11207 24364
rect 11149 24355 11207 24361
rect 11606 24352 11612 24364
rect 11664 24352 11670 24404
rect 11698 24352 11704 24404
rect 11756 24392 11762 24404
rect 11793 24395 11851 24401
rect 11793 24392 11805 24395
rect 11756 24364 11805 24392
rect 11756 24352 11762 24364
rect 11793 24361 11805 24364
rect 11839 24361 11851 24395
rect 22094 24392 22100 24404
rect 11793 24355 11851 24361
rect 13924 24364 22100 24392
rect 7837 24327 7895 24333
rect 7837 24293 7849 24327
rect 7883 24324 7895 24327
rect 13722 24324 13728 24336
rect 7883 24296 13728 24324
rect 7883 24293 7895 24296
rect 7837 24287 7895 24293
rect 13722 24284 13728 24296
rect 13780 24284 13786 24336
rect 9306 24256 9312 24268
rect 9267 24228 9312 24256
rect 9306 24216 9312 24228
rect 9364 24216 9370 24268
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 12621 24259 12679 24265
rect 12621 24256 12633 24259
rect 11388 24228 12633 24256
rect 11388 24216 11394 24228
rect 12621 24225 12633 24228
rect 12667 24225 12679 24259
rect 12621 24219 12679 24225
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 7282 24188 7288 24200
rect 1627 24160 2774 24188
rect 7243 24160 7288 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 2746 24052 2774 24160
rect 7282 24148 7288 24160
rect 7340 24148 7346 24200
rect 7742 24188 7748 24200
rect 7703 24160 7748 24188
rect 7742 24148 7748 24160
rect 7800 24148 7806 24200
rect 9122 24188 9128 24200
rect 9083 24160 9128 24188
rect 9122 24148 9128 24160
rect 9180 24148 9186 24200
rect 11054 24188 11060 24200
rect 11015 24160 11060 24188
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 11698 24188 11704 24200
rect 11659 24160 11704 24188
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 13357 24191 13415 24197
rect 12483 24160 13308 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 11716 24120 11744 24148
rect 13170 24120 13176 24132
rect 11716 24092 13176 24120
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 13280 24120 13308 24160
rect 13357 24157 13369 24191
rect 13403 24188 13415 24191
rect 13924 24188 13952 24364
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 22278 24352 22284 24404
rect 22336 24392 22342 24404
rect 24394 24392 24400 24404
rect 22336 24364 24400 24392
rect 22336 24352 22342 24364
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 31941 24395 31999 24401
rect 31941 24361 31953 24395
rect 31987 24392 31999 24395
rect 32122 24392 32128 24404
rect 31987 24364 32128 24392
rect 31987 24361 31999 24364
rect 31941 24355 31999 24361
rect 32122 24352 32128 24364
rect 32180 24392 32186 24404
rect 32398 24392 32404 24404
rect 32180 24364 32404 24392
rect 32180 24352 32186 24364
rect 32398 24352 32404 24364
rect 32456 24352 32462 24404
rect 34146 24392 34152 24404
rect 34107 24364 34152 24392
rect 34146 24352 34152 24364
rect 34204 24352 34210 24404
rect 14182 24284 14188 24336
rect 14240 24324 14246 24336
rect 14369 24327 14427 24333
rect 14369 24324 14381 24327
rect 14240 24296 14381 24324
rect 14240 24284 14246 24296
rect 14369 24293 14381 24296
rect 14415 24293 14427 24327
rect 14369 24287 14427 24293
rect 19058 24284 19064 24336
rect 19116 24324 19122 24336
rect 19116 24296 20208 24324
rect 19116 24284 19122 24296
rect 16298 24216 16304 24268
rect 16356 24256 16362 24268
rect 19610 24256 19616 24268
rect 16356 24228 19616 24256
rect 16356 24216 16362 24228
rect 19610 24216 19616 24228
rect 19668 24216 19674 24268
rect 19702 24216 19708 24268
rect 19760 24256 19766 24268
rect 20073 24259 20131 24265
rect 20073 24256 20085 24259
rect 19760 24228 20085 24256
rect 19760 24216 19766 24228
rect 20073 24225 20085 24228
rect 20119 24225 20131 24259
rect 20180 24256 20208 24296
rect 31726 24296 32536 24324
rect 20806 24256 20812 24268
rect 20180 24228 20812 24256
rect 20073 24219 20131 24225
rect 20806 24216 20812 24228
rect 20864 24216 20870 24268
rect 24854 24216 24860 24268
rect 24912 24256 24918 24268
rect 24949 24259 25007 24265
rect 24949 24256 24961 24259
rect 24912 24228 24961 24256
rect 24912 24216 24918 24228
rect 24949 24225 24961 24228
rect 24995 24225 25007 24259
rect 24949 24219 25007 24225
rect 30469 24259 30527 24265
rect 30469 24225 30481 24259
rect 30515 24256 30527 24259
rect 31726 24256 31754 24296
rect 30515 24228 31754 24256
rect 30515 24225 30527 24228
rect 30469 24219 30527 24225
rect 32306 24216 32312 24268
rect 32364 24256 32370 24268
rect 32401 24259 32459 24265
rect 32401 24256 32413 24259
rect 32364 24228 32413 24256
rect 32364 24216 32370 24228
rect 32401 24225 32413 24228
rect 32447 24225 32459 24259
rect 32508 24256 32536 24296
rect 34238 24256 34244 24268
rect 32508 24228 34244 24256
rect 32401 24219 32459 24225
rect 34238 24216 34244 24228
rect 34296 24216 34302 24268
rect 35161 24259 35219 24265
rect 35161 24225 35173 24259
rect 35207 24256 35219 24259
rect 36170 24256 36176 24268
rect 35207 24228 36176 24256
rect 35207 24225 35219 24228
rect 35161 24219 35219 24225
rect 36170 24216 36176 24228
rect 36228 24216 36234 24268
rect 13403 24160 13952 24188
rect 13403 24157 13415 24160
rect 13357 24151 13415 24157
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14182 24188 14188 24200
rect 14056 24160 14188 24188
rect 14056 24148 14062 24160
rect 14182 24148 14188 24160
rect 14240 24148 14246 24200
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 14323 24160 19564 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 19242 24120 19248 24132
rect 13280 24092 19248 24120
rect 19242 24080 19248 24092
rect 19300 24080 19306 24132
rect 7101 24055 7159 24061
rect 7101 24052 7113 24055
rect 2746 24024 7113 24052
rect 7101 24021 7113 24024
rect 7147 24021 7159 24055
rect 7101 24015 7159 24021
rect 13449 24055 13507 24061
rect 13449 24021 13461 24055
rect 13495 24052 13507 24055
rect 13998 24052 14004 24064
rect 13495 24024 14004 24052
rect 13495 24021 13507 24024
rect 13449 24015 13507 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 16482 24012 16488 24064
rect 16540 24052 16546 24064
rect 19426 24052 19432 24064
rect 16540 24024 19432 24052
rect 16540 24012 16546 24024
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 19536 24052 19564 24160
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 30193 24191 30251 24197
rect 30193 24188 30205 24191
rect 29512 24160 30205 24188
rect 29512 24148 29518 24160
rect 30193 24157 30205 24160
rect 30239 24157 30251 24191
rect 30193 24151 30251 24157
rect 31570 24148 31576 24200
rect 31628 24148 31634 24200
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 37458 24188 37464 24200
rect 37419 24160 37464 24188
rect 34885 24151 34943 24157
rect 37458 24148 37464 24160
rect 37516 24148 37522 24200
rect 37737 24191 37795 24197
rect 37737 24157 37749 24191
rect 37783 24188 37795 24191
rect 38102 24188 38108 24200
rect 37783 24160 38108 24188
rect 37783 24157 37795 24160
rect 37737 24151 37795 24157
rect 38102 24148 38108 24160
rect 38160 24148 38166 24200
rect 20346 24120 20352 24132
rect 20307 24092 20352 24120
rect 20346 24080 20352 24092
rect 20404 24080 20410 24132
rect 23290 24120 23296 24132
rect 21574 24092 23296 24120
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 24670 24120 24676 24132
rect 24631 24092 24676 24120
rect 24670 24080 24676 24092
rect 24728 24080 24734 24132
rect 24765 24123 24823 24129
rect 24765 24089 24777 24123
rect 24811 24089 24823 24123
rect 32677 24123 32735 24129
rect 32677 24120 32689 24123
rect 24765 24083 24823 24089
rect 31864 24092 32689 24120
rect 20990 24052 20996 24064
rect 19536 24024 20996 24052
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 21818 24052 21824 24064
rect 21140 24024 21824 24052
rect 21140 24012 21146 24024
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 21910 24012 21916 24064
rect 21968 24052 21974 24064
rect 24780 24052 24808 24083
rect 21968 24024 24808 24052
rect 21968 24012 21974 24024
rect 31110 24012 31116 24064
rect 31168 24052 31174 24064
rect 31864 24052 31892 24092
rect 32677 24089 32689 24092
rect 32723 24089 32735 24123
rect 34422 24120 34428 24132
rect 33902 24092 34428 24120
rect 32677 24083 32735 24089
rect 34422 24080 34428 24092
rect 34480 24080 34486 24132
rect 39482 24120 39488 24132
rect 36386 24092 39488 24120
rect 39482 24080 39488 24092
rect 39540 24080 39546 24132
rect 31168 24024 31892 24052
rect 31168 24012 31174 24024
rect 35434 24012 35440 24064
rect 35492 24052 35498 24064
rect 36633 24055 36691 24061
rect 36633 24052 36645 24055
rect 35492 24024 36645 24052
rect 35492 24012 35498 24024
rect 36633 24021 36645 24024
rect 36679 24021 36691 24055
rect 36633 24015 36691 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 13372 23820 19196 23848
rect 11885 23783 11943 23789
rect 11885 23749 11897 23783
rect 11931 23780 11943 23783
rect 12434 23780 12440 23792
rect 11931 23752 12440 23780
rect 11931 23749 11943 23752
rect 11885 23743 11943 23749
rect 12434 23740 12440 23752
rect 12492 23740 12498 23792
rect 13372 23721 13400 23820
rect 13357 23715 13415 23721
rect 13357 23681 13369 23715
rect 13403 23681 13415 23715
rect 17034 23712 17040 23724
rect 16995 23684 17040 23712
rect 13357 23675 13415 23681
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 10965 23647 11023 23653
rect 10965 23613 10977 23647
rect 11011 23644 11023 23647
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11011 23616 11805 23644
rect 11011 23613 11023 23616
rect 10965 23607 11023 23613
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 12250 23644 12256 23656
rect 12211 23616 12256 23644
rect 11793 23607 11851 23613
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 17313 23647 17371 23653
rect 17313 23613 17325 23647
rect 17359 23644 17371 23647
rect 17954 23644 17960 23656
rect 17359 23616 17960 23644
rect 17359 23613 17371 23616
rect 17313 23607 17371 23613
rect 17954 23604 17960 23616
rect 18012 23604 18018 23656
rect 13170 23536 13176 23588
rect 13228 23576 13234 23588
rect 18432 23576 18460 23698
rect 19168 23644 19196 23820
rect 19334 23808 19340 23860
rect 19392 23808 19398 23860
rect 23382 23808 23388 23860
rect 23440 23848 23446 23860
rect 25222 23848 25228 23860
rect 23440 23820 25228 23848
rect 23440 23808 23446 23820
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 26970 23808 26976 23860
rect 27028 23848 27034 23860
rect 29365 23851 29423 23857
rect 29365 23848 29377 23851
rect 27028 23820 29377 23848
rect 27028 23808 27034 23820
rect 29365 23817 29377 23820
rect 29411 23817 29423 23851
rect 36906 23848 36912 23860
rect 29365 23811 29423 23817
rect 31726 23820 36912 23848
rect 19352 23780 19380 23808
rect 19260 23752 19380 23780
rect 19260 23721 19288 23752
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19521 23783 19579 23789
rect 19521 23780 19533 23783
rect 19484 23752 19533 23780
rect 19484 23740 19490 23752
rect 19521 23749 19533 23752
rect 19567 23749 19579 23783
rect 19521 23743 19579 23749
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21269 23783 21327 23789
rect 21269 23780 21281 23783
rect 21048 23752 21281 23780
rect 21048 23740 21054 23752
rect 21269 23749 21281 23752
rect 21315 23780 21327 23783
rect 23661 23783 23719 23789
rect 23661 23780 23673 23783
rect 21315 23752 23673 23780
rect 21315 23749 21327 23752
rect 21269 23743 21327 23749
rect 23661 23749 23673 23752
rect 23707 23749 23719 23783
rect 28166 23780 28172 23792
rect 24886 23752 28172 23780
rect 23661 23743 23719 23749
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 30374 23780 30380 23792
rect 29118 23752 30380 23780
rect 30374 23740 30380 23752
rect 30432 23740 30438 23792
rect 31726 23780 31754 23820
rect 36906 23808 36912 23820
rect 36964 23808 36970 23860
rect 37550 23848 37556 23860
rect 37511 23820 37556 23848
rect 37550 23808 37556 23820
rect 37608 23808 37614 23860
rect 34790 23780 34796 23792
rect 31326 23752 31754 23780
rect 34440 23752 34796 23780
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 22462 23712 22468 23724
rect 20654 23684 22468 23712
rect 19245 23675 19303 23681
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 23382 23712 23388 23724
rect 23343 23684 23388 23712
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 27154 23672 27160 23724
rect 27212 23712 27218 23724
rect 27617 23715 27675 23721
rect 27617 23712 27629 23715
rect 27212 23684 27629 23712
rect 27212 23672 27218 23684
rect 27617 23681 27629 23684
rect 27663 23681 27675 23715
rect 27617 23675 27675 23681
rect 29454 23672 29460 23724
rect 29512 23712 29518 23724
rect 29825 23715 29883 23721
rect 29825 23712 29837 23715
rect 29512 23684 29837 23712
rect 29512 23672 29518 23684
rect 29825 23681 29837 23684
rect 29871 23681 29883 23715
rect 29825 23675 29883 23681
rect 32306 23672 32312 23724
rect 32364 23712 32370 23724
rect 34440 23721 34468 23752
rect 34790 23740 34796 23752
rect 34848 23740 34854 23792
rect 37642 23780 37648 23792
rect 35926 23752 37648 23780
rect 37642 23740 37648 23752
rect 37700 23740 37706 23792
rect 34425 23715 34483 23721
rect 34425 23712 34437 23715
rect 32364 23684 34437 23712
rect 32364 23672 32370 23684
rect 34425 23681 34437 23684
rect 34471 23681 34483 23715
rect 36446 23712 36452 23724
rect 36407 23684 36452 23712
rect 34425 23675 34483 23681
rect 36446 23672 36452 23684
rect 36504 23672 36510 23724
rect 37461 23715 37519 23721
rect 37461 23681 37473 23715
rect 37507 23712 37519 23715
rect 39758 23712 39764 23724
rect 37507 23684 39764 23712
rect 37507 23681 37519 23684
rect 37461 23675 37519 23681
rect 39758 23672 39764 23684
rect 39816 23672 39822 23724
rect 19168 23616 21588 23644
rect 21560 23576 21588 23616
rect 21634 23604 21640 23656
rect 21692 23644 21698 23656
rect 21818 23644 21824 23656
rect 21692 23616 21824 23644
rect 21692 23604 21698 23616
rect 21818 23604 21824 23616
rect 21876 23604 21882 23656
rect 25130 23644 25136 23656
rect 23485 23616 25136 23644
rect 23485 23576 23513 23616
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25409 23647 25467 23653
rect 25409 23613 25421 23647
rect 25455 23644 25467 23647
rect 26326 23644 26332 23656
rect 25455 23616 26332 23644
rect 25455 23613 25467 23616
rect 25409 23607 25467 23613
rect 26326 23604 26332 23616
rect 26384 23604 26390 23656
rect 27893 23647 27951 23653
rect 27893 23613 27905 23647
rect 27939 23644 27951 23647
rect 28258 23644 28264 23656
rect 27939 23616 28264 23644
rect 27939 23613 27951 23616
rect 27893 23607 27951 23613
rect 28258 23604 28264 23616
rect 28316 23644 28322 23656
rect 28902 23644 28908 23656
rect 28316 23616 28908 23644
rect 28316 23604 28322 23616
rect 28902 23604 28908 23616
rect 28960 23604 28966 23656
rect 30098 23644 30104 23656
rect 30059 23616 30104 23644
rect 30098 23604 30104 23616
rect 30156 23604 30162 23656
rect 34330 23604 34336 23656
rect 34388 23644 34394 23656
rect 34701 23647 34759 23653
rect 34701 23644 34713 23647
rect 34388 23616 34713 23644
rect 34388 23604 34394 23616
rect 34701 23613 34713 23616
rect 34747 23613 34759 23647
rect 34701 23607 34759 23613
rect 13228 23548 17172 23576
rect 18432 23548 19334 23576
rect 21560 23548 23513 23576
rect 13228 23536 13234 23548
rect 12710 23468 12716 23520
rect 12768 23508 12774 23520
rect 13449 23511 13507 23517
rect 13449 23508 13461 23511
rect 12768 23480 13461 23508
rect 12768 23468 12774 23480
rect 13449 23477 13461 23480
rect 13495 23477 13507 23511
rect 17144 23508 17172 23548
rect 18598 23508 18604 23520
rect 17144 23480 18604 23508
rect 13449 23471 13507 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 18782 23508 18788 23520
rect 18743 23480 18788 23508
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 19306 23508 19334 23548
rect 25590 23536 25596 23588
rect 25648 23576 25654 23588
rect 27614 23576 27620 23588
rect 25648 23548 27620 23576
rect 25648 23536 25654 23548
rect 27614 23536 27620 23548
rect 27672 23536 27678 23588
rect 29270 23536 29276 23588
rect 29328 23576 29334 23588
rect 29328 23548 29960 23576
rect 29328 23536 29334 23548
rect 21450 23508 21456 23520
rect 19306 23480 21456 23508
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 23750 23468 23756 23520
rect 23808 23508 23814 23520
rect 28534 23508 28540 23520
rect 23808 23480 28540 23508
rect 23808 23468 23814 23480
rect 28534 23468 28540 23480
rect 28592 23468 28598 23520
rect 29932 23508 29960 23548
rect 31386 23508 31392 23520
rect 29932 23480 31392 23508
rect 31386 23468 31392 23480
rect 31444 23508 31450 23520
rect 31573 23511 31631 23517
rect 31573 23508 31585 23511
rect 31444 23480 31585 23508
rect 31444 23468 31450 23480
rect 31573 23477 31585 23480
rect 31619 23477 31631 23511
rect 31573 23471 31631 23477
rect 32950 23468 32956 23520
rect 33008 23508 33014 23520
rect 34514 23508 34520 23520
rect 33008 23480 34520 23508
rect 33008 23468 33014 23480
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 9122 23264 9128 23316
rect 9180 23304 9186 23316
rect 9493 23307 9551 23313
rect 9493 23304 9505 23307
rect 9180 23276 9505 23304
rect 9180 23264 9186 23276
rect 9493 23273 9505 23276
rect 9539 23273 9551 23307
rect 9493 23267 9551 23273
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12492 23276 12537 23304
rect 12492 23264 12498 23276
rect 15102 23264 15108 23316
rect 15160 23304 15166 23316
rect 15565 23307 15623 23313
rect 15565 23304 15577 23307
rect 15160 23276 15577 23304
rect 15160 23264 15166 23276
rect 15565 23273 15577 23276
rect 15611 23273 15623 23307
rect 15565 23267 15623 23273
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 20070 23304 20076 23316
rect 19484 23276 20076 23304
rect 19484 23264 19490 23276
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 20180 23276 21772 23304
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20180 23236 20208 23276
rect 19944 23208 20208 23236
rect 19944 23196 19950 23208
rect 14918 23168 14924 23180
rect 11532 23140 14924 23168
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8904 23072 9137 23100
rect 8904 23060 8910 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9306 23100 9312 23112
rect 9267 23072 9312 23100
rect 9125 23063 9183 23069
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 11532 23109 11560 23140
rect 14918 23128 14924 23140
rect 14976 23128 14982 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 20714 23168 20720 23180
rect 19392 23140 20392 23168
rect 20675 23140 20720 23168
rect 19392 23128 19398 23140
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23100 12403 23103
rect 12986 23100 12992 23112
rect 12391 23072 12992 23100
rect 12391 23069 12403 23072
rect 12345 23063 12403 23069
rect 12986 23060 12992 23072
rect 13044 23060 13050 23112
rect 15746 23100 15752 23112
rect 15707 23072 15752 23100
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 19886 23100 19892 23112
rect 17460 23072 19892 23100
rect 17460 23060 17466 23072
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 20364 23100 20392 23140
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 21744 23168 21772 23276
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 23750 23304 23756 23316
rect 22888 23276 23756 23304
rect 22888 23264 22894 23276
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 24210 23264 24216 23316
rect 24268 23304 24274 23316
rect 31110 23304 31116 23316
rect 24268 23276 31116 23304
rect 24268 23264 24274 23276
rect 31110 23264 31116 23276
rect 31168 23264 31174 23316
rect 31220 23276 33548 23304
rect 27614 23196 27620 23248
rect 27672 23236 27678 23248
rect 31220 23236 31248 23276
rect 27672 23208 31248 23236
rect 27672 23196 27678 23208
rect 23385 23171 23443 23177
rect 23385 23168 23397 23171
rect 21744 23140 23397 23168
rect 23385 23137 23397 23140
rect 23431 23137 23443 23171
rect 23385 23131 23443 23137
rect 24029 23171 24087 23177
rect 24029 23137 24041 23171
rect 24075 23168 24087 23171
rect 29362 23168 29368 23180
rect 24075 23140 29368 23168
rect 24075 23137 24087 23140
rect 24029 23131 24087 23137
rect 29362 23128 29368 23140
rect 29420 23128 29426 23180
rect 29454 23128 29460 23180
rect 29512 23168 29518 23180
rect 30469 23171 30527 23177
rect 30469 23168 30481 23171
rect 29512 23140 30481 23168
rect 29512 23128 29518 23140
rect 30469 23137 30481 23140
rect 30515 23137 30527 23171
rect 30469 23131 30527 23137
rect 31481 23171 31539 23177
rect 31481 23137 31493 23171
rect 31527 23168 31539 23171
rect 32306 23168 32312 23180
rect 31527 23140 32312 23168
rect 31527 23137 31539 23140
rect 31481 23131 31539 23137
rect 32306 23128 32312 23140
rect 32364 23128 32370 23180
rect 33520 23177 33548 23276
rect 33505 23171 33563 23177
rect 33505 23137 33517 23171
rect 33551 23137 33563 23171
rect 33505 23131 33563 23137
rect 34790 23128 34796 23180
rect 34848 23168 34854 23180
rect 34885 23171 34943 23177
rect 34885 23168 34897 23171
rect 34848 23140 34897 23168
rect 34848 23128 34854 23140
rect 34885 23137 34897 23140
rect 34931 23137 34943 23171
rect 34885 23131 34943 23137
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20364 23072 20453 23100
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 24762 23060 24768 23112
rect 24820 23100 24826 23112
rect 25222 23100 25228 23112
rect 24820 23072 25228 23100
rect 24820 23060 24826 23072
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 29730 23100 29736 23112
rect 29691 23072 29736 23100
rect 29730 23060 29736 23072
rect 29788 23060 29794 23112
rect 37458 23060 37464 23112
rect 37516 23100 37522 23112
rect 37553 23103 37611 23109
rect 37553 23100 37565 23103
rect 37516 23072 37565 23100
rect 37516 23060 37522 23072
rect 37553 23069 37565 23072
rect 37599 23069 37611 23103
rect 37553 23063 37611 23069
rect 19978 22992 19984 23044
rect 20036 23032 20042 23044
rect 20036 23004 20668 23032
rect 21942 23004 23428 23032
rect 20036 22992 20042 23004
rect 11609 22967 11667 22973
rect 11609 22933 11621 22967
rect 11655 22964 11667 22967
rect 11882 22964 11888 22976
rect 11655 22936 11888 22964
rect 11655 22933 11667 22936
rect 11609 22927 11667 22933
rect 11882 22924 11888 22936
rect 11940 22924 11946 22976
rect 17862 22924 17868 22976
rect 17920 22964 17926 22976
rect 20530 22964 20536 22976
rect 17920 22936 20536 22964
rect 17920 22924 17926 22936
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 20640 22964 20668 23004
rect 22189 22967 22247 22973
rect 22189 22964 22201 22967
rect 20640 22936 22201 22964
rect 22189 22933 22201 22936
rect 22235 22933 22247 22967
rect 23400 22964 23428 23004
rect 23474 22992 23480 23044
rect 23532 23032 23538 23044
rect 25498 23032 25504 23044
rect 23532 23004 23577 23032
rect 25459 23004 25504 23032
rect 23532 22992 23538 23004
rect 25498 22992 25504 23004
rect 25556 22992 25562 23044
rect 27522 23032 27528 23044
rect 26726 23004 27528 23032
rect 27522 22992 27528 23004
rect 27580 22992 27586 23044
rect 31757 23035 31815 23041
rect 31757 23001 31769 23035
rect 31803 23032 31815 23035
rect 31846 23032 31852 23044
rect 31803 23004 31852 23032
rect 31803 23001 31815 23004
rect 31757 22995 31815 23001
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 35066 23032 35072 23044
rect 32982 23004 35072 23032
rect 35066 22992 35072 23004
rect 35124 22992 35130 23044
rect 35161 23035 35219 23041
rect 35161 23001 35173 23035
rect 35207 23001 35219 23035
rect 36998 23032 37004 23044
rect 36386 23004 37004 23032
rect 35161 22995 35219 23001
rect 25038 22964 25044 22976
rect 23400 22936 25044 22964
rect 22189 22927 22247 22933
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 25516 22964 25544 22992
rect 26418 22964 26424 22976
rect 25516 22936 26424 22964
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 26786 22924 26792 22976
rect 26844 22964 26850 22976
rect 26973 22967 27031 22973
rect 26973 22964 26985 22967
rect 26844 22936 26985 22964
rect 26844 22924 26850 22936
rect 26973 22933 26985 22936
rect 27019 22933 27031 22967
rect 26973 22927 27031 22933
rect 32674 22924 32680 22976
rect 32732 22964 32738 22976
rect 35176 22964 35204 22995
rect 36998 22992 37004 23004
rect 37056 22992 37062 23044
rect 36630 22964 36636 22976
rect 32732 22936 35204 22964
rect 36591 22936 36636 22964
rect 32732 22924 32738 22936
rect 36630 22924 36636 22936
rect 36688 22924 36694 22976
rect 37274 22924 37280 22976
rect 37332 22964 37338 22976
rect 37645 22967 37703 22973
rect 37645 22964 37657 22967
rect 37332 22936 37657 22964
rect 37332 22924 37338 22936
rect 37645 22933 37657 22936
rect 37691 22933 37703 22967
rect 37645 22927 37703 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 14734 22760 14740 22772
rect 12452 22732 14740 22760
rect 12342 22692 12348 22704
rect 12303 22664 12348 22692
rect 12342 22652 12348 22664
rect 12400 22652 12406 22704
rect 12452 22701 12480 22732
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 20070 22760 20076 22772
rect 15068 22732 20076 22760
rect 15068 22720 15074 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 24118 22760 24124 22772
rect 20588 22732 24124 22760
rect 20588 22720 20594 22732
rect 24118 22720 24124 22732
rect 24176 22720 24182 22772
rect 25590 22720 25596 22772
rect 25648 22760 25654 22772
rect 25648 22732 25728 22760
rect 25648 22720 25654 22732
rect 12437 22695 12495 22701
rect 12437 22661 12449 22695
rect 12483 22661 12495 22695
rect 13998 22692 14004 22704
rect 13959 22664 14004 22692
rect 12437 22655 12495 22661
rect 13998 22652 14004 22664
rect 14056 22652 14062 22704
rect 18230 22652 18236 22704
rect 18288 22692 18294 22704
rect 18782 22692 18788 22704
rect 18288 22664 18788 22692
rect 18288 22652 18294 22664
rect 18782 22652 18788 22664
rect 18840 22652 18846 22704
rect 22002 22692 22008 22704
rect 20010 22664 22008 22692
rect 22002 22652 22008 22664
rect 22060 22652 22066 22704
rect 23937 22695 23995 22701
rect 23937 22692 23949 22695
rect 23032 22664 23949 22692
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 7340 22596 9137 22624
rect 7340 22584 7346 22596
rect 9125 22593 9137 22596
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 9272 22596 10241 22624
rect 9272 22584 9278 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22624 11023 22627
rect 11698 22624 11704 22636
rect 11011 22596 11704 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 15286 22584 15292 22636
rect 15344 22624 15350 22636
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 15344 22596 15853 22624
rect 15344 22584 15350 22596
rect 15841 22593 15853 22596
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 21358 22584 21364 22636
rect 21416 22624 21422 22636
rect 23032 22624 23060 22664
rect 23937 22661 23949 22664
rect 23983 22661 23995 22695
rect 23937 22655 23995 22661
rect 24489 22695 24547 22701
rect 24489 22661 24501 22695
rect 24535 22692 24547 22695
rect 24854 22692 24860 22704
rect 24535 22664 24860 22692
rect 24535 22661 24547 22664
rect 24489 22655 24547 22661
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 25700 22701 25728 22732
rect 26142 22720 26148 22772
rect 26200 22760 26206 22772
rect 26200 22732 27476 22760
rect 26200 22720 26206 22732
rect 27448 22701 27476 22732
rect 31110 22720 31116 22772
rect 31168 22760 31174 22772
rect 31665 22763 31723 22769
rect 31665 22760 31677 22763
rect 31168 22732 31677 22760
rect 31168 22720 31174 22732
rect 31665 22729 31677 22732
rect 31711 22729 31723 22763
rect 36078 22760 36084 22772
rect 31665 22723 31723 22729
rect 35452 22732 36084 22760
rect 25685 22695 25743 22701
rect 25685 22661 25697 22695
rect 25731 22661 25743 22695
rect 25685 22655 25743 22661
rect 27433 22695 27491 22701
rect 27433 22661 27445 22695
rect 27479 22661 27491 22695
rect 30466 22692 30472 22704
rect 28658 22664 30472 22692
rect 27433 22655 27491 22661
rect 30466 22652 30472 22664
rect 30524 22652 30530 22704
rect 31846 22692 31852 22704
rect 31418 22664 31852 22692
rect 31846 22652 31852 22664
rect 31904 22652 31910 22704
rect 35452 22692 35480 22732
rect 36078 22720 36084 22732
rect 36136 22720 36142 22772
rect 36446 22720 36452 22772
rect 36504 22760 36510 22772
rect 36541 22763 36599 22769
rect 36541 22760 36553 22763
rect 36504 22732 36553 22760
rect 36504 22720 36510 22732
rect 36541 22729 36553 22732
rect 36587 22729 36599 22763
rect 36541 22723 36599 22729
rect 37182 22692 37188 22704
rect 33810 22664 35480 22692
rect 36294 22664 37188 22692
rect 37182 22652 37188 22664
rect 37240 22652 37246 22704
rect 21416 22596 23060 22624
rect 25409 22627 25467 22633
rect 21416 22584 21422 22596
rect 25409 22593 25421 22627
rect 25455 22624 25467 22627
rect 25774 22624 25780 22636
rect 25455 22596 25780 22624
rect 25455 22593 25467 22596
rect 25409 22587 25467 22593
rect 25774 22584 25780 22596
rect 25832 22584 25838 22636
rect 26329 22627 26387 22633
rect 26329 22593 26341 22627
rect 26375 22593 26387 22627
rect 27154 22624 27160 22636
rect 27115 22596 27160 22624
rect 26329 22587 26387 22593
rect 8297 22559 8355 22565
rect 8297 22525 8309 22559
rect 8343 22556 8355 22559
rect 8941 22559 8999 22565
rect 8941 22556 8953 22559
rect 8343 22528 8953 22556
rect 8343 22525 8355 22528
rect 8297 22519 8355 22525
rect 8941 22525 8953 22528
rect 8987 22525 8999 22559
rect 11054 22556 11060 22568
rect 8941 22519 8999 22525
rect 9048 22528 11060 22556
rect 1857 22491 1915 22497
rect 1857 22457 1869 22491
rect 1903 22488 1915 22491
rect 9048 22488 9076 22528
rect 11054 22516 11060 22528
rect 11112 22556 11118 22568
rect 11606 22556 11612 22568
rect 11112 22528 11612 22556
rect 11112 22516 11118 22528
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 13354 22556 13360 22568
rect 13315 22528 13360 22556
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 13909 22559 13967 22565
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 14366 22556 14372 22568
rect 13955 22528 14372 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 14918 22556 14924 22568
rect 14879 22528 14924 22556
rect 14918 22516 14924 22528
rect 14976 22516 14982 22568
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22556 18567 22559
rect 19334 22556 19340 22568
rect 18555 22528 19340 22556
rect 18555 22525 18567 22528
rect 18509 22519 18567 22525
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23624 22528 23857 22556
rect 23624 22516 23630 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 26344 22556 26372 22587
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 29454 22584 29460 22636
rect 29512 22624 29518 22636
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29512 22596 29929 22624
rect 29512 22584 29518 22596
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 34238 22584 34244 22636
rect 34296 22624 34302 22636
rect 34333 22627 34391 22633
rect 34333 22624 34345 22627
rect 34296 22596 34345 22624
rect 34296 22584 34302 22596
rect 34333 22593 34345 22596
rect 34379 22593 34391 22627
rect 34790 22624 34796 22636
rect 34751 22596 34796 22624
rect 34333 22587 34391 22593
rect 34790 22584 34796 22596
rect 34848 22584 34854 22636
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 37608 22596 38025 22624
rect 37608 22584 37614 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 23845 22519 23903 22525
rect 25240 22528 26372 22556
rect 26421 22559 26479 22565
rect 1903 22460 9076 22488
rect 1903 22457 1915 22460
rect 1857 22451 1915 22457
rect 9122 22448 9128 22500
rect 9180 22488 9186 22500
rect 9309 22491 9367 22497
rect 9309 22488 9321 22491
rect 9180 22460 9321 22488
rect 9180 22448 9186 22460
rect 9309 22457 9321 22460
rect 9355 22457 9367 22491
rect 9309 22451 9367 22457
rect 10321 22491 10379 22497
rect 10321 22457 10333 22491
rect 10367 22488 10379 22491
rect 14826 22488 14832 22500
rect 10367 22460 14832 22488
rect 10367 22457 10379 22460
rect 10321 22451 10379 22457
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 20254 22488 20260 22500
rect 20215 22460 20260 22488
rect 20254 22448 20260 22460
rect 20312 22448 20318 22500
rect 21266 22448 21272 22500
rect 21324 22488 21330 22500
rect 25240 22488 25268 22528
rect 26421 22525 26433 22559
rect 26467 22556 26479 22559
rect 26602 22556 26608 22568
rect 26467 22528 26608 22556
rect 26467 22525 26479 22528
rect 26421 22519 26479 22525
rect 26602 22516 26608 22528
rect 26660 22516 26666 22568
rect 30190 22556 30196 22568
rect 29932 22528 30196 22556
rect 21324 22460 25268 22488
rect 28905 22491 28963 22497
rect 21324 22448 21330 22460
rect 28905 22457 28917 22491
rect 28951 22488 28963 22491
rect 29822 22488 29828 22500
rect 28951 22460 29828 22488
rect 28951 22457 28963 22460
rect 28905 22451 28963 22457
rect 29822 22448 29828 22460
rect 29880 22448 29886 22500
rect 11054 22420 11060 22432
rect 11015 22392 11060 22420
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 15933 22423 15991 22429
rect 15933 22389 15945 22423
rect 15979 22420 15991 22423
rect 17310 22420 17316 22432
rect 15979 22392 17316 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 18598 22380 18604 22432
rect 18656 22420 18662 22432
rect 20714 22420 20720 22432
rect 18656 22392 20720 22420
rect 18656 22380 18662 22392
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 24118 22380 24124 22432
rect 24176 22420 24182 22432
rect 29549 22423 29607 22429
rect 29549 22420 29561 22423
rect 24176 22392 29561 22420
rect 24176 22380 24182 22392
rect 29549 22389 29561 22392
rect 29595 22420 29607 22423
rect 29932 22420 29960 22528
rect 30190 22516 30196 22528
rect 30248 22516 30254 22568
rect 30558 22516 30564 22568
rect 30616 22556 30622 22568
rect 30616 22528 32260 22556
rect 30616 22516 30622 22528
rect 29595 22392 29960 22420
rect 32232 22420 32260 22528
rect 32306 22516 32312 22568
rect 32364 22556 32370 22568
rect 32585 22559 32643 22565
rect 32364 22528 32409 22556
rect 32364 22516 32370 22528
rect 32585 22525 32597 22559
rect 32631 22556 32643 22559
rect 32674 22556 32680 22568
rect 32631 22528 32680 22556
rect 32631 22525 32643 22528
rect 32585 22519 32643 22525
rect 32674 22516 32680 22528
rect 32732 22516 32738 22568
rect 35069 22559 35127 22565
rect 35069 22556 35081 22559
rect 33612 22528 35081 22556
rect 33612 22420 33640 22528
rect 35069 22525 35081 22528
rect 35115 22556 35127 22559
rect 35434 22556 35440 22568
rect 35115 22528 35440 22556
rect 35115 22525 35127 22528
rect 35069 22519 35127 22525
rect 35434 22516 35440 22528
rect 35492 22516 35498 22568
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 32232 22392 33640 22420
rect 29595 22389 29607 22392
rect 29549 22383 29607 22389
rect 34330 22380 34336 22432
rect 34388 22420 34394 22432
rect 35618 22420 35624 22432
rect 34388 22392 35624 22420
rect 34388 22380 34394 22392
rect 35618 22380 35624 22392
rect 35676 22380 35682 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 9217 22219 9275 22225
rect 9217 22185 9229 22219
rect 9263 22216 9275 22219
rect 9306 22216 9312 22228
rect 9263 22188 9312 22216
rect 9263 22185 9275 22188
rect 9217 22179 9275 22185
rect 9306 22176 9312 22188
rect 9364 22176 9370 22228
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 15010 22216 15016 22228
rect 14884 22188 15016 22216
rect 14884 22176 14890 22188
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15746 22176 15752 22228
rect 15804 22216 15810 22228
rect 15841 22219 15899 22225
rect 15841 22216 15853 22219
rect 15804 22188 15853 22216
rect 15804 22176 15810 22188
rect 15841 22185 15853 22188
rect 15887 22185 15899 22219
rect 15841 22179 15899 22185
rect 15930 22176 15936 22228
rect 15988 22216 15994 22228
rect 25498 22216 25504 22228
rect 15988 22188 25504 22216
rect 15988 22176 15994 22188
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 26132 22219 26190 22225
rect 26132 22185 26144 22219
rect 26178 22216 26190 22219
rect 26786 22216 26792 22228
rect 26178 22188 26792 22216
rect 26178 22185 26190 22188
rect 26132 22179 26190 22185
rect 26786 22176 26792 22188
rect 26844 22176 26850 22228
rect 32214 22176 32220 22228
rect 32272 22216 32278 22228
rect 32398 22216 32404 22228
rect 32272 22188 32404 22216
rect 32272 22176 32278 22188
rect 32398 22176 32404 22188
rect 32456 22176 32462 22228
rect 36630 22216 36636 22228
rect 34624 22188 36636 22216
rect 21450 22108 21456 22160
rect 21508 22148 21514 22160
rect 25130 22148 25136 22160
rect 21508 22120 25136 22148
rect 21508 22108 21514 22120
rect 25130 22108 25136 22120
rect 25188 22108 25194 22160
rect 25332 22120 26004 22148
rect 7742 22080 7748 22092
rect 1964 22052 7748 22080
rect 1964 22024 1992 22052
rect 7742 22040 7748 22052
rect 7800 22040 7806 22092
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11609 22083 11667 22089
rect 11609 22080 11621 22083
rect 11296 22052 11621 22080
rect 11296 22040 11302 22052
rect 11609 22049 11621 22052
rect 11655 22049 11667 22083
rect 12066 22080 12072 22092
rect 12027 22052 12072 22080
rect 11609 22043 11667 22049
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22080 15439 22083
rect 18874 22080 18880 22092
rect 15427 22052 18880 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 24949 22083 25007 22089
rect 24949 22080 24961 22083
rect 22066 22052 24961 22080
rect 1946 22012 1952 22024
rect 1907 21984 1952 22012
rect 1946 21972 1952 21984
rect 2004 21972 2010 22024
rect 6822 21972 6828 22024
rect 6880 22012 6886 22024
rect 8205 22015 8263 22021
rect 8205 22012 8217 22015
rect 6880 21984 8217 22012
rect 6880 21972 6886 21984
rect 8205 21981 8217 21984
rect 8251 21981 8263 22015
rect 8205 21975 8263 21981
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 10873 22015 10931 22021
rect 10873 21981 10885 22015
rect 10919 22012 10931 22015
rect 11422 22012 11428 22024
rect 10919 21984 11428 22012
rect 10919 21981 10931 21984
rect 10873 21975 10931 21981
rect 6638 21904 6644 21956
rect 6696 21944 6702 21956
rect 9140 21944 9168 21975
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 6696 21916 9168 21944
rect 11701 21947 11759 21953
rect 6696 21904 6702 21916
rect 6886 21888 6914 21916
rect 11701 21913 11713 21947
rect 11747 21913 11759 21947
rect 14366 21944 14372 21956
rect 14327 21916 14372 21944
rect 11701 21907 11759 21913
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 1765 21879 1823 21885
rect 1765 21876 1777 21879
rect 1636 21848 1777 21876
rect 1636 21836 1642 21848
rect 1765 21845 1777 21848
rect 1811 21845 1823 21879
rect 1765 21839 1823 21845
rect 6822 21836 6828 21888
rect 6880 21848 6914 21888
rect 8297 21879 8355 21885
rect 6880 21836 6886 21848
rect 8297 21845 8309 21879
rect 8343 21876 8355 21879
rect 10870 21876 10876 21888
rect 8343 21848 10876 21876
rect 8343 21845 8355 21848
rect 8297 21839 8355 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 10965 21879 11023 21885
rect 10965 21845 10977 21879
rect 11011 21876 11023 21879
rect 11716 21876 11744 21907
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14461 21947 14519 21953
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 15286 21944 15292 21956
rect 14507 21916 15292 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 16040 21944 16068 21975
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 17402 22012 17408 22024
rect 16632 21984 17408 22012
rect 16632 21972 16638 21984
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 21726 21972 21732 22024
rect 21784 22012 21790 22024
rect 22066 22012 22094 22052
rect 24949 22049 24961 22052
rect 24995 22049 25007 22083
rect 25332 22080 25360 22120
rect 24949 22043 25007 22049
rect 25148 22052 25360 22080
rect 25869 22083 25927 22089
rect 21784 21984 22094 22012
rect 24857 22015 24915 22021
rect 21784 21972 21790 21984
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25148 22012 25176 22052
rect 25869 22049 25881 22083
rect 25915 22049 25927 22083
rect 25976 22080 26004 22120
rect 31294 22108 31300 22160
rect 31352 22148 31358 22160
rect 31352 22120 32720 22148
rect 31352 22108 31358 22120
rect 26602 22080 26608 22092
rect 25976 22052 26608 22080
rect 25869 22043 25927 22049
rect 24903 21984 25176 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 22830 21944 22836 21956
rect 16040 21916 22836 21944
rect 22830 21904 22836 21916
rect 22888 21904 22894 21956
rect 24762 21904 24768 21956
rect 24820 21944 24826 21956
rect 25884 21944 25912 22043
rect 26602 22040 26608 22052
rect 26660 22080 26666 22092
rect 28261 22083 28319 22089
rect 28261 22080 28273 22083
rect 26660 22052 28273 22080
rect 26660 22040 26666 22052
rect 28261 22049 28273 22052
rect 28307 22049 28319 22083
rect 28261 22043 28319 22049
rect 32306 22040 32312 22092
rect 32364 22080 32370 22092
rect 32585 22083 32643 22089
rect 32585 22080 32597 22083
rect 32364 22052 32597 22080
rect 32364 22040 32370 22052
rect 32585 22049 32597 22052
rect 32631 22049 32643 22083
rect 32692 22080 32720 22120
rect 34624 22080 34652 22188
rect 36630 22176 36636 22188
rect 36688 22176 36694 22228
rect 36998 22176 37004 22228
rect 37056 22216 37062 22228
rect 37461 22219 37519 22225
rect 37461 22216 37473 22219
rect 37056 22188 37473 22216
rect 37056 22176 37062 22188
rect 37461 22185 37473 22188
rect 37507 22185 37519 22219
rect 37461 22179 37519 22185
rect 39850 22108 39856 22160
rect 39908 22148 39914 22160
rect 39908 22120 39988 22148
rect 39908 22108 39914 22120
rect 32692 22052 34652 22080
rect 32585 22043 32643 22049
rect 27982 21972 27988 22024
rect 28040 22012 28046 22024
rect 28077 22015 28135 22021
rect 28077 22012 28089 22015
rect 28040 21984 28089 22012
rect 28040 21972 28046 21984
rect 28077 21981 28089 21984
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 28997 22015 29055 22021
rect 28997 21981 29009 22015
rect 29043 22012 29055 22015
rect 29914 22012 29920 22024
rect 29043 21984 29920 22012
rect 29043 21981 29055 21984
rect 28997 21975 29055 21981
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 27430 21944 27436 21956
rect 24820 21916 25912 21944
rect 27370 21916 27436 21944
rect 24820 21904 24826 21916
rect 27430 21904 27436 21916
rect 27488 21904 27494 21956
rect 32861 21947 32919 21953
rect 32861 21913 32873 21947
rect 32907 21944 32919 21947
rect 32950 21944 32956 21956
rect 32907 21916 32956 21944
rect 32907 21913 32919 21916
rect 32861 21907 32919 21913
rect 32950 21904 32956 21916
rect 33008 21904 33014 21956
rect 34624 21944 34652 22052
rect 34790 22040 34796 22092
rect 34848 22080 34854 22092
rect 34885 22083 34943 22089
rect 34885 22080 34897 22083
rect 34848 22052 34897 22080
rect 34848 22040 34854 22052
rect 34885 22049 34897 22052
rect 34931 22049 34943 22083
rect 34885 22043 34943 22049
rect 35618 22040 35624 22092
rect 35676 22080 35682 22092
rect 36633 22083 36691 22089
rect 36633 22080 36645 22083
rect 35676 22052 36645 22080
rect 35676 22040 35682 22052
rect 36633 22049 36645 22052
rect 36679 22049 36691 22083
rect 39960 22080 39988 22120
rect 36633 22043 36691 22049
rect 37568 22052 39988 22080
rect 37369 22017 37427 22023
rect 37369 21983 37381 22017
rect 37415 22012 37427 22017
rect 37458 22012 37464 22024
rect 37415 21984 37464 22012
rect 37415 21983 37427 21984
rect 37369 21977 37427 21983
rect 37458 21972 37464 21984
rect 37516 21972 37522 22024
rect 35161 21947 35219 21953
rect 35161 21944 35173 21947
rect 34086 21916 34560 21944
rect 34624 21916 35173 21944
rect 11011 21848 11744 21876
rect 11011 21845 11023 21848
rect 10965 21839 11023 21845
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 17218 21876 17224 21888
rect 12032 21848 17224 21876
rect 12032 21836 12038 21848
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 17402 21836 17408 21888
rect 17460 21876 17466 21888
rect 23934 21876 23940 21888
rect 17460 21848 23940 21876
rect 17460 21836 17466 21848
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 24302 21836 24308 21888
rect 24360 21876 24366 21888
rect 25866 21876 25872 21888
rect 24360 21848 25872 21876
rect 24360 21836 24366 21848
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 27617 21879 27675 21885
rect 27617 21845 27629 21879
rect 27663 21876 27675 21879
rect 28718 21876 28724 21888
rect 27663 21848 28724 21876
rect 27663 21845 27675 21848
rect 27617 21839 27675 21845
rect 28718 21836 28724 21848
rect 28776 21836 28782 21888
rect 29089 21879 29147 21885
rect 29089 21845 29101 21879
rect 29135 21876 29147 21879
rect 29914 21876 29920 21888
rect 29135 21848 29920 21876
rect 29135 21845 29147 21848
rect 29089 21839 29147 21845
rect 29914 21836 29920 21848
rect 29972 21836 29978 21888
rect 33778 21836 33784 21888
rect 33836 21876 33842 21888
rect 34333 21879 34391 21885
rect 34333 21876 34345 21879
rect 33836 21848 34345 21876
rect 33836 21836 33842 21848
rect 34333 21845 34345 21848
rect 34379 21845 34391 21879
rect 34532 21876 34560 21916
rect 35161 21913 35173 21916
rect 35207 21913 35219 21947
rect 36998 21944 37004 21956
rect 36386 21916 37004 21944
rect 35161 21907 35219 21913
rect 36998 21904 37004 21916
rect 37056 21904 37062 21956
rect 37568 21876 37596 22052
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 34532 21848 37596 21876
rect 34333 21839 34391 21845
rect 37826 21836 37832 21888
rect 37884 21876 37890 21888
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 37884 21848 38117 21876
rect 37884 21836 37890 21848
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 14734 21672 14740 21684
rect 14695 21644 14740 21672
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 15381 21675 15439 21681
rect 15381 21672 15393 21675
rect 15344 21644 15393 21672
rect 15344 21632 15350 21644
rect 15381 21641 15393 21644
rect 15427 21641 15439 21675
rect 15381 21635 15439 21641
rect 20530 21632 20536 21684
rect 20588 21672 20594 21684
rect 20898 21672 20904 21684
rect 20588 21644 20904 21672
rect 20588 21632 20594 21644
rect 20898 21632 20904 21644
rect 20956 21632 20962 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 23477 21675 23535 21681
rect 23477 21672 23489 21675
rect 22520 21644 23489 21672
rect 22520 21632 22526 21644
rect 23477 21641 23489 21644
rect 23523 21641 23535 21675
rect 23477 21635 23535 21641
rect 24394 21632 24400 21684
rect 24452 21672 24458 21684
rect 24489 21675 24547 21681
rect 24489 21672 24501 21675
rect 24452 21644 24501 21672
rect 24452 21632 24458 21644
rect 24489 21641 24501 21644
rect 24535 21641 24547 21675
rect 25130 21672 25136 21684
rect 25091 21644 25136 21672
rect 24489 21635 24547 21641
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 25866 21632 25872 21684
rect 25924 21672 25930 21684
rect 25924 21644 28028 21672
rect 25924 21632 25930 21644
rect 10137 21607 10195 21613
rect 10137 21573 10149 21607
rect 10183 21604 10195 21607
rect 11054 21604 11060 21616
rect 10183 21576 11060 21604
rect 10183 21573 10195 21576
rect 10137 21567 10195 21573
rect 11054 21564 11060 21576
rect 11112 21564 11118 21616
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17276 21576 22094 21604
rect 17276 21564 17282 21576
rect 1578 21536 1584 21548
rect 1539 21508 1584 21536
rect 1578 21496 1584 21508
rect 1636 21496 1642 21548
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 6788 21508 8217 21536
rect 6788 21496 6794 21508
rect 8205 21505 8217 21508
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 12526 21536 12532 21548
rect 10735 21508 12532 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14691 21508 15301 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 15289 21505 15301 21508
rect 15335 21536 15347 21539
rect 20346 21536 20352 21548
rect 15335 21508 20352 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 22066 21536 22094 21576
rect 23290 21564 23296 21616
rect 23348 21604 23354 21616
rect 28000 21613 28028 21644
rect 33962 21632 33968 21684
rect 34020 21672 34026 21684
rect 34020 21644 37688 21672
rect 34020 21632 34026 21644
rect 26421 21607 26479 21613
rect 26421 21604 26433 21607
rect 23348 21576 26433 21604
rect 23348 21564 23354 21576
rect 26421 21573 26433 21576
rect 26467 21573 26479 21607
rect 26421 21567 26479 21573
rect 27985 21607 28043 21613
rect 27985 21573 27997 21607
rect 28031 21604 28043 21607
rect 28074 21604 28080 21616
rect 28031 21576 28080 21604
rect 28031 21573 28043 21576
rect 27985 21567 28043 21573
rect 28074 21564 28080 21576
rect 28132 21564 28138 21616
rect 28902 21604 28908 21616
rect 28863 21576 28908 21604
rect 28902 21564 28908 21576
rect 28960 21564 28966 21616
rect 34238 21564 34244 21616
rect 34296 21604 34302 21616
rect 35434 21604 35440 21616
rect 34296 21576 35440 21604
rect 34296 21564 34302 21576
rect 35434 21564 35440 21576
rect 35492 21564 35498 21616
rect 37274 21604 37280 21616
rect 36386 21576 37280 21604
rect 37274 21564 37280 21576
rect 37332 21564 37338 21616
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 22066 21508 23397 21536
rect 23385 21505 23397 21508
rect 23431 21536 23443 21539
rect 24302 21536 24308 21548
rect 23431 21508 24308 21536
rect 23431 21505 23443 21508
rect 23385 21499 23443 21505
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24397 21539 24455 21545
rect 24397 21505 24409 21539
rect 24443 21536 24455 21539
rect 24854 21536 24860 21548
rect 24443 21508 24860 21536
rect 24443 21505 24455 21508
rect 24397 21499 24455 21505
rect 24854 21496 24860 21508
rect 24912 21536 24918 21548
rect 25041 21539 25099 21545
rect 25041 21536 25053 21539
rect 24912 21508 25053 21536
rect 24912 21496 24918 21508
rect 25041 21505 25053 21508
rect 25087 21536 25099 21539
rect 25590 21536 25596 21548
rect 25087 21508 25596 21536
rect 25087 21505 25099 21508
rect 25041 21499 25099 21505
rect 25590 21496 25596 21508
rect 25648 21536 25654 21548
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 25648 21508 25697 21536
rect 25648 21496 25654 21508
rect 25685 21505 25697 21508
rect 25731 21536 25743 21539
rect 26329 21539 26387 21545
rect 26329 21536 26341 21539
rect 25731 21508 26341 21536
rect 25731 21505 25743 21508
rect 25685 21499 25743 21505
rect 26329 21505 26341 21508
rect 26375 21505 26387 21539
rect 26329 21499 26387 21505
rect 27062 21496 27068 21548
rect 27120 21536 27126 21548
rect 27617 21539 27675 21545
rect 27617 21536 27629 21539
rect 27120 21508 27629 21536
rect 27120 21496 27126 21508
rect 27617 21505 27629 21508
rect 27663 21505 27675 21539
rect 27617 21499 27675 21505
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21468 10103 21471
rect 10134 21468 10140 21480
rect 10091 21440 10140 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10134 21428 10140 21440
rect 10192 21428 10198 21480
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 17862 21468 17868 21480
rect 10928 21440 17868 21468
rect 10928 21428 10934 21440
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 22002 21428 22008 21480
rect 22060 21468 22066 21480
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 22060 21440 25789 21468
rect 22060 21428 22066 21440
rect 25777 21437 25789 21440
rect 25823 21437 25835 21471
rect 27632 21468 27660 21499
rect 34330 21496 34336 21548
rect 34388 21536 34394 21548
rect 34606 21536 34612 21548
rect 34388 21508 34612 21536
rect 34388 21496 34394 21508
rect 34606 21496 34612 21508
rect 34664 21496 34670 21548
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 37660 21545 37688 21644
rect 34885 21539 34943 21545
rect 34885 21536 34897 21539
rect 34848 21508 34897 21536
rect 34848 21496 34854 21508
rect 34885 21505 34897 21508
rect 34931 21505 34943 21539
rect 34885 21499 34943 21505
rect 37645 21539 37703 21545
rect 37645 21505 37657 21539
rect 37691 21505 37703 21539
rect 37645 21499 37703 21505
rect 27982 21468 27988 21480
rect 27632 21440 27988 21468
rect 25777 21431 25835 21437
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 28813 21471 28871 21477
rect 28813 21437 28825 21471
rect 28859 21437 28871 21471
rect 28813 21431 28871 21437
rect 23106 21360 23112 21412
rect 23164 21400 23170 21412
rect 23566 21400 23572 21412
rect 23164 21372 23572 21400
rect 23164 21360 23170 21372
rect 23566 21360 23572 21372
rect 23624 21400 23630 21412
rect 23624 21372 26556 21400
rect 23624 21360 23630 21372
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 8297 21335 8355 21341
rect 8297 21301 8309 21335
rect 8343 21332 8355 21335
rect 16942 21332 16948 21344
rect 8343 21304 16948 21332
rect 8343 21301 8355 21304
rect 8297 21295 8355 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 26418 21332 26424 21344
rect 21232 21304 26424 21332
rect 21232 21292 21238 21304
rect 26418 21292 26424 21304
rect 26476 21292 26482 21344
rect 26528 21332 26556 21372
rect 27614 21360 27620 21412
rect 27672 21400 27678 21412
rect 28828 21400 28856 21431
rect 29822 21428 29828 21480
rect 29880 21468 29886 21480
rect 31386 21468 31392 21480
rect 29880 21440 31392 21468
rect 29880 21428 29886 21440
rect 31386 21428 31392 21440
rect 31444 21468 31450 21480
rect 35161 21471 35219 21477
rect 35161 21468 35173 21471
rect 31444 21440 35173 21468
rect 31444 21428 31450 21440
rect 35161 21437 35173 21440
rect 35207 21437 35219 21471
rect 35161 21431 35219 21437
rect 37274 21428 37280 21480
rect 37332 21468 37338 21480
rect 38105 21471 38163 21477
rect 38105 21468 38117 21471
rect 37332 21440 38117 21468
rect 37332 21428 37338 21440
rect 38105 21437 38117 21440
rect 38151 21437 38163 21471
rect 38105 21431 38163 21437
rect 29362 21400 29368 21412
rect 27672 21372 28856 21400
rect 29323 21372 29368 21400
rect 27672 21360 27678 21372
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 29730 21360 29736 21412
rect 29788 21400 29794 21412
rect 30650 21400 30656 21412
rect 29788 21372 30656 21400
rect 29788 21360 29794 21372
rect 30650 21360 30656 21372
rect 30708 21360 30714 21412
rect 31846 21360 31852 21412
rect 31904 21400 31910 21412
rect 34330 21400 34336 21412
rect 31904 21372 34336 21400
rect 31904 21360 31910 21372
rect 34330 21360 34336 21372
rect 34388 21360 34394 21412
rect 36998 21360 37004 21412
rect 37056 21400 37062 21412
rect 37734 21400 37740 21412
rect 37056 21372 37740 21400
rect 37056 21360 37062 21372
rect 37734 21360 37740 21372
rect 37792 21360 37798 21412
rect 33962 21332 33968 21344
rect 26528 21304 33968 21332
rect 33962 21292 33968 21304
rect 34020 21292 34026 21344
rect 36170 21292 36176 21344
rect 36228 21332 36234 21344
rect 36630 21332 36636 21344
rect 36228 21304 36636 21332
rect 36228 21292 36234 21304
rect 36630 21292 36636 21304
rect 36688 21292 36694 21344
rect 37461 21335 37519 21341
rect 37461 21301 37473 21335
rect 37507 21332 37519 21335
rect 38286 21332 38292 21344
rect 37507 21304 38292 21332
rect 37507 21301 37519 21304
rect 37461 21295 37519 21301
rect 38286 21292 38292 21304
rect 38344 21292 38350 21344
rect 39666 21292 39672 21344
rect 39724 21292 39730 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 39684 21208 39712 21292
rect 1104 21168 38824 21190
rect 39666 21156 39672 21208
rect 39724 21156 39730 21208
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 9214 21128 9220 21140
rect 1627 21100 9220 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 11422 21088 11428 21140
rect 11480 21128 11486 21140
rect 19426 21128 19432 21140
rect 11480 21100 19432 21128
rect 11480 21088 11486 21100
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 20625 21131 20683 21137
rect 20625 21097 20637 21131
rect 20671 21128 20683 21131
rect 21910 21128 21916 21140
rect 20671 21100 21916 21128
rect 20671 21097 20683 21100
rect 20625 21091 20683 21097
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 22189 21131 22247 21137
rect 22189 21097 22201 21131
rect 22235 21128 22247 21131
rect 23382 21128 23388 21140
rect 22235 21100 23388 21128
rect 22235 21097 22247 21100
rect 22189 21091 22247 21097
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 25038 21088 25044 21140
rect 25096 21128 25102 21140
rect 25869 21131 25927 21137
rect 25869 21128 25881 21131
rect 25096 21100 25881 21128
rect 25096 21088 25102 21100
rect 25869 21097 25881 21100
rect 25915 21097 25927 21131
rect 25869 21091 25927 21097
rect 26142 21088 26148 21140
rect 26200 21088 26206 21140
rect 26418 21088 26424 21140
rect 26476 21128 26482 21140
rect 26513 21131 26571 21137
rect 26513 21128 26525 21131
rect 26476 21100 26525 21128
rect 26476 21088 26482 21100
rect 26513 21097 26525 21100
rect 26559 21097 26571 21131
rect 26513 21091 26571 21097
rect 30834 21088 30840 21140
rect 30892 21128 30898 21140
rect 32217 21131 32275 21137
rect 32217 21128 32229 21131
rect 30892 21100 32229 21128
rect 30892 21088 30898 21100
rect 32217 21097 32229 21100
rect 32263 21097 32275 21131
rect 33962 21128 33968 21140
rect 33923 21100 33968 21128
rect 32217 21091 32275 21097
rect 33962 21088 33968 21100
rect 34020 21088 34026 21140
rect 35894 21128 35900 21140
rect 35855 21100 35900 21128
rect 35894 21088 35900 21100
rect 35952 21088 35958 21140
rect 37274 21088 37280 21140
rect 37332 21088 37338 21140
rect 37458 21088 37464 21140
rect 37516 21128 37522 21140
rect 39574 21128 39580 21140
rect 37516 21100 39580 21128
rect 37516 21088 37522 21100
rect 39574 21088 39580 21100
rect 39632 21088 39638 21140
rect 3418 21020 3424 21072
rect 3476 21060 3482 21072
rect 23934 21060 23940 21072
rect 3476 21032 6914 21060
rect 3476 21020 3482 21032
rect 6886 20992 6914 21032
rect 17512 21032 23796 21060
rect 23895 21032 23940 21060
rect 17512 21001 17540 21032
rect 17497 20995 17555 21001
rect 17497 20992 17509 20995
rect 6886 20964 17509 20992
rect 17497 20961 17509 20964
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 21266 20952 21272 21004
rect 21324 20992 21330 21004
rect 21361 20995 21419 21001
rect 21361 20992 21373 20995
rect 21324 20964 21373 20992
rect 21324 20952 21330 20964
rect 21361 20961 21373 20964
rect 21407 20961 21419 20995
rect 23768 20992 23796 21032
rect 23934 21020 23940 21032
rect 23992 21060 23998 21072
rect 25225 21063 25283 21069
rect 25225 21060 25237 21063
rect 23992 21032 25237 21060
rect 23992 21020 23998 21032
rect 25225 21029 25237 21032
rect 25271 21029 25283 21063
rect 25225 21023 25283 21029
rect 25406 21020 25412 21072
rect 25464 21060 25470 21072
rect 26160 21060 26188 21088
rect 25464 21032 26188 21060
rect 25464 21020 25470 21032
rect 27338 21020 27344 21072
rect 27396 21060 27402 21072
rect 27396 21032 30972 21060
rect 27396 21020 27402 21032
rect 28169 20995 28227 21001
rect 28169 20992 28181 20995
rect 23768 20964 28181 20992
rect 21361 20955 21419 20961
rect 28169 20961 28181 20964
rect 28215 20961 28227 20995
rect 28442 20992 28448 21004
rect 28403 20964 28448 20992
rect 28169 20955 28227 20961
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 30653 20995 30711 21001
rect 30653 20961 30665 20995
rect 30699 20992 30711 20995
rect 30742 20992 30748 21004
rect 30699 20964 30748 20992
rect 30699 20961 30711 20964
rect 30653 20955 30711 20961
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 30944 21001 30972 21032
rect 33134 21020 33140 21072
rect 33192 21060 33198 21072
rect 33870 21060 33876 21072
rect 33192 21032 33876 21060
rect 33192 21020 33198 21032
rect 33870 21020 33876 21032
rect 33928 21020 33934 21072
rect 34238 21020 34244 21072
rect 34296 21060 34302 21072
rect 34422 21060 34428 21072
rect 34296 21032 34428 21060
rect 34296 21020 34302 21032
rect 34422 21020 34428 21032
rect 34480 21020 34486 21072
rect 30929 20995 30987 21001
rect 30929 20961 30941 20995
rect 30975 20992 30987 20995
rect 30975 20964 31616 20992
rect 30975 20961 30987 20964
rect 30929 20955 30987 20961
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 16482 20924 16488 20936
rect 16443 20896 16488 20924
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 20530 20924 20536 20936
rect 20491 20896 20536 20924
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22186 20924 22192 20936
rect 22143 20896 22192 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 17221 20859 17279 20865
rect 17221 20825 17233 20859
rect 17267 20825 17279 20859
rect 17221 20819 17279 20825
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 16577 20791 16635 20797
rect 16577 20788 16589 20791
rect 15252 20760 16589 20788
rect 15252 20748 15258 20760
rect 16577 20757 16589 20760
rect 16623 20757 16635 20791
rect 16577 20751 16635 20757
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17236 20788 17264 20819
rect 17310 20816 17316 20868
rect 17368 20856 17374 20868
rect 17368 20828 17413 20856
rect 17368 20816 17374 20828
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 21192 20856 21220 20887
rect 22186 20884 22192 20896
rect 22244 20884 22250 20936
rect 25777 20927 25835 20933
rect 25777 20893 25789 20927
rect 25823 20893 25835 20927
rect 25777 20887 25835 20893
rect 22646 20856 22652 20868
rect 19300 20828 22652 20856
rect 19300 20816 19306 20828
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 23106 20816 23112 20868
rect 23164 20856 23170 20868
rect 23374 20859 23432 20865
rect 23374 20856 23386 20859
rect 23164 20828 23386 20856
rect 23164 20816 23170 20828
rect 23374 20825 23386 20828
rect 23420 20825 23432 20859
rect 23374 20819 23432 20825
rect 23470 20859 23528 20865
rect 23470 20825 23482 20859
rect 23516 20856 23528 20859
rect 23658 20856 23664 20868
rect 23516 20828 23664 20856
rect 23516 20825 23528 20828
rect 23470 20819 23528 20825
rect 23658 20816 23664 20828
rect 23716 20816 23722 20868
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 24670 20856 24676 20868
rect 24176 20828 24676 20856
rect 24176 20816 24182 20828
rect 24670 20816 24676 20828
rect 24728 20816 24734 20868
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20825 24823 20859
rect 24765 20819 24823 20825
rect 17184 20760 17264 20788
rect 17184 20748 17190 20760
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 20346 20788 20352 20800
rect 19484 20760 20352 20788
rect 19484 20748 19490 20760
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 22922 20748 22928 20800
rect 22980 20788 22986 20800
rect 24780 20788 24808 20819
rect 24854 20816 24860 20868
rect 24912 20856 24918 20868
rect 25792 20856 25820 20887
rect 25866 20884 25872 20936
rect 25924 20924 25930 20936
rect 25924 20896 26280 20924
rect 25924 20884 25930 20896
rect 24912 20828 25820 20856
rect 26252 20856 26280 20896
rect 26326 20884 26332 20936
rect 26384 20924 26390 20936
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26384 20896 26433 20924
rect 26384 20884 26390 20896
rect 26421 20893 26433 20896
rect 26467 20924 26479 20927
rect 26602 20924 26608 20936
rect 26467 20896 26608 20924
rect 26467 20893 26479 20896
rect 26421 20887 26479 20893
rect 26602 20884 26608 20896
rect 26660 20884 26666 20936
rect 27062 20924 27068 20936
rect 27023 20896 27068 20924
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 27341 20859 27399 20865
rect 27341 20856 27353 20859
rect 26252 20828 27353 20856
rect 24912 20816 24918 20828
rect 27341 20825 27353 20828
rect 27387 20825 27399 20859
rect 27341 20819 27399 20825
rect 28261 20859 28319 20865
rect 28261 20825 28273 20859
rect 28307 20856 28319 20859
rect 28994 20856 29000 20868
rect 28307 20828 29000 20856
rect 28307 20825 28319 20828
rect 28261 20819 28319 20825
rect 22980 20760 24808 20788
rect 27356 20788 27384 20819
rect 28994 20816 29000 20828
rect 29052 20816 29058 20868
rect 29546 20816 29552 20868
rect 29604 20856 29610 20868
rect 30745 20859 30803 20865
rect 30745 20856 30757 20859
rect 29604 20828 30757 20856
rect 29604 20816 29610 20828
rect 30745 20825 30757 20828
rect 30791 20825 30803 20859
rect 30745 20819 30803 20825
rect 28442 20788 28448 20800
rect 27356 20760 28448 20788
rect 22980 20748 22986 20760
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 29825 20791 29883 20797
rect 29825 20757 29837 20791
rect 29871 20788 29883 20791
rect 30834 20788 30840 20800
rect 29871 20760 30840 20788
rect 29871 20757 29883 20760
rect 29825 20751 29883 20757
rect 30834 20748 30840 20760
rect 30892 20748 30898 20800
rect 31588 20788 31616 20964
rect 31662 20952 31668 21004
rect 31720 20992 31726 21004
rect 37292 21001 37320 21088
rect 36541 20995 36599 21001
rect 36541 20992 36553 20995
rect 31720 20964 36553 20992
rect 31720 20952 31726 20964
rect 36541 20961 36553 20964
rect 36587 20961 36599 20995
rect 36541 20955 36599 20961
rect 37277 20995 37335 21001
rect 37277 20961 37289 20995
rect 37323 20961 37335 20995
rect 37277 20955 37335 20961
rect 37458 20952 37464 21004
rect 37516 20992 37522 21004
rect 37553 20995 37611 21001
rect 37553 20992 37565 20995
rect 37516 20964 37565 20992
rect 37516 20952 37522 20964
rect 37553 20961 37565 20964
rect 37599 20961 37611 20995
rect 37553 20955 37611 20961
rect 38102 20952 38108 21004
rect 38160 20992 38166 21004
rect 38746 20992 38752 21004
rect 38160 20964 38752 20992
rect 38160 20952 38166 20964
rect 38746 20952 38752 20964
rect 38804 20952 38810 21004
rect 32122 20924 32128 20936
rect 32083 20896 32128 20924
rect 32122 20884 32128 20896
rect 32180 20884 32186 20936
rect 32490 20884 32496 20936
rect 32548 20924 32554 20936
rect 33229 20927 33287 20933
rect 33229 20924 33241 20927
rect 32548 20896 33241 20924
rect 32548 20884 32554 20896
rect 33229 20893 33241 20896
rect 33275 20893 33287 20927
rect 33229 20887 33287 20893
rect 33502 20884 33508 20936
rect 33560 20924 33566 20936
rect 33778 20924 33784 20936
rect 33560 20896 33784 20924
rect 33560 20884 33566 20896
rect 33778 20884 33784 20896
rect 33836 20884 33842 20936
rect 33870 20884 33876 20936
rect 33928 20924 33934 20936
rect 33928 20896 33973 20924
rect 33928 20884 33934 20896
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 35161 20927 35219 20933
rect 35161 20924 35173 20927
rect 34204 20896 35173 20924
rect 34204 20884 34210 20896
rect 35161 20893 35173 20896
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 35805 20927 35863 20933
rect 35805 20893 35817 20927
rect 35851 20924 35863 20927
rect 35986 20924 35992 20936
rect 35851 20896 35992 20924
rect 35851 20893 35863 20896
rect 35805 20887 35863 20893
rect 35986 20884 35992 20896
rect 36044 20884 36050 20936
rect 36446 20924 36452 20936
rect 36407 20896 36452 20924
rect 36446 20884 36452 20896
rect 36504 20884 36510 20936
rect 33321 20859 33379 20865
rect 33321 20825 33333 20859
rect 33367 20856 33379 20859
rect 34790 20856 34796 20868
rect 33367 20828 34796 20856
rect 33367 20825 33379 20828
rect 33321 20819 33379 20825
rect 34790 20816 34796 20828
rect 34848 20816 34854 20868
rect 37366 20856 37372 20868
rect 37327 20828 37372 20856
rect 37366 20816 37372 20828
rect 37424 20816 37430 20868
rect 35158 20788 35164 20800
rect 31588 20760 35164 20788
rect 35158 20748 35164 20760
rect 35216 20748 35222 20800
rect 35253 20791 35311 20797
rect 35253 20757 35265 20791
rect 35299 20788 35311 20791
rect 35802 20788 35808 20800
rect 35299 20760 35808 20788
rect 35299 20757 35311 20760
rect 35253 20751 35311 20757
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 20990 20584 20996 20596
rect 6687 20556 7512 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7484 20457 7512 20556
rect 18432 20556 20996 20584
rect 16942 20516 16948 20528
rect 16903 20488 16948 20516
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 17037 20519 17095 20525
rect 17037 20485 17049 20519
rect 17083 20516 17095 20519
rect 18322 20516 18328 20528
rect 17083 20488 18328 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 18432 20457 18460 20556
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 21269 20587 21327 20593
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 23658 20584 23664 20596
rect 21315 20556 23664 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 23842 20584 23848 20596
rect 23803 20556 23848 20584
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 24578 20544 24584 20596
rect 24636 20584 24642 20596
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 24636 20556 25053 20584
rect 24636 20544 24642 20556
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 28902 20584 28908 20596
rect 25041 20547 25099 20553
rect 25516 20556 28764 20584
rect 28863 20556 28908 20584
rect 25516 20516 25544 20556
rect 19168 20488 25544 20516
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 14645 20383 14703 20389
rect 14645 20380 14657 20383
rect 14608 20352 14657 20380
rect 14608 20340 14614 20352
rect 14645 20349 14657 20352
rect 14691 20349 14703 20383
rect 14645 20343 14703 20349
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17644 20352 17877 20380
rect 17644 20340 17650 20352
rect 17865 20349 17877 20352
rect 17911 20380 17923 20383
rect 19168 20380 19196 20488
rect 26142 20476 26148 20528
rect 26200 20516 26206 20528
rect 26200 20488 26245 20516
rect 26200 20476 26206 20488
rect 26418 20476 26424 20528
rect 26476 20516 26482 20528
rect 27433 20519 27491 20525
rect 27433 20516 27445 20519
rect 26476 20488 27445 20516
rect 26476 20476 26482 20488
rect 27433 20485 27445 20488
rect 27479 20485 27491 20519
rect 27433 20479 27491 20485
rect 21177 20451 21235 20457
rect 21177 20417 21189 20451
rect 21223 20448 21235 20451
rect 22554 20448 22560 20460
rect 21223 20420 22560 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 22704 20420 22749 20448
rect 22704 20408 22710 20420
rect 22830 20408 22836 20460
rect 22888 20448 22894 20460
rect 23753 20451 23811 20457
rect 22888 20420 23244 20448
rect 22888 20408 22894 20420
rect 17911 20352 19196 20380
rect 17911 20349 17923 20352
rect 17865 20343 17923 20349
rect 21818 20340 21824 20392
rect 21876 20380 21882 20392
rect 23216 20389 23244 20420
rect 23753 20417 23765 20451
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 23201 20383 23259 20389
rect 21876 20352 23152 20380
rect 21876 20340 21882 20352
rect 7282 20312 7288 20324
rect 7243 20284 7288 20312
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 13262 20272 13268 20324
rect 13320 20312 13326 20324
rect 13722 20312 13728 20324
rect 13320 20284 13728 20312
rect 13320 20272 13326 20284
rect 13722 20272 13728 20284
rect 13780 20312 13786 20324
rect 22094 20312 22100 20324
rect 13780 20284 22100 20312
rect 13780 20272 13786 20284
rect 22094 20272 22100 20284
rect 22152 20272 22158 20324
rect 22370 20272 22376 20324
rect 22428 20312 22434 20324
rect 22830 20312 22836 20324
rect 22428 20284 22836 20312
rect 22428 20272 22434 20284
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 23124 20312 23152 20352
rect 23201 20349 23213 20383
rect 23247 20380 23259 20383
rect 23290 20380 23296 20392
rect 23247 20352 23296 20380
rect 23247 20349 23259 20352
rect 23201 20343 23259 20349
rect 23290 20340 23296 20352
rect 23348 20340 23354 20392
rect 23566 20340 23572 20392
rect 23624 20380 23630 20392
rect 23768 20380 23796 20411
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24912 20420 24961 20448
rect 24912 20408 24918 20420
rect 24949 20417 24961 20420
rect 24995 20417 25007 20451
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 24949 20411 25007 20417
rect 25056 20420 26065 20448
rect 25056 20380 25084 20420
rect 26053 20417 26065 20420
rect 26099 20448 26111 20451
rect 26326 20448 26332 20460
rect 26099 20420 26332 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26326 20408 26332 20420
rect 26384 20408 26390 20460
rect 23624 20352 25084 20380
rect 23624 20340 23630 20352
rect 25866 20340 25872 20392
rect 25924 20380 25930 20392
rect 27341 20383 27399 20389
rect 27341 20380 27353 20383
rect 25924 20352 27353 20380
rect 25924 20340 25930 20352
rect 27341 20349 27353 20352
rect 27387 20349 27399 20383
rect 27614 20380 27620 20392
rect 27575 20352 27620 20380
rect 27341 20343 27399 20349
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 28736 20380 28764 20556
rect 28902 20544 28908 20556
rect 28960 20544 28966 20596
rect 29546 20584 29552 20596
rect 29507 20556 29552 20584
rect 29546 20544 29552 20556
rect 29604 20544 29610 20596
rect 30374 20544 30380 20596
rect 30432 20584 30438 20596
rect 33045 20587 33103 20593
rect 33045 20584 33057 20587
rect 30432 20556 33057 20584
rect 30432 20544 30438 20556
rect 33045 20553 33057 20556
rect 33091 20553 33103 20587
rect 33045 20547 33103 20553
rect 33778 20544 33784 20596
rect 33836 20584 33842 20596
rect 34146 20584 34152 20596
rect 33836 20556 34152 20584
rect 33836 20544 33842 20556
rect 34146 20544 34152 20556
rect 34204 20544 34210 20596
rect 35342 20544 35348 20596
rect 35400 20584 35406 20596
rect 35529 20587 35587 20593
rect 35529 20584 35541 20587
rect 35400 20556 35541 20584
rect 35400 20544 35406 20556
rect 35529 20553 35541 20556
rect 35575 20553 35587 20587
rect 35529 20547 35587 20553
rect 36078 20544 36084 20596
rect 36136 20584 36142 20596
rect 36173 20587 36231 20593
rect 36173 20584 36185 20587
rect 36136 20556 36185 20584
rect 36136 20544 36142 20556
rect 36173 20553 36185 20556
rect 36219 20553 36231 20587
rect 38194 20584 38200 20596
rect 38155 20556 38200 20584
rect 36173 20547 36231 20553
rect 38194 20544 38200 20556
rect 38252 20544 38258 20596
rect 29178 20516 29184 20528
rect 28828 20488 29184 20516
rect 28828 20457 28856 20488
rect 29178 20476 29184 20488
rect 29236 20476 29242 20528
rect 30834 20516 30840 20528
rect 30795 20488 30840 20516
rect 30834 20476 30840 20488
rect 30892 20476 30898 20528
rect 32122 20476 32128 20528
rect 32180 20516 32186 20528
rect 34057 20519 34115 20525
rect 32180 20488 32996 20516
rect 32180 20476 32186 20488
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 29086 20408 29092 20460
rect 29144 20448 29150 20460
rect 29457 20451 29515 20457
rect 29457 20448 29469 20451
rect 29144 20420 29469 20448
rect 29144 20408 29150 20420
rect 29457 20417 29469 20420
rect 29503 20417 29515 20451
rect 29457 20411 29515 20417
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20448 32367 20451
rect 32398 20448 32404 20460
rect 32355 20420 32404 20448
rect 32355 20417 32367 20420
rect 32309 20411 32367 20417
rect 32398 20408 32404 20420
rect 32456 20408 32462 20460
rect 32968 20457 32996 20488
rect 34057 20485 34069 20519
rect 34103 20516 34115 20519
rect 35618 20516 35624 20528
rect 34103 20488 35624 20516
rect 34103 20485 34115 20488
rect 34057 20479 34115 20485
rect 35618 20476 35624 20488
rect 35676 20476 35682 20528
rect 32953 20451 33011 20457
rect 32953 20417 32965 20451
rect 32999 20448 33011 20451
rect 35437 20451 35495 20457
rect 32999 20420 33088 20448
rect 32999 20417 33011 20420
rect 32953 20411 33011 20417
rect 29730 20380 29736 20392
rect 28736 20352 29736 20380
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 30742 20380 30748 20392
rect 30703 20352 30748 20380
rect 30742 20340 30748 20352
rect 30800 20340 30806 20392
rect 31757 20383 31815 20389
rect 31757 20349 31769 20383
rect 31803 20380 31815 20383
rect 31846 20380 31852 20392
rect 31803 20352 31852 20380
rect 31803 20349 31815 20352
rect 31757 20343 31815 20349
rect 31772 20312 31800 20343
rect 31846 20340 31852 20352
rect 31904 20340 31910 20392
rect 23124 20284 31800 20312
rect 33060 20312 33088 20420
rect 35437 20417 35449 20451
rect 35483 20417 35495 20451
rect 35437 20411 35495 20417
rect 36081 20451 36139 20457
rect 36081 20417 36093 20451
rect 36127 20448 36139 20451
rect 36446 20448 36452 20460
rect 36127 20420 36452 20448
rect 36127 20417 36139 20420
rect 36081 20411 36139 20417
rect 33962 20380 33968 20392
rect 33923 20352 33968 20380
rect 33962 20340 33968 20352
rect 34020 20340 34026 20392
rect 34146 20340 34152 20392
rect 34204 20380 34210 20392
rect 34241 20383 34299 20389
rect 34241 20380 34253 20383
rect 34204 20352 34253 20380
rect 34204 20340 34210 20352
rect 34241 20349 34253 20352
rect 34287 20349 34299 20383
rect 34241 20343 34299 20349
rect 35452 20312 35480 20411
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 36722 20448 36728 20460
rect 36556 20420 36728 20448
rect 35526 20340 35532 20392
rect 35584 20380 35590 20392
rect 36556 20380 36584 20420
rect 36722 20408 36728 20420
rect 36780 20408 36786 20460
rect 38010 20448 38016 20460
rect 37971 20420 38016 20448
rect 38010 20408 38016 20420
rect 38068 20408 38074 20460
rect 35584 20352 36584 20380
rect 35584 20340 35590 20352
rect 33060 20284 35480 20312
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 18138 20244 18144 20256
rect 11756 20216 18144 20244
rect 11756 20204 11762 20216
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 19610 20244 19616 20256
rect 18555 20216 19616 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 32306 20244 32312 20256
rect 20128 20216 32312 20244
rect 20128 20204 20134 20216
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 32401 20247 32459 20253
rect 32401 20213 32413 20247
rect 32447 20244 32459 20247
rect 32490 20244 32496 20256
rect 32447 20216 32496 20244
rect 32447 20213 32459 20216
rect 32401 20207 32459 20213
rect 32490 20204 32496 20216
rect 32548 20204 32554 20256
rect 33686 20204 33692 20256
rect 33744 20244 33750 20256
rect 36817 20247 36875 20253
rect 36817 20244 36829 20247
rect 33744 20216 36829 20244
rect 33744 20204 33750 20216
rect 36817 20213 36829 20216
rect 36863 20213 36875 20247
rect 36817 20207 36875 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 14090 20000 14096 20052
rect 14148 20040 14154 20052
rect 21726 20040 21732 20052
rect 14148 20012 21732 20040
rect 14148 20000 14154 20012
rect 21726 20000 21732 20012
rect 21784 20000 21790 20052
rect 21818 20000 21824 20052
rect 21876 20040 21882 20052
rect 22922 20040 22928 20052
rect 21876 20012 22928 20040
rect 21876 20000 21882 20012
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 23017 20043 23075 20049
rect 23017 20009 23029 20043
rect 23063 20040 23075 20043
rect 23198 20040 23204 20052
rect 23063 20012 23204 20040
rect 23063 20009 23075 20012
rect 23017 20003 23075 20009
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 23661 20043 23719 20049
rect 23661 20009 23673 20043
rect 23707 20040 23719 20043
rect 23750 20040 23756 20052
rect 23707 20012 23756 20040
rect 23707 20009 23719 20012
rect 23661 20003 23719 20009
rect 23750 20000 23756 20012
rect 23808 20000 23814 20052
rect 25958 20000 25964 20052
rect 26016 20040 26022 20052
rect 26145 20043 26203 20049
rect 26145 20040 26157 20043
rect 26016 20012 26157 20040
rect 26016 20000 26022 20012
rect 26145 20009 26157 20012
rect 26191 20009 26203 20043
rect 26145 20003 26203 20009
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 28813 20043 28871 20049
rect 28813 20040 28825 20043
rect 27580 20012 28825 20040
rect 27580 20000 27586 20012
rect 28813 20009 28825 20012
rect 28859 20009 28871 20043
rect 28813 20003 28871 20009
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 32122 20040 32128 20052
rect 28960 20012 32128 20040
rect 28960 20000 28966 20012
rect 32122 20000 32128 20012
rect 32180 20000 32186 20052
rect 34146 20000 34152 20052
rect 34204 20040 34210 20052
rect 34204 20012 38148 20040
rect 34204 20000 34210 20012
rect 13630 19932 13636 19984
rect 13688 19972 13694 19984
rect 19426 19972 19432 19984
rect 13688 19944 19432 19972
rect 13688 19932 13694 19944
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 14844 19913 14872 19944
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 20070 19972 20076 19984
rect 20031 19944 20076 19972
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 22940 19944 30052 19972
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 22940 19904 22968 19944
rect 17552 19876 22968 19904
rect 17552 19864 17558 19876
rect 23014 19864 23020 19916
rect 23072 19904 23078 19916
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 23072 19876 24685 19904
rect 23072 19864 23078 19876
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 27154 19864 27160 19916
rect 27212 19904 27218 19916
rect 27433 19907 27491 19913
rect 27433 19904 27445 19907
rect 27212 19876 27445 19904
rect 27212 19864 27218 19876
rect 27433 19873 27445 19876
rect 27479 19873 27491 19907
rect 28166 19904 28172 19916
rect 28127 19876 28172 19904
rect 27433 19867 27491 19873
rect 20622 19836 20628 19848
rect 20583 19808 20628 19836
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 20772 19808 21557 19836
rect 20772 19796 20778 19808
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19836 21695 19839
rect 21818 19836 21824 19848
rect 21683 19808 21824 19836
rect 21683 19805 21695 19808
rect 21637 19799 21695 19805
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 22925 19839 22983 19845
rect 22925 19805 22937 19839
rect 22971 19836 22983 19839
rect 23566 19836 23572 19848
rect 22971 19808 23572 19836
rect 22971 19805 22983 19808
rect 22925 19799 22983 19805
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 24854 19836 24860 19848
rect 24627 19808 24860 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 26053 19839 26111 19845
rect 26053 19805 26065 19839
rect 26099 19836 26111 19839
rect 26326 19836 26332 19848
rect 26099 19808 26332 19836
rect 26099 19805 26111 19808
rect 26053 19799 26111 19805
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 11790 19768 11796 19780
rect 11751 19740 11796 19768
rect 11790 19728 11796 19740
rect 11848 19728 11854 19780
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 12802 19768 12808 19780
rect 11940 19740 11985 19768
rect 12763 19740 12808 19768
rect 11940 19728 11946 19740
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 14645 19771 14703 19777
rect 14645 19737 14657 19771
rect 14691 19768 14703 19771
rect 15194 19768 15200 19780
rect 14691 19740 15200 19768
rect 14691 19737 14703 19740
rect 14645 19731 14703 19737
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 17920 19740 19533 19768
rect 17920 19728 17926 19740
rect 19521 19737 19533 19740
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 11698 19700 11704 19712
rect 1912 19672 11704 19700
rect 1912 19660 1918 19672
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 13078 19660 13084 19712
rect 13136 19700 13142 19712
rect 13265 19703 13323 19709
rect 13265 19700 13277 19703
rect 13136 19672 13277 19700
rect 13136 19660 13142 19672
rect 13265 19669 13277 19672
rect 13311 19669 13323 19703
rect 19536 19700 19564 19731
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 26694 19768 26700 19780
rect 19668 19740 19713 19768
rect 26655 19740 26700 19768
rect 19668 19728 19674 19740
rect 26694 19728 26700 19740
rect 26752 19728 26758 19780
rect 27448 19768 27476 19867
rect 28166 19864 28172 19876
rect 28224 19864 28230 19916
rect 29730 19904 29736 19916
rect 29691 19876 29736 19904
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 29914 19904 29920 19916
rect 29875 19876 29920 19904
rect 29914 19864 29920 19876
rect 29972 19864 29978 19916
rect 30024 19904 30052 19944
rect 31846 19932 31852 19984
rect 31904 19972 31910 19984
rect 35342 19972 35348 19984
rect 31904 19944 35348 19972
rect 31904 19932 31910 19944
rect 35342 19932 35348 19944
rect 35400 19972 35406 19984
rect 37458 19972 37464 19984
rect 35400 19944 37464 19972
rect 35400 19932 35406 19944
rect 37458 19932 37464 19944
rect 37516 19932 37522 19984
rect 31573 19907 31631 19913
rect 30024 19876 31156 19904
rect 28074 19836 28080 19848
rect 28035 19808 28080 19836
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 28721 19839 28779 19845
rect 28721 19836 28733 19839
rect 28500 19808 28733 19836
rect 28500 19796 28506 19808
rect 28721 19805 28733 19808
rect 28767 19836 28779 19839
rect 28902 19836 28908 19848
rect 28767 19808 28908 19836
rect 28767 19805 28779 19808
rect 28721 19799 28779 19805
rect 28902 19796 28908 19808
rect 28960 19796 28966 19848
rect 31128 19836 31156 19876
rect 31573 19873 31585 19907
rect 31619 19904 31631 19907
rect 33870 19904 33876 19916
rect 31619 19876 33876 19904
rect 31619 19873 31631 19876
rect 31573 19867 31631 19873
rect 33870 19864 33876 19876
rect 33928 19864 33934 19916
rect 34977 19907 35035 19913
rect 34977 19904 34989 19907
rect 34808 19876 34989 19904
rect 34808 19848 34836 19876
rect 34977 19873 34989 19876
rect 35023 19873 35035 19907
rect 35250 19904 35256 19916
rect 35211 19876 35256 19904
rect 34977 19867 35035 19873
rect 35250 19864 35256 19876
rect 35308 19904 35314 19916
rect 35308 19876 35756 19904
rect 35308 19864 35314 19876
rect 31662 19836 31668 19848
rect 31128 19808 31668 19836
rect 31662 19796 31668 19808
rect 31720 19796 31726 19848
rect 32030 19836 32036 19848
rect 31991 19808 32036 19836
rect 32030 19796 32036 19808
rect 32088 19796 32094 19848
rect 34790 19796 34796 19848
rect 34848 19796 34854 19848
rect 35728 19836 35756 19876
rect 35802 19864 35808 19916
rect 35860 19904 35866 19916
rect 38120 19913 38148 20012
rect 36449 19907 36507 19913
rect 36449 19904 36461 19907
rect 35860 19876 36461 19904
rect 35860 19864 35866 19876
rect 36449 19873 36461 19876
rect 36495 19873 36507 19907
rect 36449 19867 36507 19873
rect 38105 19907 38163 19913
rect 38105 19873 38117 19907
rect 38151 19904 38163 19907
rect 39390 19904 39396 19916
rect 38151 19876 39396 19904
rect 38151 19873 38163 19876
rect 38105 19867 38163 19873
rect 39390 19864 39396 19876
rect 39448 19864 39454 19916
rect 36170 19836 36176 19848
rect 35728 19808 36176 19836
rect 36170 19796 36176 19808
rect 36228 19796 36234 19848
rect 36265 19839 36323 19845
rect 36265 19805 36277 19839
rect 36311 19805 36323 19839
rect 36265 19799 36323 19805
rect 28092 19768 28120 19796
rect 29454 19768 29460 19780
rect 27448 19740 27660 19768
rect 28092 19740 29460 19768
rect 20070 19700 20076 19712
rect 19536 19672 20076 19700
rect 13265 19663 13323 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20714 19700 20720 19712
rect 20675 19672 20720 19700
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 27632 19700 27660 19740
rect 29454 19728 29460 19740
rect 29512 19728 29518 19780
rect 32214 19768 32220 19780
rect 32175 19740 32220 19768
rect 32214 19728 32220 19740
rect 32272 19728 32278 19780
rect 35069 19771 35127 19777
rect 35069 19737 35081 19771
rect 35115 19768 35127 19771
rect 35158 19768 35164 19780
rect 35115 19740 35164 19768
rect 35115 19737 35127 19740
rect 35069 19731 35127 19737
rect 35158 19728 35164 19740
rect 35216 19728 35222 19780
rect 35894 19728 35900 19780
rect 35952 19768 35958 19780
rect 36280 19768 36308 19799
rect 35952 19740 36308 19768
rect 35952 19728 35958 19740
rect 29086 19700 29092 19712
rect 27632 19672 29092 19700
rect 29086 19660 29092 19672
rect 29144 19700 29150 19712
rect 30834 19700 30840 19712
rect 29144 19672 30840 19700
rect 29144 19660 29150 19672
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 31570 19660 31576 19712
rect 31628 19700 31634 19712
rect 33778 19700 33784 19712
rect 31628 19672 33784 19700
rect 31628 19660 31634 19672
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 34422 19660 34428 19712
rect 34480 19700 34486 19712
rect 34606 19700 34612 19712
rect 34480 19672 34612 19700
rect 34480 19660 34486 19672
rect 34606 19660 34612 19672
rect 34664 19660 34670 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 21358 19496 21364 19508
rect 21319 19468 21364 19496
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 21450 19456 21456 19508
rect 21508 19496 21514 19508
rect 26234 19496 26240 19508
rect 21508 19468 26096 19496
rect 26195 19468 26240 19496
rect 21508 19456 21514 19468
rect 13078 19428 13084 19440
rect 13039 19400 13084 19428
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 13173 19431 13231 19437
rect 13173 19397 13185 19431
rect 13219 19428 13231 19431
rect 16482 19428 16488 19440
rect 13219 19400 16488 19428
rect 13219 19397 13231 19400
rect 13173 19391 13231 19397
rect 16482 19388 16488 19400
rect 16540 19388 16546 19440
rect 16942 19428 16948 19440
rect 16903 19400 16948 19428
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 17037 19431 17095 19437
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 19150 19428 19156 19440
rect 17083 19400 19156 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 19245 19431 19303 19437
rect 19245 19397 19257 19431
rect 19291 19428 19303 19431
rect 19291 19400 20576 19428
rect 19291 19397 19303 19400
rect 19245 19391 19303 19397
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 9769 19363 9827 19369
rect 9769 19360 9781 19363
rect 8352 19332 9781 19360
rect 8352 19320 8358 19332
rect 9769 19329 9781 19332
rect 9815 19329 9827 19363
rect 9769 19323 9827 19329
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 12342 19360 12348 19372
rect 9907 19332 12348 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 17862 19360 17868 19372
rect 17604 19332 17868 19360
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 13722 19292 13728 19304
rect 13683 19264 13728 19292
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 17604 19292 17632 19332
rect 17862 19320 17868 19332
rect 17920 19360 17926 19372
rect 17920 19332 19012 19360
rect 17920 19320 17926 19332
rect 15028 19264 17632 19292
rect 18984 19292 19012 19332
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18984 19264 19165 19292
rect 13354 19184 13360 19236
rect 13412 19224 13418 19236
rect 15028 19224 15056 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19426 19292 19432 19304
rect 19387 19264 19432 19292
rect 19153 19255 19211 19261
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 20548 19292 20576 19400
rect 20714 19388 20720 19440
rect 20772 19428 20778 19440
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 20772 19400 22201 19428
rect 20772 19388 20778 19400
rect 22189 19397 22201 19400
rect 22235 19397 22247 19431
rect 22189 19391 22247 19397
rect 25593 19431 25651 19437
rect 25593 19397 25605 19431
rect 25639 19428 25651 19431
rect 25958 19428 25964 19440
rect 25639 19400 25964 19428
rect 25639 19397 25651 19400
rect 25593 19391 25651 19397
rect 25958 19388 25964 19400
rect 26016 19388 26022 19440
rect 26068 19428 26096 19468
rect 26234 19456 26240 19468
rect 26292 19456 26298 19508
rect 26344 19468 37780 19496
rect 26344 19428 26372 19468
rect 26068 19400 26372 19428
rect 27249 19431 27307 19437
rect 27249 19397 27261 19431
rect 27295 19428 27307 19431
rect 27890 19428 27896 19440
rect 27295 19400 27896 19428
rect 27295 19397 27307 19400
rect 27249 19391 27307 19397
rect 27890 19388 27896 19400
rect 27948 19388 27954 19440
rect 28994 19388 29000 19440
rect 29052 19428 29058 19440
rect 29917 19431 29975 19437
rect 29917 19428 29929 19431
rect 29052 19400 29929 19428
rect 29052 19388 29058 19400
rect 29917 19397 29929 19400
rect 29963 19397 29975 19431
rect 30650 19428 30656 19440
rect 30611 19400 30656 19428
rect 29917 19391 29975 19397
rect 30650 19388 30656 19400
rect 30708 19388 30714 19440
rect 31570 19428 31576 19440
rect 31531 19400 31576 19428
rect 31570 19388 31576 19400
rect 31628 19388 31634 19440
rect 31662 19388 31668 19440
rect 31720 19428 31726 19440
rect 34146 19428 34152 19440
rect 31720 19400 34152 19428
rect 31720 19388 31726 19400
rect 34146 19388 34152 19400
rect 34204 19388 34210 19440
rect 34790 19428 34796 19440
rect 34751 19400 34796 19428
rect 34790 19388 34796 19400
rect 34848 19388 34854 19440
rect 35250 19388 35256 19440
rect 35308 19428 35314 19440
rect 35894 19428 35900 19440
rect 35308 19400 35900 19428
rect 35308 19388 35314 19400
rect 35894 19388 35900 19400
rect 35952 19388 35958 19440
rect 36078 19388 36084 19440
rect 36136 19428 36142 19440
rect 36265 19431 36323 19437
rect 36265 19428 36277 19431
rect 36136 19400 36277 19428
rect 36136 19388 36142 19400
rect 36265 19397 36277 19400
rect 36311 19397 36323 19431
rect 36265 19391 36323 19397
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19360 20683 19363
rect 21082 19360 21088 19372
rect 20671 19332 21088 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21266 19360 21272 19372
rect 21227 19332 21272 19360
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 25498 19360 25504 19372
rect 25459 19332 25504 19360
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 25832 19332 26157 19360
rect 25832 19320 25838 19332
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26418 19360 26424 19372
rect 26292 19332 26424 19360
rect 26292 19320 26298 19332
rect 26418 19320 26424 19332
rect 26476 19320 26482 19372
rect 27154 19360 27160 19372
rect 27115 19332 27160 19360
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 27982 19360 27988 19372
rect 27943 19332 27988 19360
rect 27982 19320 27988 19332
rect 28040 19360 28046 19372
rect 28905 19363 28963 19369
rect 28905 19360 28917 19363
rect 28040 19332 28917 19360
rect 28040 19320 28046 19332
rect 28905 19329 28917 19332
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19360 29239 19363
rect 29227 19332 29592 19360
rect 29227 19329 29239 19332
rect 29181 19323 29239 19329
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20548 19264 20729 19292
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 20717 19255 20775 19261
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 28074 19292 28080 19304
rect 22152 19264 22197 19292
rect 22572 19264 28080 19292
rect 22152 19252 22158 19264
rect 13412 19196 15056 19224
rect 13412 19184 13418 19196
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 17497 19227 17555 19233
rect 17497 19224 17509 19227
rect 15160 19196 17509 19224
rect 15160 19184 15166 19196
rect 17497 19193 17509 19196
rect 17543 19224 17555 19227
rect 22572 19224 22600 19264
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 28261 19295 28319 19301
rect 28261 19261 28273 19295
rect 28307 19292 28319 19295
rect 28350 19292 28356 19304
rect 28307 19264 28356 19292
rect 28307 19261 28319 19264
rect 28261 19255 28319 19261
rect 28350 19252 28356 19264
rect 28408 19252 28414 19304
rect 29564 19292 29592 19332
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 29825 19363 29883 19369
rect 29825 19360 29837 19363
rect 29696 19332 29837 19360
rect 29696 19320 29702 19332
rect 29825 19329 29837 19332
rect 29871 19329 29883 19363
rect 30374 19360 30380 19372
rect 29825 19323 29883 19329
rect 29932 19332 30380 19360
rect 29932 19292 29960 19332
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 32030 19320 32036 19372
rect 32088 19360 32094 19372
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 32088 19332 32321 19360
rect 32088 19320 32094 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 36170 19360 36176 19372
rect 36131 19332 36176 19360
rect 32309 19323 32367 19329
rect 36170 19320 36176 19332
rect 36228 19320 36234 19372
rect 37752 19369 37780 19468
rect 37737 19363 37795 19369
rect 37737 19329 37749 19363
rect 37783 19329 37795 19363
rect 37737 19323 37795 19329
rect 29564 19264 29960 19292
rect 30561 19295 30619 19301
rect 30561 19261 30573 19295
rect 30607 19261 30619 19295
rect 32490 19292 32496 19304
rect 32451 19264 32496 19292
rect 30561 19255 30619 19261
rect 17543 19196 22600 19224
rect 22649 19227 22707 19233
rect 17543 19193 17555 19196
rect 17497 19187 17555 19193
rect 22649 19193 22661 19227
rect 22695 19224 22707 19227
rect 27338 19224 27344 19236
rect 22695 19196 27344 19224
rect 22695 19193 22707 19196
rect 22649 19187 22707 19193
rect 27338 19184 27344 19196
rect 27396 19184 27402 19236
rect 27522 19184 27528 19236
rect 27580 19224 27586 19236
rect 27580 19196 29224 19224
rect 27580 19184 27586 19196
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 23934 19156 23940 19168
rect 20128 19128 23940 19156
rect 20128 19116 20134 19128
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 29086 19156 29092 19168
rect 25740 19128 29092 19156
rect 25740 19116 25746 19128
rect 29086 19116 29092 19128
rect 29144 19116 29150 19168
rect 29196 19156 29224 19196
rect 29914 19184 29920 19236
rect 29972 19224 29978 19236
rect 30576 19224 30604 19255
rect 32490 19252 32496 19264
rect 32548 19252 32554 19304
rect 34701 19295 34759 19301
rect 34701 19292 34713 19295
rect 32876 19264 34713 19292
rect 29972 19196 30604 19224
rect 29972 19184 29978 19196
rect 32306 19184 32312 19236
rect 32364 19224 32370 19236
rect 32766 19224 32772 19236
rect 32364 19196 32772 19224
rect 32364 19184 32370 19196
rect 32766 19184 32772 19196
rect 32824 19184 32830 19236
rect 31294 19156 31300 19168
rect 29196 19128 31300 19156
rect 31294 19116 31300 19128
rect 31352 19116 31358 19168
rect 31662 19116 31668 19168
rect 31720 19156 31726 19168
rect 32876 19156 32904 19264
rect 34624 19236 34652 19264
rect 34701 19261 34713 19264
rect 34747 19261 34759 19295
rect 34974 19292 34980 19304
rect 34935 19264 34980 19292
rect 34701 19255 34759 19261
rect 34974 19252 34980 19264
rect 35032 19252 35038 19304
rect 37458 19292 37464 19304
rect 37419 19264 37464 19292
rect 37458 19252 37464 19264
rect 37516 19252 37522 19304
rect 34606 19184 34612 19236
rect 34664 19184 34670 19236
rect 35250 19224 35256 19236
rect 34716 19196 35256 19224
rect 31720 19128 32904 19156
rect 31720 19116 31726 19128
rect 34146 19116 34152 19168
rect 34204 19156 34210 19168
rect 34716 19156 34744 19196
rect 35250 19184 35256 19196
rect 35308 19184 35314 19236
rect 34204 19128 34744 19156
rect 34204 19116 34210 19128
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 14366 18952 14372 18964
rect 13679 18924 14372 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18417 18955 18475 18961
rect 18417 18952 18429 18955
rect 18380 18924 18429 18952
rect 18380 18912 18386 18924
rect 18417 18921 18429 18924
rect 18463 18921 18475 18955
rect 18417 18915 18475 18921
rect 19150 18912 19156 18964
rect 19208 18952 19214 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19208 18924 19533 18952
rect 19208 18912 19214 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 20070 18912 20076 18964
rect 20128 18952 20134 18964
rect 20346 18952 20352 18964
rect 20128 18924 20352 18952
rect 20128 18912 20134 18924
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 25130 18912 25136 18964
rect 25188 18952 25194 18964
rect 27338 18952 27344 18964
rect 25188 18924 27344 18952
rect 25188 18912 25194 18924
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 27430 18912 27436 18964
rect 27488 18952 27494 18964
rect 29825 18955 29883 18961
rect 29825 18952 29837 18955
rect 27488 18924 29837 18952
rect 27488 18912 27494 18924
rect 29825 18921 29837 18924
rect 29871 18921 29883 18955
rect 29825 18915 29883 18921
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 31113 18955 31171 18961
rect 31113 18952 31125 18955
rect 30524 18924 31125 18952
rect 30524 18912 30530 18924
rect 31113 18921 31125 18924
rect 31159 18921 31171 18955
rect 31113 18915 31171 18921
rect 31757 18955 31815 18961
rect 31757 18921 31769 18955
rect 31803 18952 31815 18955
rect 33226 18952 33232 18964
rect 31803 18924 33232 18952
rect 31803 18921 31815 18924
rect 31757 18915 31815 18921
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 33686 18952 33692 18964
rect 33647 18924 33692 18952
rect 33686 18912 33692 18924
rect 33744 18912 33750 18964
rect 36906 18952 36912 18964
rect 36867 18924 36912 18952
rect 36906 18912 36912 18924
rect 36964 18912 36970 18964
rect 37642 18912 37648 18964
rect 37700 18952 37706 18964
rect 38197 18955 38255 18961
rect 38197 18952 38209 18955
rect 37700 18924 38209 18952
rect 37700 18912 37706 18924
rect 38197 18921 38209 18924
rect 38243 18921 38255 18955
rect 38197 18915 38255 18921
rect 12526 18884 12532 18896
rect 11808 18856 12532 18884
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 11808 18757 11836 18856
rect 12526 18844 12532 18856
rect 12584 18884 12590 18896
rect 13170 18884 13176 18896
rect 12584 18856 13176 18884
rect 12584 18844 12590 18856
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 15102 18884 15108 18896
rect 15063 18856 15108 18884
rect 15102 18844 15108 18856
rect 15160 18844 15166 18896
rect 15562 18844 15568 18896
rect 15620 18884 15626 18896
rect 32398 18884 32404 18896
rect 15620 18856 31754 18884
rect 32359 18856 32404 18884
rect 15620 18844 15626 18856
rect 12342 18776 12348 18828
rect 12400 18816 12406 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 12400 18788 14565 18816
rect 12400 18776 12406 18788
rect 14553 18785 14565 18788
rect 14599 18816 14611 18819
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 14599 18788 16589 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 17586 18816 17592 18828
rect 17547 18788 17592 18816
rect 16577 18779 16635 18785
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 19518 18776 19524 18828
rect 19576 18816 19582 18828
rect 20714 18816 20720 18828
rect 19576 18788 20720 18816
rect 19576 18776 19582 18788
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 23934 18776 23940 18828
rect 23992 18816 23998 18828
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 23992 18788 25881 18816
rect 23992 18776 23998 18788
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 25869 18779 25927 18785
rect 26326 18776 26332 18828
rect 26384 18816 26390 18828
rect 27154 18816 27160 18828
rect 26384 18788 27160 18816
rect 26384 18776 26390 18788
rect 27154 18776 27160 18788
rect 27212 18816 27218 18828
rect 31726 18816 31754 18856
rect 32398 18844 32404 18856
rect 32456 18844 32462 18896
rect 32766 18844 32772 18896
rect 32824 18884 32830 18896
rect 33042 18884 33048 18896
rect 32824 18856 33048 18884
rect 32824 18844 32830 18856
rect 33042 18844 33048 18856
rect 33100 18844 33106 18896
rect 34698 18844 34704 18896
rect 34756 18884 34762 18896
rect 35710 18884 35716 18896
rect 34756 18856 35716 18884
rect 34756 18844 34762 18856
rect 35710 18844 35716 18856
rect 35768 18844 35774 18896
rect 37553 18887 37611 18893
rect 37553 18853 37565 18887
rect 37599 18884 37611 18887
rect 38930 18884 38936 18896
rect 37599 18856 38936 18884
rect 37599 18853 37611 18856
rect 37553 18847 37611 18853
rect 38930 18844 38936 18856
rect 38988 18844 38994 18896
rect 35621 18819 35679 18825
rect 35621 18816 35633 18819
rect 27212 18788 30420 18816
rect 31726 18788 35633 18816
rect 27212 18776 27218 18788
rect 30392 18760 30420 18788
rect 35621 18785 35633 18788
rect 35667 18816 35679 18819
rect 35894 18816 35900 18828
rect 35667 18788 35900 18816
rect 35667 18785 35679 18788
rect 35621 18779 35679 18785
rect 35894 18776 35900 18788
rect 35952 18776 35958 18828
rect 35986 18776 35992 18828
rect 36044 18816 36050 18828
rect 36044 18788 36860 18816
rect 36044 18776 36050 18788
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1728 18720 1961 18748
rect 1728 18708 1734 18720
rect 1949 18717 1961 18720
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 12676 18720 13553 18748
rect 12676 18708 12682 18720
rect 13541 18717 13553 18720
rect 13587 18717 13599 18751
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 13541 18711 13599 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 24762 18748 24768 18760
rect 19475 18720 24768 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25130 18748 25136 18760
rect 25091 18720 25136 18748
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 27062 18708 27068 18760
rect 27120 18748 27126 18760
rect 27430 18748 27436 18760
rect 27120 18720 27436 18748
rect 27120 18708 27126 18720
rect 27430 18708 27436 18720
rect 27488 18708 27494 18760
rect 28534 18748 28540 18760
rect 28495 18720 28540 18748
rect 28534 18708 28540 18720
rect 28592 18708 28598 18760
rect 28902 18708 28908 18760
rect 28960 18748 28966 18760
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 28960 18720 29745 18748
rect 28960 18708 28966 18720
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 30374 18748 30380 18760
rect 30335 18720 30380 18748
rect 29733 18711 29791 18717
rect 30374 18708 30380 18720
rect 30432 18708 30438 18760
rect 30466 18708 30472 18760
rect 30524 18748 30530 18760
rect 31021 18751 31079 18757
rect 31021 18748 31033 18751
rect 30524 18720 31033 18748
rect 30524 18708 30530 18720
rect 31021 18717 31033 18720
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 9306 18640 9312 18692
rect 9364 18680 9370 18692
rect 10597 18683 10655 18689
rect 10597 18680 10609 18683
rect 9364 18652 10609 18680
rect 9364 18640 9370 18652
rect 10597 18649 10609 18652
rect 10643 18649 10655 18683
rect 10597 18643 10655 18649
rect 10689 18683 10747 18689
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 11054 18680 11060 18692
rect 10735 18652 11060 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 11241 18683 11299 18689
rect 11241 18649 11253 18683
rect 11287 18680 11299 18683
rect 13722 18680 13728 18692
rect 11287 18652 13728 18680
rect 11287 18649 11299 18652
rect 11241 18643 11299 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 14642 18640 14648 18692
rect 14700 18680 14706 18692
rect 16669 18683 16727 18689
rect 14700 18652 14745 18680
rect 14700 18640 14706 18652
rect 16669 18649 16681 18683
rect 16715 18680 16727 18683
rect 17494 18680 17500 18692
rect 16715 18652 17500 18680
rect 16715 18649 16727 18652
rect 16669 18643 16727 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 20162 18640 20168 18692
rect 20220 18680 20226 18692
rect 20346 18680 20352 18692
rect 20220 18652 20352 18680
rect 20220 18640 20226 18652
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 25682 18680 25688 18692
rect 22066 18652 25688 18680
rect 11885 18615 11943 18621
rect 11885 18581 11897 18615
rect 11931 18612 11943 18615
rect 12158 18612 12164 18624
rect 11931 18584 12164 18612
rect 11931 18581 11943 18584
rect 11885 18575 11943 18581
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 14366 18612 14372 18624
rect 14240 18584 14372 18612
rect 14240 18572 14246 18584
rect 14366 18572 14372 18584
rect 14424 18612 14430 18624
rect 22066 18612 22094 18652
rect 25682 18640 25688 18652
rect 25740 18640 25746 18692
rect 25961 18683 26019 18689
rect 25961 18649 25973 18683
rect 26007 18649 26019 18683
rect 26878 18680 26884 18692
rect 26839 18652 26884 18680
rect 25961 18643 26019 18649
rect 14424 18584 22094 18612
rect 25225 18615 25283 18621
rect 14424 18572 14430 18584
rect 25225 18581 25237 18615
rect 25271 18612 25283 18615
rect 25976 18612 26004 18643
rect 26878 18640 26884 18652
rect 26936 18640 26942 18692
rect 27890 18680 27896 18692
rect 27851 18652 27896 18680
rect 27890 18640 27896 18652
rect 27948 18680 27954 18692
rect 28442 18680 28448 18692
rect 27948 18652 28448 18680
rect 27948 18640 27954 18652
rect 28442 18640 28448 18652
rect 28500 18640 28506 18692
rect 28810 18640 28816 18692
rect 28868 18680 28874 18692
rect 31036 18680 31064 18711
rect 31570 18708 31576 18760
rect 31628 18748 31634 18760
rect 31665 18753 31723 18759
rect 31665 18748 31677 18753
rect 31628 18720 31677 18748
rect 31628 18708 31634 18720
rect 31665 18719 31677 18720
rect 31711 18719 31723 18753
rect 31665 18713 31723 18719
rect 32309 18751 32367 18757
rect 32309 18717 32321 18751
rect 32355 18748 32367 18751
rect 32950 18748 32956 18760
rect 32355 18720 32956 18748
rect 32355 18717 32367 18720
rect 32309 18711 32367 18717
rect 32950 18708 32956 18720
rect 33008 18708 33014 18760
rect 33226 18708 33232 18760
rect 33284 18748 33290 18760
rect 36832 18757 36860 18788
rect 33597 18751 33655 18757
rect 33597 18748 33609 18751
rect 33284 18720 33609 18748
rect 33284 18708 33290 18720
rect 33597 18717 33609 18720
rect 33643 18717 33655 18751
rect 33597 18711 33655 18717
rect 36817 18751 36875 18757
rect 36817 18717 36829 18751
rect 36863 18748 36875 18751
rect 37461 18751 37519 18757
rect 37461 18748 37473 18751
rect 36863 18720 37473 18748
rect 36863 18717 36875 18720
rect 36817 18711 36875 18717
rect 37461 18717 37473 18720
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 38010 18708 38016 18760
rect 38068 18748 38074 18760
rect 38105 18751 38163 18757
rect 38105 18748 38117 18751
rect 38068 18720 38117 18748
rect 38068 18708 38074 18720
rect 38105 18717 38117 18720
rect 38151 18748 38163 18751
rect 39574 18748 39580 18760
rect 38151 18720 39580 18748
rect 38151 18717 38163 18720
rect 38105 18711 38163 18717
rect 39574 18708 39580 18720
rect 39632 18708 39638 18760
rect 31110 18680 31116 18692
rect 28868 18652 30512 18680
rect 31036 18652 31116 18680
rect 28868 18640 28874 18652
rect 25271 18584 26004 18612
rect 25271 18581 25283 18584
rect 25225 18575 25283 18581
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 30484 18621 30512 18652
rect 31110 18640 31116 18652
rect 31168 18640 31174 18692
rect 32582 18640 32588 18692
rect 32640 18680 32646 18692
rect 33045 18683 33103 18689
rect 33045 18680 33057 18683
rect 32640 18652 33057 18680
rect 32640 18640 32646 18652
rect 33045 18649 33057 18652
rect 33091 18649 33103 18683
rect 33045 18643 33103 18649
rect 34606 18640 34612 18692
rect 34664 18680 34670 18692
rect 35345 18683 35403 18689
rect 35345 18680 35357 18683
rect 34664 18652 35357 18680
rect 34664 18640 34670 18652
rect 35345 18649 35357 18652
rect 35391 18649 35403 18683
rect 35345 18643 35403 18649
rect 35437 18683 35495 18689
rect 35437 18649 35449 18683
rect 35483 18680 35495 18683
rect 36262 18680 36268 18692
rect 35483 18652 36268 18680
rect 35483 18649 35495 18652
rect 35437 18643 35495 18649
rect 36262 18640 36268 18652
rect 36320 18640 36326 18692
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 27396 18584 28641 18612
rect 27396 18572 27402 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 28629 18575 28687 18581
rect 30469 18615 30527 18621
rect 30469 18581 30481 18615
rect 30515 18581 30527 18615
rect 30469 18575 30527 18581
rect 30834 18572 30840 18624
rect 30892 18612 30898 18624
rect 31570 18612 31576 18624
rect 30892 18584 31576 18612
rect 30892 18572 30898 18584
rect 31570 18572 31576 18584
rect 31628 18572 31634 18624
rect 33870 18572 33876 18624
rect 33928 18612 33934 18624
rect 36170 18612 36176 18624
rect 33928 18584 36176 18612
rect 33928 18572 33934 18584
rect 36170 18572 36176 18584
rect 36228 18572 36234 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 8294 18408 8300 18420
rect 1627 18380 8300 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 16025 18411 16083 18417
rect 16025 18408 16037 18411
rect 14700 18380 16037 18408
rect 14700 18368 14706 18380
rect 16025 18377 16037 18380
rect 16071 18377 16083 18411
rect 17494 18408 17500 18420
rect 17455 18380 17500 18408
rect 16025 18371 16083 18377
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 26418 18408 26424 18420
rect 18380 18380 26424 18408
rect 18380 18368 18386 18380
rect 26418 18368 26424 18380
rect 26476 18368 26482 18420
rect 26510 18368 26516 18420
rect 26568 18408 26574 18420
rect 28445 18411 28503 18417
rect 28445 18408 28457 18411
rect 26568 18380 28457 18408
rect 26568 18368 26574 18380
rect 28445 18377 28457 18380
rect 28491 18377 28503 18411
rect 29086 18408 29092 18420
rect 29047 18380 29092 18408
rect 28445 18371 28503 18377
rect 29086 18368 29092 18380
rect 29144 18368 29150 18420
rect 30190 18408 30196 18420
rect 30024 18380 30196 18408
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 11974 18340 11980 18352
rect 11848 18312 11980 18340
rect 11848 18300 11854 18312
rect 11974 18300 11980 18312
rect 12032 18340 12038 18352
rect 12345 18343 12403 18349
rect 12345 18340 12357 18343
rect 12032 18312 12357 18340
rect 12032 18300 12038 18312
rect 12345 18309 12357 18312
rect 12391 18309 12403 18343
rect 12345 18303 12403 18309
rect 12437 18343 12495 18349
rect 12437 18309 12449 18343
rect 12483 18340 12495 18343
rect 14182 18340 14188 18352
rect 12483 18312 14188 18340
rect 12483 18309 12495 18312
rect 12437 18303 12495 18309
rect 14182 18300 14188 18312
rect 14240 18300 14246 18352
rect 14461 18343 14519 18349
rect 14461 18309 14473 18343
rect 14507 18340 14519 18343
rect 14826 18340 14832 18352
rect 14507 18312 14832 18340
rect 14507 18309 14519 18312
rect 14461 18303 14519 18309
rect 14826 18300 14832 18312
rect 14884 18300 14890 18352
rect 18874 18300 18880 18352
rect 18932 18340 18938 18352
rect 19797 18343 19855 18349
rect 19797 18340 19809 18343
rect 18932 18312 19809 18340
rect 18932 18300 18938 18312
rect 19797 18309 19809 18312
rect 19843 18309 19855 18343
rect 19797 18303 19855 18309
rect 19889 18343 19947 18349
rect 19889 18309 19901 18343
rect 19935 18340 19947 18343
rect 20162 18340 20168 18352
rect 19935 18312 20168 18340
rect 19935 18309 19947 18312
rect 19889 18303 19947 18309
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 20714 18300 20720 18352
rect 20772 18340 20778 18352
rect 20809 18343 20867 18349
rect 20809 18340 20821 18343
rect 20772 18312 20821 18340
rect 20772 18300 20778 18312
rect 20809 18309 20821 18312
rect 20855 18309 20867 18343
rect 24854 18340 24860 18352
rect 24767 18312 24860 18340
rect 20809 18303 20867 18309
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 15930 18272 15936 18284
rect 15843 18244 15936 18272
rect 15930 18232 15936 18244
rect 15988 18272 15994 18284
rect 16390 18272 16396 18284
rect 15988 18244 16396 18272
rect 15988 18232 15994 18244
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18272 17463 18275
rect 19426 18272 19432 18284
rect 17451 18244 19432 18272
rect 17451 18241 17463 18244
rect 17405 18235 17463 18241
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 24780 18281 24808 18312
rect 24854 18300 24860 18312
rect 24912 18340 24918 18352
rect 27062 18340 27068 18352
rect 24912 18312 27068 18340
rect 24912 18300 24918 18312
rect 27062 18300 27068 18312
rect 27120 18300 27126 18352
rect 27338 18340 27344 18352
rect 27299 18312 27344 18340
rect 27338 18300 27344 18312
rect 27396 18300 27402 18352
rect 29178 18300 29184 18352
rect 29236 18340 29242 18352
rect 30024 18349 30052 18380
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 31573 18411 31631 18417
rect 31573 18408 31585 18411
rect 30708 18380 31585 18408
rect 30708 18368 30714 18380
rect 31573 18377 31585 18380
rect 31619 18377 31631 18411
rect 31573 18371 31631 18377
rect 32214 18368 32220 18420
rect 32272 18408 32278 18420
rect 32401 18411 32459 18417
rect 32401 18408 32413 18411
rect 32272 18380 32413 18408
rect 32272 18368 32278 18380
rect 32401 18377 32413 18380
rect 32447 18377 32459 18411
rect 34330 18408 34336 18420
rect 34291 18380 34336 18408
rect 32401 18371 32459 18377
rect 34330 18368 34336 18380
rect 34388 18368 34394 18420
rect 34790 18368 34796 18420
rect 34848 18408 34854 18420
rect 34977 18411 35035 18417
rect 34977 18408 34989 18411
rect 34848 18380 34989 18408
rect 34848 18368 34854 18380
rect 34977 18377 34989 18380
rect 35023 18377 35035 18411
rect 35618 18408 35624 18420
rect 35579 18380 35624 18408
rect 34977 18371 35035 18377
rect 35618 18368 35624 18380
rect 35676 18368 35682 18420
rect 36262 18408 36268 18420
rect 36223 18380 36268 18408
rect 36262 18368 36268 18380
rect 36320 18368 36326 18420
rect 37461 18411 37519 18417
rect 37461 18377 37473 18411
rect 37507 18408 37519 18411
rect 37550 18408 37556 18420
rect 37507 18380 37556 18408
rect 37507 18377 37519 18380
rect 37461 18371 37519 18377
rect 37550 18368 37556 18380
rect 37608 18368 37614 18420
rect 30009 18343 30067 18349
rect 30009 18340 30021 18343
rect 29236 18312 30021 18340
rect 29236 18300 29242 18312
rect 30009 18309 30021 18312
rect 30055 18309 30067 18343
rect 30009 18303 30067 18309
rect 30101 18343 30159 18349
rect 30101 18309 30113 18343
rect 30147 18340 30159 18343
rect 30466 18340 30472 18352
rect 30147 18312 30472 18340
rect 30147 18309 30159 18312
rect 30101 18303 30159 18309
rect 30466 18300 30472 18312
rect 30524 18300 30530 18352
rect 31938 18300 31944 18352
rect 31996 18340 32002 18352
rect 33689 18343 33747 18349
rect 33689 18340 33701 18343
rect 31996 18312 33701 18340
rect 31996 18300 32002 18312
rect 33689 18309 33701 18312
rect 33735 18309 33747 18343
rect 36630 18340 36636 18352
rect 33689 18303 33747 18309
rect 35544 18312 36636 18340
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18241 24823 18275
rect 24765 18235 24823 18241
rect 26237 18275 26295 18281
rect 26237 18241 26249 18275
rect 26283 18272 26295 18275
rect 26970 18272 26976 18284
rect 26283 18244 26976 18272
rect 26283 18241 26295 18244
rect 26237 18235 26295 18241
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 28350 18272 28356 18284
rect 28311 18244 28356 18272
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29052 18244 29097 18272
rect 29052 18232 29058 18244
rect 31386 18232 31392 18284
rect 31444 18272 31450 18284
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31444 18244 31493 18272
rect 31444 18232 31450 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 31846 18232 31852 18284
rect 31904 18272 31910 18284
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 31904 18244 32321 18272
rect 31904 18232 31910 18244
rect 32309 18241 32321 18244
rect 32355 18241 32367 18275
rect 32950 18272 32956 18284
rect 32911 18244 32956 18272
rect 32309 18235 32367 18241
rect 32950 18232 32956 18244
rect 33008 18232 33014 18284
rect 33597 18275 33655 18281
rect 33597 18241 33609 18275
rect 33643 18272 33655 18275
rect 33870 18272 33876 18284
rect 33643 18244 33876 18272
rect 33643 18241 33655 18244
rect 33597 18235 33655 18241
rect 33870 18232 33876 18244
rect 33928 18232 33934 18284
rect 35544 18281 35572 18312
rect 36630 18300 36636 18312
rect 36688 18300 36694 18352
rect 34241 18275 34299 18281
rect 34241 18241 34253 18275
rect 34287 18241 34299 18275
rect 34241 18235 34299 18241
rect 34885 18275 34943 18281
rect 34885 18241 34897 18275
rect 34931 18241 34943 18275
rect 34885 18235 34943 18241
rect 35529 18275 35587 18281
rect 35529 18241 35541 18275
rect 35575 18241 35587 18275
rect 35529 18235 35587 18241
rect 13354 18204 13360 18216
rect 13315 18176 13360 18204
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 16298 18164 16304 18216
rect 16356 18204 16362 18216
rect 23566 18204 23572 18216
rect 16356 18176 23572 18204
rect 16356 18164 16362 18176
rect 23566 18164 23572 18176
rect 23624 18164 23630 18216
rect 25317 18207 25375 18213
rect 25317 18173 25329 18207
rect 25363 18204 25375 18207
rect 27062 18204 27068 18216
rect 25363 18176 27068 18204
rect 25363 18173 25375 18176
rect 25317 18167 25375 18173
rect 27062 18164 27068 18176
rect 27120 18164 27126 18216
rect 27249 18207 27307 18213
rect 27249 18173 27261 18207
rect 27295 18173 27307 18207
rect 27249 18167 27307 18173
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 20438 18068 20444 18080
rect 19484 18040 20444 18068
rect 19484 18028 19490 18040
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 25130 18028 25136 18080
rect 25188 18068 25194 18080
rect 26329 18071 26387 18077
rect 26329 18068 26341 18071
rect 25188 18040 26341 18068
rect 25188 18028 25194 18040
rect 26329 18037 26341 18040
rect 26375 18037 26387 18071
rect 27264 18068 27292 18167
rect 27522 18164 27528 18216
rect 27580 18204 27586 18216
rect 28368 18204 28396 18232
rect 27580 18176 27625 18204
rect 28368 18176 29592 18204
rect 27580 18164 27586 18176
rect 29564 18136 29592 18176
rect 29730 18164 29736 18216
rect 29788 18204 29794 18216
rect 30377 18207 30435 18213
rect 30377 18204 30389 18207
rect 29788 18176 30389 18204
rect 29788 18164 29794 18176
rect 30377 18173 30389 18176
rect 30423 18173 30435 18207
rect 30377 18167 30435 18173
rect 31110 18164 31116 18216
rect 31168 18204 31174 18216
rect 34256 18204 34284 18235
rect 31168 18176 34284 18204
rect 34900 18204 34928 18235
rect 35710 18232 35716 18284
rect 35768 18272 35774 18284
rect 36173 18275 36231 18281
rect 36173 18272 36185 18275
rect 35768 18244 36185 18272
rect 35768 18232 35774 18244
rect 36173 18241 36185 18244
rect 36219 18241 36231 18275
rect 37642 18272 37648 18284
rect 37603 18244 37648 18272
rect 36173 18235 36231 18241
rect 37642 18232 37648 18244
rect 37700 18232 37706 18284
rect 38105 18275 38163 18281
rect 38105 18241 38117 18275
rect 38151 18241 38163 18275
rect 38105 18235 38163 18241
rect 36354 18204 36360 18216
rect 34900 18176 36360 18204
rect 31168 18164 31174 18176
rect 33870 18136 33876 18148
rect 29564 18108 33876 18136
rect 33870 18096 33876 18108
rect 33928 18096 33934 18148
rect 31846 18068 31852 18080
rect 27264 18040 31852 18068
rect 26329 18031 26387 18037
rect 31846 18028 31852 18040
rect 31904 18028 31910 18080
rect 33045 18071 33103 18077
rect 33045 18037 33057 18071
rect 33091 18068 33103 18071
rect 33226 18068 33232 18080
rect 33091 18040 33232 18068
rect 33091 18037 33103 18040
rect 33045 18031 33103 18037
rect 33226 18028 33232 18040
rect 33284 18028 33290 18080
rect 34164 18068 34192 18176
rect 36354 18164 36360 18176
rect 36412 18164 36418 18216
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 38010 18204 38016 18216
rect 37516 18176 38016 18204
rect 37516 18164 37522 18176
rect 38010 18164 38016 18176
rect 38068 18204 38074 18216
rect 38120 18204 38148 18235
rect 38068 18176 38148 18204
rect 38068 18164 38074 18176
rect 34238 18096 34244 18148
rect 34296 18136 34302 18148
rect 38197 18139 38255 18145
rect 38197 18136 38209 18139
rect 34296 18108 38209 18136
rect 34296 18096 34302 18108
rect 38197 18105 38209 18108
rect 38243 18105 38255 18139
rect 38197 18099 38255 18105
rect 37458 18068 37464 18080
rect 34164 18040 37464 18068
rect 37458 18028 37464 18040
rect 37516 18028 37522 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4062 17864 4068 17876
rect 4023 17836 4068 17864
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 17773 17867 17831 17873
rect 17773 17864 17785 17867
rect 11112 17836 17785 17864
rect 11112 17824 11118 17836
rect 17773 17833 17785 17836
rect 17819 17833 17831 17867
rect 17773 17827 17831 17833
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18012 17836 26924 17864
rect 18012 17824 18018 17836
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 14274 17796 14280 17808
rect 1912 17768 14280 17796
rect 1912 17756 1918 17768
rect 14274 17756 14280 17768
rect 14332 17756 14338 17808
rect 18417 17799 18475 17805
rect 18417 17796 18429 17799
rect 14384 17768 18429 17796
rect 10226 17728 10232 17740
rect 10187 17700 10232 17728
rect 10226 17688 10232 17700
rect 10284 17728 10290 17740
rect 10594 17728 10600 17740
rect 10284 17700 10600 17728
rect 10284 17688 10290 17700
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 12066 17728 12072 17740
rect 12027 17700 12072 17728
rect 12066 17688 12072 17700
rect 12124 17728 12130 17740
rect 12250 17728 12256 17740
rect 12124 17700 12256 17728
rect 12124 17688 12130 17700
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 14384 17728 14412 17768
rect 18417 17765 18429 17768
rect 18463 17765 18475 17799
rect 26896 17796 26924 17836
rect 27062 17824 27068 17876
rect 27120 17864 27126 17876
rect 29825 17867 29883 17873
rect 27120 17836 29776 17864
rect 27120 17824 27126 17836
rect 29638 17796 29644 17808
rect 18417 17759 18475 17765
rect 20088 17768 26832 17796
rect 26896 17768 29644 17796
rect 19978 17728 19984 17740
rect 13596 17700 14412 17728
rect 18340 17700 19984 17728
rect 13596 17688 13602 17700
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 2004 17632 4261 17660
rect 2004 17620 2010 17632
rect 4249 17629 4261 17632
rect 4295 17660 4307 17663
rect 9122 17660 9128 17672
rect 4295 17632 9128 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 17678 17660 17684 17672
rect 17639 17632 17684 17660
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 18340 17669 18368 17700
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 18325 17623 18383 17629
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 20088 17669 20116 17768
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 22830 17728 22836 17740
rect 20947 17700 22836 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 22922 17688 22928 17740
rect 22980 17728 22986 17740
rect 25038 17728 25044 17740
rect 22980 17700 25044 17728
rect 22980 17688 22986 17700
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 26804 17728 26832 17768
rect 29638 17756 29644 17768
rect 29696 17756 29702 17808
rect 29748 17796 29776 17836
rect 29825 17833 29837 17867
rect 29871 17864 29883 17867
rect 30006 17864 30012 17876
rect 29871 17836 30012 17864
rect 29871 17833 29883 17836
rect 29825 17827 29883 17833
rect 30006 17824 30012 17836
rect 30064 17824 30070 17876
rect 30190 17824 30196 17876
rect 30248 17864 30254 17876
rect 35621 17867 35679 17873
rect 35621 17864 35633 17867
rect 30248 17836 35633 17864
rect 30248 17824 30254 17836
rect 35621 17833 35633 17836
rect 35667 17833 35679 17867
rect 35621 17827 35679 17833
rect 36909 17867 36967 17873
rect 36909 17833 36921 17867
rect 36955 17864 36967 17867
rect 37366 17864 37372 17876
rect 36955 17836 37372 17864
rect 36955 17833 36967 17836
rect 36909 17827 36967 17833
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 37553 17867 37611 17873
rect 37553 17833 37565 17867
rect 37599 17864 37611 17867
rect 37734 17864 37740 17876
rect 37599 17836 37740 17864
rect 37599 17833 37611 17836
rect 37553 17827 37611 17833
rect 37734 17824 37740 17836
rect 37792 17824 37798 17876
rect 29748 17768 30328 17796
rect 27154 17728 27160 17740
rect 26804 17700 27160 17728
rect 27154 17688 27160 17700
rect 27212 17688 27218 17740
rect 27433 17731 27491 17737
rect 27433 17697 27445 17731
rect 27479 17728 27491 17731
rect 29086 17728 29092 17740
rect 27479 17700 29092 17728
rect 27479 17697 27491 17700
rect 27433 17691 27491 17697
rect 29086 17688 29092 17700
rect 29144 17688 29150 17740
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17660 21603 17663
rect 22462 17660 22468 17672
rect 21591 17632 22468 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 22462 17620 22468 17632
rect 22520 17620 22526 17672
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 26697 17663 26755 17669
rect 26697 17660 26709 17663
rect 26660 17632 26709 17660
rect 26660 17620 26666 17632
rect 26697 17629 26709 17632
rect 26743 17629 26755 17663
rect 26697 17623 26755 17629
rect 28074 17620 28080 17672
rect 28132 17660 28138 17672
rect 28534 17660 28540 17672
rect 28132 17632 28177 17660
rect 28495 17632 28540 17660
rect 28132 17620 28138 17632
rect 28534 17620 28540 17632
rect 28592 17660 28598 17672
rect 29178 17660 29184 17672
rect 28592 17632 29184 17660
rect 28592 17620 28598 17632
rect 29178 17620 29184 17632
rect 29236 17620 29242 17672
rect 29454 17620 29460 17672
rect 29512 17660 29518 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29512 17632 29745 17660
rect 29512 17620 29518 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 30300 17660 30328 17768
rect 30374 17756 30380 17808
rect 30432 17796 30438 17808
rect 30469 17799 30527 17805
rect 30469 17796 30481 17799
rect 30432 17768 30481 17796
rect 30432 17756 30438 17768
rect 30469 17765 30481 17768
rect 30515 17765 30527 17799
rect 34977 17799 35035 17805
rect 30469 17759 30527 17765
rect 31726 17768 34928 17796
rect 31573 17731 31631 17737
rect 31573 17697 31585 17731
rect 31619 17728 31631 17731
rect 31726 17728 31754 17768
rect 31938 17728 31944 17740
rect 31619 17700 31754 17728
rect 31899 17700 31944 17728
rect 31619 17697 31631 17700
rect 31573 17691 31631 17697
rect 31938 17688 31944 17700
rect 31996 17728 32002 17740
rect 32122 17728 32128 17740
rect 31996 17700 32128 17728
rect 31996 17688 32002 17700
rect 32122 17688 32128 17700
rect 32180 17688 32186 17740
rect 33962 17728 33968 17740
rect 33923 17700 33968 17728
rect 33962 17688 33968 17700
rect 34020 17688 34026 17740
rect 34514 17688 34520 17740
rect 34572 17728 34578 17740
rect 34698 17728 34704 17740
rect 34572 17700 34704 17728
rect 34572 17688 34578 17700
rect 34698 17688 34704 17700
rect 34756 17688 34762 17740
rect 34900 17728 34928 17768
rect 34977 17765 34989 17799
rect 35023 17796 35035 17799
rect 37642 17796 37648 17808
rect 35023 17768 37648 17796
rect 35023 17765 35035 17768
rect 34977 17759 35035 17765
rect 37642 17756 37648 17768
rect 37700 17756 37706 17808
rect 35710 17728 35716 17740
rect 34900 17700 35716 17728
rect 35710 17688 35716 17700
rect 35768 17688 35774 17740
rect 37182 17688 37188 17740
rect 37240 17728 37246 17740
rect 38197 17731 38255 17737
rect 38197 17728 38209 17731
rect 37240 17700 38209 17728
rect 37240 17688 37246 17700
rect 38197 17697 38209 17700
rect 38243 17697 38255 17731
rect 38197 17691 38255 17697
rect 30374 17660 30380 17672
rect 30287 17632 30380 17660
rect 29733 17623 29791 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 34885 17663 34943 17669
rect 34885 17629 34897 17663
rect 34931 17660 34943 17663
rect 35342 17660 35348 17672
rect 34931 17632 35348 17660
rect 34931 17629 34943 17632
rect 34885 17623 34943 17629
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 35529 17663 35587 17669
rect 35529 17629 35541 17663
rect 35575 17629 35587 17663
rect 36170 17660 36176 17672
rect 36131 17632 36176 17660
rect 35529 17623 35587 17629
rect 9950 17592 9956 17604
rect 9911 17564 9956 17592
rect 9950 17552 9956 17564
rect 10008 17552 10014 17604
rect 10045 17595 10103 17601
rect 10045 17561 10057 17595
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 10060 17524 10088 17555
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 11020 17564 12112 17592
rect 11020 17552 11026 17564
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10060 17496 11069 17524
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 12084 17524 12112 17564
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 12713 17595 12771 17601
rect 12216 17564 12261 17592
rect 12216 17552 12222 17564
rect 12713 17561 12725 17595
rect 12759 17592 12771 17595
rect 13446 17592 13452 17604
rect 12759 17564 13452 17592
rect 12759 17561 12771 17564
rect 12713 17555 12771 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 19521 17595 19579 17601
rect 16540 17564 18552 17592
rect 16540 17552 16546 17564
rect 17954 17524 17960 17536
rect 12084 17496 17960 17524
rect 11057 17487 11115 17493
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18524 17524 18552 17564
rect 19521 17561 19533 17595
rect 19567 17592 19579 17595
rect 20714 17592 20720 17604
rect 19567 17564 20720 17592
rect 19567 17561 19579 17564
rect 19521 17555 19579 17561
rect 20714 17552 20720 17564
rect 20772 17552 20778 17604
rect 20993 17595 21051 17601
rect 20993 17561 21005 17595
rect 21039 17592 21051 17595
rect 21358 17592 21364 17604
rect 21039 17564 21364 17592
rect 21039 17561 21051 17564
rect 20993 17555 21051 17561
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22649 17595 22707 17601
rect 22649 17592 22661 17595
rect 21692 17564 22661 17592
rect 21692 17552 21698 17564
rect 22649 17561 22661 17564
rect 22695 17561 22707 17595
rect 22649 17555 22707 17561
rect 22738 17552 22744 17604
rect 22796 17592 22802 17604
rect 22796 17564 22841 17592
rect 22796 17552 22802 17564
rect 26970 17552 26976 17604
rect 27028 17592 27034 17604
rect 27502 17595 27560 17601
rect 27502 17592 27514 17595
rect 27028 17564 27514 17592
rect 27028 17552 27034 17564
rect 27502 17561 27514 17564
rect 27548 17561 27560 17595
rect 28626 17592 28632 17604
rect 28587 17564 28632 17592
rect 27502 17555 27560 17561
rect 28626 17552 28632 17564
rect 28684 17552 28690 17604
rect 31665 17595 31723 17601
rect 31665 17561 31677 17595
rect 31711 17561 31723 17595
rect 31665 17555 31723 17561
rect 33137 17595 33195 17601
rect 33137 17561 33149 17595
rect 33183 17561 33195 17595
rect 33137 17555 33195 17561
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 18524 17496 20177 17524
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20165 17487 20223 17493
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 25314 17524 25320 17536
rect 22612 17496 25320 17524
rect 22612 17484 22618 17496
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 26789 17527 26847 17533
rect 26789 17493 26801 17527
rect 26835 17524 26847 17527
rect 31680 17524 31708 17555
rect 26835 17496 31708 17524
rect 33152 17524 33180 17555
rect 33226 17552 33232 17604
rect 33284 17592 33290 17604
rect 33284 17564 33329 17592
rect 33284 17552 33290 17564
rect 33778 17552 33784 17604
rect 33836 17592 33842 17604
rect 34330 17592 34336 17604
rect 33836 17564 34336 17592
rect 33836 17552 33842 17564
rect 34330 17552 34336 17564
rect 34388 17552 34394 17604
rect 35544 17592 35572 17623
rect 36170 17620 36176 17632
rect 36228 17620 36234 17672
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17660 36875 17663
rect 37274 17660 37280 17672
rect 36863 17632 37280 17660
rect 36863 17629 36875 17632
rect 36817 17623 36875 17629
rect 37274 17620 37280 17632
rect 37332 17620 37338 17672
rect 37458 17660 37464 17672
rect 37419 17632 37464 17660
rect 37458 17620 37464 17632
rect 37516 17660 37522 17672
rect 38105 17663 38163 17669
rect 38105 17660 38117 17663
rect 37516 17632 38117 17660
rect 37516 17620 37522 17632
rect 38105 17629 38117 17632
rect 38151 17629 38163 17663
rect 38105 17623 38163 17629
rect 37826 17592 37832 17604
rect 35544 17564 37832 17592
rect 37826 17552 37832 17564
rect 37884 17552 37890 17604
rect 35986 17524 35992 17536
rect 33152 17496 35992 17524
rect 26835 17493 26847 17496
rect 26789 17487 26847 17493
rect 35986 17484 35992 17496
rect 36044 17484 36050 17536
rect 36262 17524 36268 17536
rect 36223 17496 36268 17524
rect 36262 17484 36268 17496
rect 36320 17484 36326 17536
rect 36446 17484 36452 17536
rect 36504 17524 36510 17536
rect 36630 17524 36636 17536
rect 36504 17496 36636 17524
rect 36504 17484 36510 17496
rect 36630 17484 36636 17496
rect 36688 17484 36694 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 11238 17280 11244 17332
rect 11296 17320 11302 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 11296 17292 13093 17320
rect 11296 17280 11302 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13081 17283 13139 17289
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 17497 17323 17555 17329
rect 17497 17320 17509 17323
rect 14240 17292 17509 17320
rect 14240 17280 14246 17292
rect 17497 17289 17509 17292
rect 17543 17289 17555 17323
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 17497 17283 17555 17289
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 25038 17280 25044 17332
rect 25096 17320 25102 17332
rect 27062 17320 27068 17332
rect 25096 17292 27068 17320
rect 25096 17280 25102 17292
rect 27062 17280 27068 17292
rect 27120 17280 27126 17332
rect 27246 17320 27252 17332
rect 27207 17292 27252 17320
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 28442 17320 28448 17332
rect 28184 17292 28448 17320
rect 9217 17255 9275 17261
rect 9217 17221 9229 17255
rect 9263 17252 9275 17255
rect 9950 17252 9956 17264
rect 9263 17224 9956 17252
rect 9263 17221 9275 17224
rect 9217 17215 9275 17221
rect 9950 17212 9956 17224
rect 10008 17252 10014 17264
rect 10137 17255 10195 17261
rect 10137 17252 10149 17255
rect 10008 17224 10149 17252
rect 10008 17212 10014 17224
rect 10137 17221 10149 17224
rect 10183 17221 10195 17255
rect 10137 17215 10195 17221
rect 10229 17255 10287 17261
rect 10229 17221 10241 17255
rect 10275 17252 10287 17255
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 10275 17224 14289 17252
rect 10275 17221 10287 17224
rect 10229 17215 10287 17221
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 17678 17212 17684 17264
rect 17736 17252 17742 17264
rect 17736 17224 22416 17252
rect 17736 17212 17742 17224
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12584 17156 12633 17184
rect 12584 17144 12590 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 12621 17147 12679 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 17405 17187 17463 17193
rect 17405 17153 17417 17187
rect 17451 17184 17463 17187
rect 17954 17184 17960 17196
rect 17451 17156 17960 17184
rect 17451 17153 17463 17156
rect 17405 17147 17463 17153
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 10962 17116 10968 17128
rect 10923 17088 10968 17116
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 14200 17048 14228 17147
rect 17954 17144 17960 17156
rect 18012 17184 18018 17196
rect 18230 17184 18236 17196
rect 18012 17156 18236 17184
rect 18012 17144 18018 17156
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20806 17184 20812 17196
rect 20119 17156 20812 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 21048 17156 21281 17184
rect 21048 17144 21054 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 22278 17184 22284 17196
rect 22239 17156 22284 17184
rect 21269 17147 21327 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 22388 17184 22416 17224
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 28184 17252 28212 17292
rect 28442 17280 28448 17292
rect 28500 17280 28506 17332
rect 30837 17323 30895 17329
rect 30837 17320 30849 17323
rect 29380 17292 30849 17320
rect 22520 17224 28212 17252
rect 28261 17255 28319 17261
rect 22520 17212 22526 17224
rect 28261 17221 28273 17255
rect 28307 17252 28319 17255
rect 29178 17252 29184 17264
rect 28307 17224 29184 17252
rect 28307 17221 28319 17224
rect 28261 17215 28319 17221
rect 29178 17212 29184 17224
rect 29236 17212 29242 17264
rect 29380 17261 29408 17292
rect 30837 17289 30849 17292
rect 30883 17289 30895 17323
rect 33962 17320 33968 17332
rect 30837 17283 30895 17289
rect 30944 17292 33968 17320
rect 29365 17255 29423 17261
rect 29365 17221 29377 17255
rect 29411 17221 29423 17255
rect 29365 17215 29423 17221
rect 29454 17212 29460 17264
rect 29512 17252 29518 17264
rect 29512 17224 29557 17252
rect 29512 17212 29518 17224
rect 29638 17212 29644 17264
rect 29696 17252 29702 17264
rect 30944 17252 30972 17292
rect 33962 17280 33968 17292
rect 34020 17280 34026 17332
rect 29696 17224 30972 17252
rect 31573 17255 31631 17261
rect 29696 17212 29702 17224
rect 31573 17221 31585 17255
rect 31619 17252 31631 17255
rect 32677 17255 32735 17261
rect 32677 17252 32689 17255
rect 31619 17224 32689 17252
rect 31619 17221 31631 17224
rect 31573 17215 31631 17221
rect 32677 17221 32689 17224
rect 32723 17221 32735 17255
rect 34146 17252 34152 17264
rect 32677 17215 32735 17221
rect 33980 17224 34152 17252
rect 25222 17184 25228 17196
rect 22388 17156 25228 17184
rect 25222 17144 25228 17156
rect 25280 17144 25286 17196
rect 25406 17184 25412 17196
rect 25367 17156 25412 17184
rect 25406 17144 25412 17156
rect 25464 17144 25470 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27430 17184 27436 17196
rect 27203 17156 27436 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 30282 17144 30288 17196
rect 30340 17184 30346 17196
rect 31481 17187 31539 17193
rect 31481 17184 31493 17187
rect 30340 17156 31493 17184
rect 30340 17144 30346 17156
rect 31481 17153 31493 17156
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 23293 17119 23351 17125
rect 23293 17116 23305 17119
rect 17828 17088 23305 17116
rect 17828 17076 17834 17088
rect 23293 17085 23305 17088
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17085 23535 17119
rect 23477 17079 23535 17085
rect 14200 17020 18184 17048
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12986 16980 12992 16992
rect 12483 16952 12992 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 18156 16980 18184 17020
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 21634 17048 21640 17060
rect 20220 17020 21640 17048
rect 20220 17008 20226 17020
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 22097 17051 22155 17057
rect 22097 17017 22109 17051
rect 22143 17048 22155 17051
rect 23492 17048 23520 17079
rect 27982 17076 27988 17128
rect 28040 17116 28046 17128
rect 28169 17119 28227 17125
rect 28169 17116 28181 17119
rect 28040 17088 28181 17116
rect 28040 17076 28046 17088
rect 28169 17085 28181 17088
rect 28215 17085 28227 17119
rect 28442 17116 28448 17128
rect 28403 17088 28448 17116
rect 28169 17079 28227 17085
rect 22143 17020 23520 17048
rect 23937 17051 23995 17057
rect 22143 17017 22155 17020
rect 22097 17011 22155 17017
rect 23937 17017 23949 17051
rect 23983 17048 23995 17051
rect 27246 17048 27252 17060
rect 23983 17020 27252 17048
rect 23983 17017 23995 17020
rect 23937 17011 23995 17017
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 25406 16980 25412 16992
rect 18156 16952 25412 16980
rect 25406 16940 25412 16952
rect 25464 16940 25470 16992
rect 25501 16983 25559 16989
rect 25501 16949 25513 16983
rect 25547 16980 25559 16983
rect 25590 16980 25596 16992
rect 25547 16952 25596 16980
rect 25547 16949 25559 16952
rect 25501 16943 25559 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 28184 16980 28212 17079
rect 28442 17076 28448 17088
rect 28500 17076 28506 17128
rect 28534 17076 28540 17128
rect 28592 17116 28598 17128
rect 29641 17119 29699 17125
rect 29641 17116 29653 17119
rect 28592 17088 29653 17116
rect 28592 17076 28598 17088
rect 29641 17085 29653 17088
rect 29687 17085 29699 17119
rect 29641 17079 29699 17085
rect 31846 17076 31852 17128
rect 31904 17116 31910 17128
rect 32585 17119 32643 17125
rect 32585 17116 32597 17119
rect 31904 17088 32597 17116
rect 31904 17076 31910 17088
rect 32585 17085 32597 17088
rect 32631 17085 32643 17119
rect 32585 17079 32643 17085
rect 32861 17119 32919 17125
rect 32861 17085 32873 17119
rect 32907 17085 32919 17119
rect 32861 17079 32919 17085
rect 28460 17048 28488 17076
rect 30742 17048 30748 17060
rect 28460 17020 30748 17048
rect 30742 17008 30748 17020
rect 30800 17048 30806 17060
rect 30926 17048 30932 17060
rect 30800 17020 30932 17048
rect 30800 17008 30806 17020
rect 30926 17008 30932 17020
rect 30984 17008 30990 17060
rect 31938 17008 31944 17060
rect 31996 17048 32002 17060
rect 32876 17048 32904 17079
rect 33980 17060 34008 17224
rect 34146 17212 34152 17224
rect 34204 17212 34210 17264
rect 34241 17255 34299 17261
rect 34241 17221 34253 17255
rect 34287 17252 34299 17255
rect 34790 17252 34796 17264
rect 34287 17224 34796 17252
rect 34287 17221 34299 17224
rect 34241 17215 34299 17221
rect 34790 17212 34796 17224
rect 34848 17212 34854 17264
rect 35342 17212 35348 17264
rect 35400 17252 35406 17264
rect 35805 17255 35863 17261
rect 35805 17252 35817 17255
rect 35400 17224 35817 17252
rect 35400 17212 35406 17224
rect 35805 17221 35817 17224
rect 35851 17221 35863 17255
rect 35805 17215 35863 17221
rect 37366 17212 37372 17264
rect 37424 17252 37430 17264
rect 37645 17255 37703 17261
rect 37645 17252 37657 17255
rect 37424 17224 37657 17252
rect 37424 17212 37430 17224
rect 37645 17221 37657 17224
rect 37691 17221 37703 17255
rect 37645 17215 37703 17221
rect 38470 17212 38476 17264
rect 38528 17252 38534 17264
rect 38838 17252 38844 17264
rect 38528 17224 38844 17252
rect 38528 17212 38534 17224
rect 38838 17212 38844 17224
rect 38896 17212 38902 17264
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 34425 17119 34483 17125
rect 34425 17085 34437 17119
rect 34471 17085 34483 17119
rect 35710 17116 35716 17128
rect 35671 17088 35716 17116
rect 34425 17079 34483 17085
rect 31996 17020 32904 17048
rect 31996 17008 32002 17020
rect 33962 17008 33968 17060
rect 34020 17048 34026 17060
rect 34440 17048 34468 17079
rect 35710 17076 35716 17088
rect 35768 17076 35774 17128
rect 35894 17076 35900 17128
rect 35952 17116 35958 17128
rect 35989 17119 36047 17125
rect 35989 17116 36001 17119
rect 35952 17088 36001 17116
rect 35952 17076 35958 17088
rect 35989 17085 36001 17088
rect 36035 17085 36047 17119
rect 37550 17116 37556 17128
rect 37511 17088 37556 17116
rect 35989 17079 36047 17085
rect 37550 17076 37556 17088
rect 37608 17076 37614 17128
rect 38197 17119 38255 17125
rect 38197 17085 38209 17119
rect 38243 17116 38255 17119
rect 38286 17116 38292 17128
rect 38243 17088 38292 17116
rect 38243 17085 38255 17088
rect 38197 17079 38255 17085
rect 38286 17076 38292 17088
rect 38344 17076 38350 17128
rect 34020 17020 34468 17048
rect 34020 17008 34026 17020
rect 36262 16980 36268 16992
rect 28184 16952 36268 16980
rect 36262 16940 36268 16952
rect 36320 16940 36326 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 17034 16776 17040 16788
rect 12860 16748 17040 16776
rect 12860 16736 12866 16748
rect 17034 16736 17040 16748
rect 17092 16776 17098 16788
rect 17586 16776 17592 16788
rect 17092 16748 17592 16776
rect 17092 16736 17098 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 22373 16779 22431 16785
rect 22373 16745 22385 16779
rect 22419 16776 22431 16779
rect 22738 16776 22744 16788
rect 22419 16748 22744 16776
rect 22419 16745 22431 16748
rect 22373 16739 22431 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27065 16779 27123 16785
rect 27065 16776 27077 16779
rect 27028 16748 27077 16776
rect 27028 16736 27034 16748
rect 27065 16745 27077 16748
rect 27111 16745 27123 16779
rect 27065 16739 27123 16745
rect 29178 16736 29184 16788
rect 29236 16776 29242 16788
rect 29825 16779 29883 16785
rect 29825 16776 29837 16779
rect 29236 16748 29837 16776
rect 29236 16736 29242 16748
rect 29825 16745 29837 16748
rect 29871 16745 29883 16779
rect 35526 16776 35532 16788
rect 29825 16739 29883 16745
rect 29932 16748 35532 16776
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 13320 16680 17448 16708
rect 13320 16668 13326 16680
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 15933 16643 15991 16649
rect 1636 16612 10180 16640
rect 1636 16600 1642 16612
rect 10152 16581 10180 16612
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16850 16640 16856 16652
rect 15979 16612 16856 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17034 16640 17040 16652
rect 16991 16612 17040 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17420 16640 17448 16680
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 20806 16708 20812 16720
rect 19024 16680 19932 16708
rect 20767 16680 20812 16708
rect 19024 16668 19030 16680
rect 19058 16640 19064 16652
rect 17420 16612 19064 16640
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16574 10195 16575
rect 10183 16546 10217 16574
rect 12618 16572 12624 16584
rect 10183 16541 10195 16546
rect 12579 16544 12624 16572
rect 10137 16535 10195 16541
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14918 16572 14924 16584
rect 14056 16544 14924 16572
rect 14056 16532 14062 16544
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 17420 16581 17448 16612
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19904 16581 19932 16680
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 20916 16680 23060 16708
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20916 16640 20944 16680
rect 23032 16649 23060 16680
rect 26142 16668 26148 16720
rect 26200 16708 26206 16720
rect 28629 16711 28687 16717
rect 28629 16708 28641 16711
rect 26200 16680 28641 16708
rect 26200 16668 26206 16680
rect 28629 16677 28641 16680
rect 28675 16677 28687 16711
rect 29932 16708 29960 16748
rect 35526 16736 35532 16748
rect 35584 16736 35590 16788
rect 28629 16671 28687 16677
rect 29748 16680 29960 16708
rect 20036 16612 20944 16640
rect 23017 16643 23075 16649
rect 20036 16600 20042 16612
rect 23017 16609 23029 16643
rect 23063 16609 23075 16643
rect 25498 16640 25504 16652
rect 25459 16612 25504 16640
rect 23017 16603 23075 16609
rect 25498 16600 25504 16612
rect 25556 16600 25562 16652
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 26844 16612 27016 16640
rect 26844 16600 26850 16612
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 21542 16572 21548 16584
rect 21503 16544 21548 16572
rect 19889 16535 19947 16541
rect 21542 16532 21548 16544
rect 21600 16532 21606 16584
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22554 16572 22560 16584
rect 22327 16544 22560 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 26988 16581 27016 16612
rect 27154 16600 27160 16652
rect 27212 16640 27218 16652
rect 29748 16640 29776 16680
rect 30374 16668 30380 16720
rect 30432 16708 30438 16720
rect 35158 16708 35164 16720
rect 30432 16680 35164 16708
rect 30432 16668 30438 16680
rect 35158 16668 35164 16680
rect 35216 16668 35222 16720
rect 35894 16668 35900 16720
rect 35952 16708 35958 16720
rect 35952 16680 36400 16708
rect 35952 16668 35958 16680
rect 27212 16612 29776 16640
rect 27212 16600 27218 16612
rect 29748 16581 29776 16612
rect 30098 16600 30104 16652
rect 30156 16640 30162 16652
rect 31754 16640 31760 16652
rect 30156 16612 30420 16640
rect 30156 16600 30162 16612
rect 30392 16581 30420 16612
rect 31680 16612 31760 16640
rect 26973 16575 27031 16581
rect 26973 16541 26985 16575
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 30377 16575 30435 16581
rect 30377 16541 30389 16575
rect 30423 16541 30435 16575
rect 30377 16535 30435 16541
rect 30466 16532 30472 16584
rect 30524 16572 30530 16584
rect 31018 16572 31024 16584
rect 30524 16544 30569 16572
rect 30979 16544 31024 16572
rect 30524 16532 30530 16544
rect 31018 16532 31024 16544
rect 31076 16532 31082 16584
rect 31110 16532 31116 16584
rect 31168 16572 31174 16584
rect 31680 16581 31708 16612
rect 31754 16600 31760 16612
rect 31812 16640 31818 16652
rect 32674 16640 32680 16652
rect 31812 16612 32680 16640
rect 31812 16600 31818 16612
rect 32324 16581 32352 16612
rect 32674 16600 32680 16612
rect 32732 16600 32738 16652
rect 33042 16600 33048 16652
rect 33100 16640 33106 16652
rect 35805 16643 35863 16649
rect 33100 16612 34928 16640
rect 33100 16600 33106 16612
rect 31665 16575 31723 16581
rect 31168 16544 31213 16572
rect 31168 16532 31174 16544
rect 31665 16541 31677 16575
rect 31711 16541 31723 16575
rect 31665 16535 31723 16541
rect 32309 16575 32367 16581
rect 32309 16541 32321 16575
rect 32355 16541 32367 16575
rect 32309 16535 32367 16541
rect 32398 16532 32404 16584
rect 32456 16572 32462 16584
rect 32766 16572 32772 16584
rect 32456 16544 32772 16572
rect 32456 16532 32462 16544
rect 32766 16532 32772 16544
rect 32824 16572 32830 16584
rect 32953 16575 33011 16581
rect 32953 16572 32965 16575
rect 32824 16544 32965 16572
rect 32824 16532 32830 16544
rect 32953 16541 32965 16544
rect 32999 16541 33011 16575
rect 32953 16535 33011 16541
rect 33502 16532 33508 16584
rect 33560 16572 33566 16584
rect 34900 16581 34928 16612
rect 35805 16609 35817 16643
rect 35851 16640 35863 16643
rect 36262 16640 36268 16652
rect 35851 16612 36268 16640
rect 35851 16609 35863 16612
rect 35805 16603 35863 16609
rect 36262 16600 36268 16612
rect 36320 16600 36326 16652
rect 36372 16649 36400 16680
rect 36357 16643 36415 16649
rect 36357 16609 36369 16643
rect 36403 16609 36415 16643
rect 37458 16640 37464 16652
rect 36357 16603 36415 16609
rect 37384 16612 37464 16640
rect 37384 16581 37412 16612
rect 37458 16600 37464 16612
rect 37516 16640 37522 16652
rect 37516 16612 38056 16640
rect 37516 16600 37522 16612
rect 38028 16581 38056 16612
rect 33597 16575 33655 16581
rect 33597 16572 33609 16575
rect 33560 16544 33609 16572
rect 33560 16532 33566 16544
rect 33597 16541 33609 16544
rect 33643 16541 33655 16575
rect 33597 16535 33655 16541
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 37369 16575 37427 16581
rect 37369 16541 37381 16575
rect 37415 16541 37427 16575
rect 37369 16535 37427 16541
rect 38013 16575 38071 16581
rect 38013 16541 38025 16575
rect 38059 16541 38071 16575
rect 38013 16535 38071 16541
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 10229 16507 10287 16513
rect 10229 16504 10241 16507
rect 10100 16476 10241 16504
rect 10100 16464 10106 16476
rect 10229 16473 10241 16476
rect 10275 16473 10287 16507
rect 10229 16467 10287 16473
rect 16025 16507 16083 16513
rect 16025 16473 16037 16507
rect 16071 16504 16083 16507
rect 16758 16504 16764 16516
rect 16071 16476 16764 16504
rect 16071 16473 16083 16476
rect 16025 16467 16083 16473
rect 16758 16464 16764 16476
rect 16816 16464 16822 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 19981 16507 20039 16513
rect 19981 16504 19993 16507
rect 17000 16476 19993 16504
rect 17000 16464 17006 16476
rect 19981 16473 19993 16476
rect 20027 16473 20039 16507
rect 19981 16467 20039 16473
rect 20530 16464 20536 16516
rect 20588 16504 20594 16516
rect 20625 16507 20683 16513
rect 20625 16504 20637 16507
rect 20588 16476 20637 16504
rect 20588 16464 20594 16476
rect 20625 16473 20637 16476
rect 20671 16473 20683 16507
rect 20625 16467 20683 16473
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 23109 16507 23167 16513
rect 20772 16476 22600 16504
rect 20772 16464 20778 16476
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 12437 16439 12495 16445
rect 12437 16436 12449 16439
rect 10836 16408 12449 16436
rect 10836 16396 10842 16408
rect 12437 16405 12449 16408
rect 12483 16405 12495 16439
rect 12437 16399 12495 16405
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 17092 16408 17509 16436
rect 17092 16396 17098 16408
rect 17497 16405 17509 16408
rect 17543 16405 17555 16439
rect 17497 16399 17555 16405
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 20070 16436 20076 16448
rect 19484 16408 20076 16436
rect 19484 16396 19490 16408
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 21361 16439 21419 16445
rect 21361 16405 21373 16439
rect 21407 16436 21419 16439
rect 22278 16436 22284 16448
rect 21407 16408 22284 16436
rect 21407 16405 21419 16408
rect 21361 16399 21419 16405
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 22572 16436 22600 16476
rect 23109 16473 23121 16507
rect 23155 16473 23167 16507
rect 23109 16467 23167 16473
rect 24029 16507 24087 16513
rect 24029 16473 24041 16507
rect 24075 16473 24087 16507
rect 24029 16467 24087 16473
rect 23124 16436 23152 16467
rect 22572 16408 23152 16436
rect 24044 16436 24072 16467
rect 25590 16464 25596 16516
rect 25648 16504 25654 16516
rect 26510 16504 26516 16516
rect 25648 16476 25693 16504
rect 26423 16476 26516 16504
rect 25648 16464 25654 16476
rect 26510 16464 26516 16476
rect 26568 16504 26574 16516
rect 28074 16504 28080 16516
rect 26568 16476 27752 16504
rect 28035 16476 28080 16504
rect 26568 16464 26574 16476
rect 27614 16436 27620 16448
rect 24044 16408 27620 16436
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 27724 16436 27752 16476
rect 28074 16464 28080 16476
rect 28132 16464 28138 16516
rect 28166 16464 28172 16516
rect 28224 16504 28230 16516
rect 28224 16476 28269 16504
rect 28224 16464 28230 16476
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 30190 16504 30196 16516
rect 29328 16476 30196 16504
rect 29328 16464 29334 16476
rect 30190 16464 30196 16476
rect 30248 16464 30254 16516
rect 31294 16464 31300 16516
rect 31352 16504 31358 16516
rect 33045 16507 33103 16513
rect 33045 16504 33057 16507
rect 31352 16476 33057 16504
rect 31352 16464 31358 16476
rect 33045 16473 33057 16476
rect 33091 16473 33103 16507
rect 33045 16467 33103 16473
rect 35894 16464 35900 16516
rect 35952 16504 35958 16516
rect 35952 16476 35997 16504
rect 35952 16464 35958 16476
rect 37918 16464 37924 16516
rect 37976 16504 37982 16516
rect 38105 16507 38163 16513
rect 38105 16504 38117 16507
rect 37976 16476 38117 16504
rect 37976 16464 37982 16476
rect 38105 16473 38117 16476
rect 38151 16473 38163 16507
rect 38105 16467 38163 16473
rect 29914 16436 29920 16448
rect 27724 16408 29920 16436
rect 29914 16396 29920 16408
rect 29972 16396 29978 16448
rect 31754 16436 31760 16448
rect 31715 16408 31760 16436
rect 31754 16396 31760 16408
rect 31812 16396 31818 16448
rect 32401 16439 32459 16445
rect 32401 16405 32413 16439
rect 32447 16436 32459 16439
rect 32490 16436 32496 16448
rect 32447 16408 32496 16436
rect 32447 16405 32459 16408
rect 32401 16399 32459 16405
rect 32490 16396 32496 16408
rect 32548 16396 32554 16448
rect 33686 16436 33692 16448
rect 33647 16408 33692 16436
rect 33686 16396 33692 16408
rect 33744 16396 33750 16448
rect 34974 16436 34980 16448
rect 34935 16408 34980 16436
rect 34974 16396 34980 16408
rect 35032 16396 35038 16448
rect 37461 16439 37519 16445
rect 37461 16405 37473 16439
rect 37507 16436 37519 16439
rect 39482 16436 39488 16448
rect 37507 16408 39488 16436
rect 37507 16405 37519 16408
rect 37461 16399 37519 16405
rect 39482 16396 39488 16408
rect 39540 16396 39546 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11974 16232 11980 16244
rect 11011 16204 11980 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 14108 16204 14688 16232
rect 12529 16167 12587 16173
rect 12529 16133 12541 16167
rect 12575 16164 12587 16167
rect 12710 16164 12716 16176
rect 12575 16136 12716 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 13449 16167 13507 16173
rect 13449 16133 13461 16167
rect 13495 16164 13507 16167
rect 13998 16164 14004 16176
rect 13495 16136 14004 16164
rect 13495 16133 13507 16136
rect 13449 16127 13507 16133
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 10778 16096 10784 16108
rect 1627 16068 10784 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 10226 16028 10232 16040
rect 10187 16000 10232 16028
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 10888 15960 10916 16059
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11480 16000 12449 16028
rect 11480 15988 11486 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 14108 16028 14136 16204
rect 14366 16164 14372 16176
rect 14327 16136 14372 16164
rect 14366 16124 14372 16136
rect 14424 16124 14430 16176
rect 14660 16164 14688 16204
rect 14734 16192 14740 16244
rect 14792 16232 14798 16244
rect 19521 16235 19579 16241
rect 14792 16204 17172 16232
rect 14792 16192 14798 16204
rect 16298 16164 16304 16176
rect 14660 16136 16304 16164
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 17034 16164 17040 16176
rect 16995 16136 17040 16164
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17144 16164 17172 16204
rect 19521 16201 19533 16235
rect 19567 16232 19579 16235
rect 19978 16232 19984 16244
rect 19567 16204 19984 16232
rect 19567 16201 19579 16204
rect 19521 16195 19579 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 20088 16204 26556 16232
rect 20088 16164 20116 16204
rect 17144 16136 20116 16164
rect 22646 16124 22652 16176
rect 22704 16164 22710 16176
rect 22741 16167 22799 16173
rect 22741 16164 22753 16167
rect 22704 16136 22753 16164
rect 22704 16124 22710 16136
rect 22741 16133 22753 16136
rect 22787 16133 22799 16167
rect 26528 16164 26556 16204
rect 28166 16192 28172 16244
rect 28224 16232 28230 16244
rect 28997 16235 29055 16241
rect 28997 16232 29009 16235
rect 28224 16204 29009 16232
rect 28224 16192 28230 16204
rect 28997 16201 29009 16204
rect 29043 16201 29055 16235
rect 28997 16195 29055 16201
rect 29454 16192 29460 16244
rect 29512 16232 29518 16244
rect 29641 16235 29699 16241
rect 29641 16232 29653 16235
rect 29512 16204 29653 16232
rect 29512 16192 29518 16204
rect 29641 16201 29653 16204
rect 29687 16201 29699 16235
rect 29641 16195 29699 16201
rect 31478 16192 31484 16244
rect 31536 16232 31542 16244
rect 33686 16232 33692 16244
rect 31536 16204 33692 16232
rect 31536 16192 31542 16204
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 35250 16192 35256 16244
rect 35308 16232 35314 16244
rect 35805 16235 35863 16241
rect 35805 16232 35817 16235
rect 35308 16204 35817 16232
rect 35308 16192 35314 16204
rect 35805 16201 35817 16204
rect 35851 16201 35863 16235
rect 36446 16232 36452 16244
rect 36407 16204 36452 16232
rect 35805 16195 35863 16201
rect 36446 16192 36452 16204
rect 36504 16192 36510 16244
rect 26528 16136 31156 16164
rect 22741 16127 22799 16133
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 14108 16000 14289 16028
rect 12437 15991 12495 15997
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 14553 15991 14611 15997
rect 8536 15932 10916 15960
rect 8536 15920 8542 15932
rect 13722 15920 13728 15972
rect 13780 15960 13786 15972
rect 14568 15960 14596 15991
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 15997 17279 16031
rect 19444 16028 19472 16059
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 19852 16068 20269 16096
rect 19852 16056 19858 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 20346 16056 20352 16108
rect 20404 16096 20410 16108
rect 20714 16096 20720 16108
rect 20404 16068 20720 16096
rect 20404 16056 20410 16068
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 28258 16096 28264 16108
rect 28219 16068 28264 16096
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 28718 16056 28724 16108
rect 28776 16096 28782 16108
rect 28905 16099 28963 16105
rect 28905 16096 28917 16099
rect 28776 16068 28917 16096
rect 28776 16056 28782 16068
rect 28905 16065 28917 16068
rect 28951 16065 28963 16099
rect 29546 16096 29552 16108
rect 29507 16068 29552 16096
rect 28905 16059 28963 16065
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 30190 16096 30196 16108
rect 30151 16068 30196 16096
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 31128 16105 31156 16136
rect 32214 16124 32220 16176
rect 32272 16164 32278 16176
rect 32398 16164 32404 16176
rect 32272 16136 32404 16164
rect 32272 16124 32278 16136
rect 32398 16124 32404 16136
rect 32456 16124 32462 16176
rect 32493 16167 32551 16173
rect 32493 16133 32505 16167
rect 32539 16164 32551 16167
rect 33778 16164 33784 16176
rect 32539 16136 33784 16164
rect 32539 16133 32551 16136
rect 32493 16127 32551 16133
rect 33778 16124 33784 16136
rect 33836 16124 33842 16176
rect 34057 16167 34115 16173
rect 34057 16133 34069 16167
rect 34103 16164 34115 16167
rect 35161 16167 35219 16173
rect 35161 16164 35173 16167
rect 34103 16136 35173 16164
rect 34103 16133 34115 16136
rect 34057 16127 34115 16133
rect 35161 16133 35173 16136
rect 35207 16133 35219 16167
rect 37734 16164 37740 16176
rect 37695 16136 37740 16164
rect 35161 16127 35219 16133
rect 37734 16124 37740 16136
rect 37792 16124 37798 16176
rect 31113 16099 31171 16105
rect 31113 16065 31125 16099
rect 31159 16065 31171 16099
rect 31294 16096 31300 16108
rect 31255 16068 31300 16096
rect 31113 16059 31171 16065
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 35069 16099 35127 16105
rect 35069 16065 35081 16099
rect 35115 16096 35127 16099
rect 35526 16096 35532 16108
rect 35115 16068 35532 16096
rect 35115 16065 35127 16068
rect 35069 16059 35127 16065
rect 35526 16056 35532 16068
rect 35584 16056 35590 16108
rect 35713 16099 35771 16105
rect 35713 16065 35725 16099
rect 35759 16065 35771 16099
rect 35713 16059 35771 16065
rect 36357 16099 36415 16105
rect 36357 16065 36369 16099
rect 36403 16096 36415 16099
rect 36446 16096 36452 16108
rect 36403 16068 36452 16096
rect 36403 16065 36415 16068
rect 36357 16059 36415 16065
rect 20530 16028 20536 16040
rect 19444 16000 20536 16028
rect 17221 15991 17279 15997
rect 13780 15932 14596 15960
rect 13780 15920 13786 15932
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 17236 15892 17264 15991
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 22925 16031 22983 16037
rect 22925 16028 22937 16031
rect 22704 16000 22749 16028
rect 22848 16000 22937 16028
rect 22704 15988 22710 16000
rect 17310 15920 17316 15972
rect 17368 15960 17374 15972
rect 22848 15960 22876 16000
rect 22925 15997 22937 16000
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 31662 15988 31668 16040
rect 31720 16028 31726 16040
rect 32030 16028 32036 16040
rect 31720 16000 32036 16028
rect 31720 15988 31726 16000
rect 32030 15988 32036 16000
rect 32088 15988 32094 16040
rect 32398 16028 32404 16040
rect 32359 16000 32404 16028
rect 32398 15988 32404 16000
rect 32456 15988 32462 16040
rect 33318 16028 33324 16040
rect 33279 16000 33324 16028
rect 33318 15988 33324 16000
rect 33376 15988 33382 16040
rect 33686 15988 33692 16040
rect 33744 16028 33750 16040
rect 33965 16031 34023 16037
rect 33965 16028 33977 16031
rect 33744 16000 33977 16028
rect 33744 15988 33750 16000
rect 33965 15997 33977 16000
rect 34011 16028 34023 16031
rect 34146 16028 34152 16040
rect 34011 16000 34152 16028
rect 34011 15997 34023 16000
rect 33965 15991 34023 15997
rect 34146 15988 34152 16000
rect 34204 15988 34210 16040
rect 34609 16031 34667 16037
rect 34609 15997 34621 16031
rect 34655 16028 34667 16031
rect 35434 16028 35440 16040
rect 34655 16000 35440 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 17368 15932 22876 15960
rect 17368 15920 17374 15932
rect 34514 15920 34520 15972
rect 34572 15960 34578 15972
rect 34624 15960 34652 15991
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 34572 15932 34652 15960
rect 34572 15920 34578 15932
rect 35158 15920 35164 15972
rect 35216 15960 35222 15972
rect 35728 15960 35756 16059
rect 36446 16056 36452 16068
rect 36504 16056 36510 16108
rect 37642 16028 37648 16040
rect 37603 16000 37648 16028
rect 37642 15988 37648 16000
rect 37700 15988 37706 16040
rect 38286 16028 38292 16040
rect 38247 16000 38292 16028
rect 38286 15988 38292 16000
rect 38344 15988 38350 16040
rect 36170 15960 36176 15972
rect 35216 15932 36176 15960
rect 35216 15920 35222 15932
rect 36170 15920 36176 15932
rect 36228 15960 36234 15972
rect 36722 15960 36728 15972
rect 36228 15932 36728 15960
rect 36228 15920 36234 15932
rect 36722 15920 36728 15932
rect 36780 15920 36786 15972
rect 10652 15864 17264 15892
rect 10652 15852 10658 15864
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 19978 15892 19984 15904
rect 17644 15864 19984 15892
rect 17644 15852 17650 15864
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20073 15895 20131 15901
rect 20073 15861 20085 15895
rect 20119 15892 20131 15895
rect 20622 15892 20628 15904
rect 20119 15864 20628 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 20806 15892 20812 15904
rect 20767 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 26326 15852 26332 15904
rect 26384 15892 26390 15904
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 26384 15864 28365 15892
rect 26384 15852 26390 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 28353 15855 28411 15861
rect 29178 15852 29184 15904
rect 29236 15892 29242 15904
rect 30285 15895 30343 15901
rect 30285 15892 30297 15895
rect 29236 15864 30297 15892
rect 29236 15852 29242 15864
rect 30285 15861 30297 15864
rect 30331 15861 30343 15895
rect 30285 15855 30343 15861
rect 31757 15895 31815 15901
rect 31757 15861 31769 15895
rect 31803 15892 31815 15895
rect 32030 15892 32036 15904
rect 31803 15864 32036 15892
rect 31803 15861 31815 15864
rect 31757 15855 31815 15861
rect 32030 15852 32036 15864
rect 32088 15852 32094 15904
rect 32582 15852 32588 15904
rect 32640 15892 32646 15904
rect 38194 15892 38200 15904
rect 32640 15864 38200 15892
rect 32640 15852 32646 15864
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 14366 15688 14372 15700
rect 14327 15660 14372 15688
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 19794 15688 19800 15700
rect 14516 15660 17448 15688
rect 19755 15660 19800 15688
rect 14516 15648 14522 15660
rect 11333 15623 11391 15629
rect 11333 15620 11345 15623
rect 10428 15592 11345 15620
rect 10226 15552 10232 15564
rect 10187 15524 10232 15552
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 10428 15561 10456 15592
rect 11333 15589 11345 15592
rect 11379 15589 11391 15623
rect 11333 15583 11391 15589
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 17310 15620 17316 15632
rect 12308 15592 17316 15620
rect 12308 15580 12314 15592
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 17420 15620 17448 15660
rect 19794 15648 19800 15660
rect 19852 15648 19858 15700
rect 24946 15688 24952 15700
rect 19904 15660 24952 15688
rect 19904 15620 19932 15660
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 28813 15691 28871 15697
rect 28813 15657 28825 15691
rect 28859 15688 28871 15691
rect 32582 15688 32588 15700
rect 28859 15660 32588 15688
rect 28859 15657 28871 15660
rect 28813 15651 28871 15657
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 32692 15660 33732 15688
rect 17420 15592 19932 15620
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 26510 15620 26516 15632
rect 20036 15592 26516 15620
rect 20036 15580 20042 15592
rect 26510 15580 26516 15592
rect 26568 15580 26574 15632
rect 27246 15580 27252 15632
rect 27304 15620 27310 15632
rect 28534 15620 28540 15632
rect 27304 15592 28540 15620
rect 27304 15580 27310 15592
rect 28534 15580 28540 15592
rect 28592 15620 28598 15632
rect 30101 15623 30159 15629
rect 30101 15620 30113 15623
rect 28592 15592 30113 15620
rect 28592 15580 28598 15592
rect 30101 15589 30113 15592
rect 30147 15589 30159 15623
rect 30926 15620 30932 15632
rect 30887 15592 30932 15620
rect 30101 15583 30159 15589
rect 30926 15580 30932 15592
rect 30984 15580 30990 15632
rect 32214 15620 32220 15632
rect 31680 15592 32220 15620
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 28077 15555 28135 15561
rect 11756 15524 25268 15552
rect 11756 15512 11762 15524
rect 11514 15484 11520 15496
rect 11475 15456 11520 15484
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 12986 15484 12992 15496
rect 12947 15456 12992 15484
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14458 15484 14464 15496
rect 14323 15456 14464 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 18104 15456 18153 15484
rect 18104 15444 18110 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19484 15456 19993 15484
rect 19484 15444 19490 15456
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 21450 15484 21456 15496
rect 21411 15456 21456 15484
rect 20625 15447 20683 15453
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 20640 15416 20668 15447
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 25240 15493 25268 15524
rect 26344 15524 26556 15552
rect 25225 15487 25283 15493
rect 21600 15456 25176 15484
rect 21600 15444 21606 15456
rect 18012 15388 20668 15416
rect 20717 15419 20775 15425
rect 18012 15376 18018 15388
rect 20717 15385 20729 15419
rect 20763 15416 20775 15419
rect 23382 15416 23388 15428
rect 20763 15388 23388 15416
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 23382 15376 23388 15388
rect 23440 15376 23446 15428
rect 25148 15416 25176 15456
rect 25225 15453 25237 15487
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 26344 15416 26372 15524
rect 26421 15487 26479 15493
rect 26421 15453 26433 15487
rect 26467 15453 26479 15487
rect 26528 15484 26556 15524
rect 28077 15521 28089 15555
rect 28123 15552 28135 15555
rect 29917 15555 29975 15561
rect 29917 15552 29929 15555
rect 28123 15524 29929 15552
rect 28123 15521 28135 15524
rect 28077 15515 28135 15521
rect 29917 15521 29929 15524
rect 29963 15521 29975 15555
rect 31570 15552 31576 15564
rect 29917 15515 29975 15521
rect 30668 15524 31576 15552
rect 27985 15487 28043 15493
rect 27985 15484 27997 15487
rect 26528 15456 27997 15484
rect 26421 15447 26479 15453
rect 27985 15453 27997 15456
rect 28031 15453 28043 15487
rect 29270 15484 29276 15496
rect 27985 15447 28043 15453
rect 28092 15456 29276 15484
rect 25148 15388 26372 15416
rect 26436 15416 26464 15447
rect 28092 15416 28120 15456
rect 29270 15444 29276 15456
rect 29328 15444 29334 15496
rect 29362 15444 29368 15496
rect 29420 15484 29426 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29420 15456 29745 15484
rect 29420 15444 29426 15456
rect 29733 15453 29745 15456
rect 29779 15484 29791 15487
rect 30668 15484 30696 15524
rect 31570 15512 31576 15524
rect 31628 15512 31634 15564
rect 29779 15456 30696 15484
rect 29779 15453 29791 15456
rect 29733 15447 29791 15453
rect 30742 15444 30748 15496
rect 30800 15484 30806 15496
rect 31680 15493 31708 15592
rect 32214 15580 32220 15592
rect 32272 15580 32278 15632
rect 32692 15561 32720 15660
rect 33226 15620 33232 15632
rect 33187 15592 33232 15620
rect 33226 15580 33232 15592
rect 33284 15580 33290 15632
rect 33704 15620 33732 15660
rect 33778 15648 33784 15700
rect 33836 15688 33842 15700
rect 33873 15691 33931 15697
rect 33873 15688 33885 15691
rect 33836 15660 33885 15688
rect 33836 15648 33842 15660
rect 33873 15657 33885 15660
rect 33919 15657 33931 15691
rect 33873 15651 33931 15657
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 34977 15691 35035 15697
rect 34977 15688 34989 15691
rect 34848 15660 34989 15688
rect 34848 15648 34854 15660
rect 34977 15657 34989 15660
rect 35023 15657 35035 15691
rect 34977 15651 35035 15657
rect 37369 15691 37427 15697
rect 37369 15657 37381 15691
rect 37415 15688 37427 15691
rect 39022 15688 39028 15700
rect 37415 15660 39028 15688
rect 37415 15657 37427 15660
rect 37369 15651 37427 15657
rect 39022 15648 39028 15660
rect 39080 15648 39086 15700
rect 35710 15620 35716 15632
rect 33704 15592 35716 15620
rect 35710 15580 35716 15592
rect 35768 15580 35774 15632
rect 32677 15555 32735 15561
rect 32677 15521 32689 15555
rect 32723 15521 32735 15555
rect 32677 15515 32735 15521
rect 32858 15512 32864 15564
rect 32916 15552 32922 15564
rect 35897 15555 35955 15561
rect 32916 15524 33824 15552
rect 32916 15512 32922 15524
rect 33796 15493 33824 15524
rect 35897 15521 35909 15555
rect 35943 15552 35955 15555
rect 36354 15552 36360 15564
rect 35943 15524 36360 15552
rect 35943 15521 35955 15524
rect 35897 15515 35955 15521
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 30837 15487 30895 15493
rect 30837 15484 30849 15487
rect 30800 15456 30849 15484
rect 30800 15444 30806 15456
rect 30837 15453 30849 15456
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 31665 15487 31723 15493
rect 31665 15453 31677 15487
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 33781 15487 33839 15493
rect 33781 15453 33793 15487
rect 33827 15453 33839 15487
rect 34882 15484 34888 15496
rect 34843 15456 34888 15484
rect 33781 15447 33839 15453
rect 34882 15444 34888 15456
rect 34940 15444 34946 15496
rect 37458 15444 37464 15496
rect 37516 15484 37522 15496
rect 37553 15487 37611 15493
rect 37553 15484 37565 15487
rect 37516 15456 37565 15484
rect 37516 15444 37522 15456
rect 37553 15453 37565 15456
rect 37599 15453 37611 15487
rect 38010 15484 38016 15496
rect 37971 15456 38016 15484
rect 37553 15447 37611 15453
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 28718 15416 28724 15428
rect 26436 15388 28120 15416
rect 28679 15388 28724 15416
rect 28718 15376 28724 15388
rect 28776 15376 28782 15428
rect 31938 15416 31944 15428
rect 28828 15388 31944 15416
rect 10870 15348 10876 15360
rect 10831 15320 10876 15348
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 12805 15351 12863 15357
rect 12805 15317 12817 15351
rect 12851 15348 12863 15351
rect 13262 15348 13268 15360
rect 12851 15320 13268 15348
rect 12851 15317 12863 15320
rect 12805 15311 12863 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 18230 15348 18236 15360
rect 18191 15320 18236 15348
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21269 15351 21327 15357
rect 21269 15348 21281 15351
rect 21232 15320 21281 15348
rect 21232 15308 21238 15320
rect 21269 15317 21281 15320
rect 21315 15317 21327 15351
rect 25038 15348 25044 15360
rect 24999 15320 25044 15348
rect 21269 15311 21327 15317
rect 25038 15308 25044 15320
rect 25096 15308 25102 15360
rect 26513 15351 26571 15357
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 27338 15348 27344 15360
rect 26559 15320 27344 15348
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27614 15308 27620 15360
rect 27672 15348 27678 15360
rect 28828 15348 28856 15388
rect 31938 15376 31944 15388
rect 31996 15376 32002 15428
rect 32769 15419 32827 15425
rect 32769 15385 32781 15419
rect 32815 15385 32827 15419
rect 32769 15379 32827 15385
rect 27672 15320 28856 15348
rect 27672 15308 27678 15320
rect 31386 15308 31392 15360
rect 31444 15348 31450 15360
rect 31481 15351 31539 15357
rect 31481 15348 31493 15351
rect 31444 15320 31493 15348
rect 31444 15308 31450 15320
rect 31481 15317 31493 15320
rect 31527 15317 31539 15351
rect 31481 15311 31539 15317
rect 31754 15308 31760 15360
rect 31812 15348 31818 15360
rect 32784 15348 32812 15379
rect 34606 15376 34612 15428
rect 34664 15416 34670 15428
rect 35989 15419 36047 15425
rect 35989 15416 36001 15419
rect 34664 15388 36001 15416
rect 34664 15376 34670 15388
rect 35989 15385 36001 15388
rect 36035 15385 36047 15419
rect 35989 15379 36047 15385
rect 36541 15419 36599 15425
rect 36541 15385 36553 15419
rect 36587 15416 36599 15419
rect 37918 15416 37924 15428
rect 36587 15388 37924 15416
rect 36587 15385 36599 15388
rect 36541 15379 36599 15385
rect 37918 15376 37924 15388
rect 37976 15376 37982 15428
rect 31812 15320 32812 15348
rect 31812 15308 31818 15320
rect 32950 15308 32956 15360
rect 33008 15348 33014 15360
rect 35434 15348 35440 15360
rect 33008 15320 35440 15348
rect 33008 15308 33014 15320
rect 35434 15308 35440 15320
rect 35492 15308 35498 15360
rect 38194 15348 38200 15360
rect 38155 15320 38200 15348
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 11422 15144 11428 15156
rect 10827 15116 11428 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 11514 15104 11520 15156
rect 11572 15144 11578 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11572 15116 11713 15144
rect 11572 15104 11578 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 11701 15107 11759 15113
rect 11808 15116 14933 15144
rect 10870 15036 10876 15088
rect 10928 15076 10934 15088
rect 11808 15076 11836 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 17770 15104 17776 15156
rect 17828 15144 17834 15156
rect 18874 15144 18880 15156
rect 17828 15116 18880 15144
rect 17828 15104 17834 15116
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19426 15144 19432 15156
rect 18932 15116 19432 15144
rect 18932 15104 18938 15116
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 24210 15144 24216 15156
rect 20036 15116 24216 15144
rect 20036 15104 20042 15116
rect 13262 15076 13268 15088
rect 10928 15048 11836 15076
rect 13223 15048 13268 15076
rect 10928 15036 10934 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 20162 15076 20168 15088
rect 14200 15048 20168 15076
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 1728 14980 9597 15008
rect 1728 14968 1734 14980
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9585 14971 9643 14977
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 14977 10747 15011
rect 11882 15008 11888 15020
rect 11843 14980 11888 15008
rect 10689 14971 10747 14977
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 10704 14940 10732 14971
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 13170 14940 13176 14952
rect 8812 14912 10732 14940
rect 13131 14912 13176 14940
rect 8812 14900 8818 14912
rect 13170 14900 13176 14912
rect 13228 14900 13234 14952
rect 13446 14940 13452 14952
rect 13407 14912 13452 14940
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 9677 14875 9735 14881
rect 9677 14841 9689 14875
rect 9723 14872 9735 14875
rect 14200 14872 14228 15048
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 20622 15076 20628 15088
rect 20312 15048 20628 15076
rect 20312 15036 20318 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 15008 17371 15011
rect 18046 15008 18052 15020
rect 17359 14980 18052 15008
rect 17359 14977 17371 14980
rect 17313 14971 17371 14977
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20128 14980 20361 15008
rect 20128 14968 20134 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 15008 20591 15011
rect 20806 15008 20812 15020
rect 20579 14980 20812 15008
rect 20579 14977 20591 14980
rect 20533 14971 20591 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 22020 15017 22048 15116
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 28350 15144 28356 15156
rect 27172 15116 28356 15144
rect 22097 15079 22155 15085
rect 22097 15045 22109 15079
rect 22143 15076 22155 15079
rect 22925 15079 22983 15085
rect 22925 15076 22937 15079
rect 22143 15048 22937 15076
rect 22143 15045 22155 15048
rect 22097 15039 22155 15045
rect 22925 15045 22937 15048
rect 22971 15045 22983 15079
rect 27172 15076 27200 15116
rect 28350 15104 28356 15116
rect 28408 15104 28414 15156
rect 33042 15104 33048 15156
rect 33100 15144 33106 15156
rect 35621 15147 35679 15153
rect 35621 15144 35633 15147
rect 33100 15116 35633 15144
rect 33100 15104 33106 15116
rect 35621 15113 35633 15116
rect 35667 15113 35679 15147
rect 35621 15107 35679 15113
rect 36170 15104 36176 15156
rect 36228 15104 36234 15156
rect 36538 15104 36544 15156
rect 36596 15144 36602 15156
rect 37553 15147 37611 15153
rect 37553 15144 37565 15147
rect 36596 15116 37565 15144
rect 36596 15104 36602 15116
rect 37553 15113 37565 15116
rect 37599 15113 37611 15147
rect 37553 15107 37611 15113
rect 38102 15104 38108 15156
rect 38160 15144 38166 15156
rect 38197 15147 38255 15153
rect 38197 15144 38209 15147
rect 38160 15116 38209 15144
rect 38160 15104 38166 15116
rect 38197 15113 38209 15116
rect 38243 15113 38255 15147
rect 38197 15107 38255 15113
rect 27338 15076 27344 15088
rect 22925 15039 22983 15045
rect 26436 15048 27200 15076
rect 27299 15048 27344 15076
rect 26436 15017 26464 15048
rect 27338 15036 27344 15048
rect 27396 15036 27402 15088
rect 29178 15076 29184 15088
rect 29139 15048 29184 15076
rect 29178 15036 29184 15048
rect 29236 15036 29242 15088
rect 32490 15076 32496 15088
rect 32451 15048 32496 15076
rect 32490 15036 32496 15048
rect 32548 15036 32554 15088
rect 34422 15076 34428 15088
rect 33060 15048 34428 15076
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 30561 15011 30619 15017
rect 30561 14977 30573 15011
rect 30607 15008 30619 15011
rect 31202 15008 31208 15020
rect 30607 14980 31208 15008
rect 30607 14977 30619 14980
rect 30561 14971 30619 14977
rect 31202 14968 31208 14980
rect 31260 14968 31266 15020
rect 31386 15008 31392 15020
rect 31347 14980 31392 15008
rect 31386 14968 31392 14980
rect 31444 14968 31450 15020
rect 33060 15017 33088 15048
rect 34422 15036 34428 15048
rect 34480 15036 34486 15088
rect 34514 15036 34520 15088
rect 34572 15076 34578 15088
rect 36188 15076 36216 15104
rect 34572 15048 36400 15076
rect 34572 15036 34578 15048
rect 33045 15011 33103 15017
rect 33045 14977 33057 15011
rect 33091 14977 33103 15011
rect 33045 14971 33103 14977
rect 33226 14968 33232 15020
rect 33284 15008 33290 15020
rect 34149 15011 34207 15017
rect 34149 15008 34161 15011
rect 33284 14980 34161 15008
rect 33284 14968 33290 14980
rect 34149 14977 34161 14980
rect 34195 15008 34207 15011
rect 34238 15008 34244 15020
rect 34195 14980 34244 15008
rect 34195 14977 34207 14980
rect 34149 14971 34207 14977
rect 34238 14968 34244 14980
rect 34296 14968 34302 15020
rect 34882 15008 34888 15020
rect 34843 14980 34888 15008
rect 34882 14968 34888 14980
rect 34940 14968 34946 15020
rect 35544 15017 35572 15048
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 14977 35587 15011
rect 35529 14971 35587 14977
rect 36173 15011 36231 15017
rect 36173 14977 36185 15011
rect 36219 14977 36231 15011
rect 36173 14971 36231 14977
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 9723 14844 14228 14872
rect 14292 14872 14320 14903
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14424 14912 14473 14940
rect 14424 14900 14430 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 22830 14940 22836 14952
rect 22791 14912 22836 14940
rect 14461 14903 14519 14909
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23845 14943 23903 14949
rect 23845 14909 23857 14943
rect 23891 14940 23903 14943
rect 26878 14940 26884 14952
rect 23891 14912 26884 14940
rect 23891 14909 23903 14912
rect 23845 14903 23903 14909
rect 26878 14900 26884 14912
rect 26936 14900 26942 14952
rect 27246 14940 27252 14952
rect 27207 14912 27252 14940
rect 27246 14900 27252 14912
rect 27304 14900 27310 14952
rect 27614 14940 27620 14952
rect 27575 14912 27620 14940
rect 27614 14900 27620 14912
rect 27672 14900 27678 14952
rect 29089 14943 29147 14949
rect 29089 14909 29101 14943
rect 29135 14909 29147 14943
rect 29730 14940 29736 14952
rect 29691 14912 29736 14940
rect 29089 14903 29147 14909
rect 19242 14872 19248 14884
rect 14292 14844 19248 14872
rect 9723 14841 9735 14844
rect 9677 14835 9735 14841
rect 19242 14832 19248 14844
rect 19300 14872 19306 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 19300 14844 20729 14872
rect 19300 14832 19306 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 13630 14804 13636 14816
rect 13504 14776 13636 14804
rect 13504 14764 13510 14776
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17184 14776 17417 14804
rect 17184 14764 17190 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 26896 14804 26924 14900
rect 26970 14832 26976 14884
rect 27028 14872 27034 14884
rect 29104 14872 29132 14903
rect 29730 14900 29736 14912
rect 29788 14900 29794 14952
rect 32214 14940 32220 14952
rect 30208 14912 32220 14940
rect 30208 14872 30236 14912
rect 32214 14900 32220 14912
rect 32272 14900 32278 14952
rect 32401 14943 32459 14949
rect 32401 14909 32413 14943
rect 32447 14940 32459 14943
rect 33318 14940 33324 14952
rect 32447 14912 33324 14940
rect 32447 14909 32459 14912
rect 32401 14903 32459 14909
rect 33318 14900 33324 14912
rect 33376 14900 33382 14952
rect 33502 14940 33508 14952
rect 33463 14912 33508 14940
rect 33502 14900 33508 14912
rect 33560 14900 33566 14952
rect 34977 14943 35035 14949
rect 34977 14909 34989 14943
rect 35023 14940 35035 14943
rect 35618 14940 35624 14952
rect 35023 14912 35624 14940
rect 35023 14909 35035 14912
rect 34977 14903 35035 14909
rect 35618 14900 35624 14912
rect 35676 14900 35682 14952
rect 32122 14872 32128 14884
rect 27028 14844 30236 14872
rect 30576 14844 32128 14872
rect 27028 14832 27034 14844
rect 30576 14804 30604 14844
rect 32122 14832 32128 14844
rect 32180 14832 32186 14884
rect 32306 14832 32312 14884
rect 32364 14872 32370 14884
rect 36188 14872 36216 14971
rect 36372 14940 36400 15048
rect 36446 15036 36452 15088
rect 36504 15076 36510 15088
rect 36504 15048 38148 15076
rect 36504 15036 36510 15048
rect 38120 15020 38148 15048
rect 36630 14968 36636 15020
rect 36688 15008 36694 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 36688 14980 37473 15008
rect 36688 14968 36694 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 38102 15008 38108 15020
rect 38015 14980 38108 15008
rect 37461 14971 37519 14977
rect 38102 14968 38108 14980
rect 38160 15008 38166 15020
rect 39758 15008 39764 15020
rect 38160 14980 39764 15008
rect 38160 14968 38166 14980
rect 39758 14968 39764 14980
rect 39816 14968 39822 15020
rect 37182 14940 37188 14952
rect 36372 14912 37188 14940
rect 37182 14900 37188 14912
rect 37240 14900 37246 14952
rect 32364 14844 36216 14872
rect 32364 14832 32370 14844
rect 26896 14776 30604 14804
rect 30653 14807 30711 14813
rect 17405 14767 17463 14773
rect 30653 14773 30665 14807
rect 30699 14804 30711 14807
rect 30834 14804 30840 14816
rect 30699 14776 30840 14804
rect 30699 14773 30711 14776
rect 30653 14767 30711 14773
rect 30834 14764 30840 14776
rect 30892 14764 30898 14816
rect 31205 14807 31263 14813
rect 31205 14773 31217 14807
rect 31251 14804 31263 14807
rect 31846 14804 31852 14816
rect 31251 14776 31852 14804
rect 31251 14773 31263 14776
rect 31205 14767 31263 14773
rect 31846 14764 31852 14776
rect 31904 14764 31910 14816
rect 33410 14764 33416 14816
rect 33468 14804 33474 14816
rect 34241 14807 34299 14813
rect 34241 14804 34253 14807
rect 33468 14776 34253 14804
rect 33468 14764 33474 14776
rect 34241 14773 34253 14776
rect 34287 14773 34299 14807
rect 34241 14767 34299 14773
rect 36265 14807 36323 14813
rect 36265 14773 36277 14807
rect 36311 14804 36323 14807
rect 36998 14804 37004 14816
rect 36311 14776 37004 14804
rect 36311 14773 36323 14776
rect 36265 14767 36323 14773
rect 36998 14764 37004 14776
rect 37056 14764 37062 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 14366 14600 14372 14612
rect 14327 14572 14372 14600
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 27798 14560 27804 14612
rect 27856 14600 27862 14612
rect 28261 14603 28319 14609
rect 28261 14600 28273 14603
rect 27856 14572 28273 14600
rect 27856 14560 27862 14572
rect 28261 14569 28273 14572
rect 28307 14569 28319 14603
rect 28261 14563 28319 14569
rect 31113 14603 31171 14609
rect 31113 14569 31125 14603
rect 31159 14600 31171 14603
rect 31754 14600 31760 14612
rect 31159 14572 31760 14600
rect 31159 14569 31171 14572
rect 31113 14563 31171 14569
rect 31754 14560 31760 14572
rect 31812 14560 31818 14612
rect 32030 14600 32036 14612
rect 31991 14572 32036 14600
rect 32030 14560 32036 14572
rect 32088 14560 32094 14612
rect 32214 14560 32220 14612
rect 32272 14600 32278 14612
rect 34977 14603 35035 14609
rect 34977 14600 34989 14603
rect 32272 14572 34989 14600
rect 32272 14560 32278 14572
rect 34977 14569 34989 14572
rect 35023 14569 35035 14603
rect 36354 14600 36360 14612
rect 36315 14572 36360 14600
rect 34977 14563 35035 14569
rect 36354 14560 36360 14572
rect 36412 14560 36418 14612
rect 37829 14603 37887 14609
rect 37829 14569 37841 14603
rect 37875 14600 37887 14603
rect 39850 14600 39856 14612
rect 37875 14572 39856 14600
rect 37875 14569 37887 14572
rect 37829 14563 37887 14569
rect 39850 14560 39856 14572
rect 39908 14560 39914 14612
rect 14921 14535 14979 14541
rect 14921 14532 14933 14535
rect 6886 14504 14933 14532
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 6886 14396 6914 14504
rect 14921 14501 14933 14504
rect 14967 14501 14979 14535
rect 14921 14495 14979 14501
rect 25682 14492 25688 14544
rect 25740 14532 25746 14544
rect 33502 14532 33508 14544
rect 25740 14504 27292 14532
rect 25740 14492 25746 14504
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 15654 14464 15660 14476
rect 11940 14436 15660 14464
rect 11940 14424 11946 14436
rect 14292 14405 14320 14436
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 16908 14436 17049 14464
rect 16908 14424 16914 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17862 14464 17868 14476
rect 17823 14436 17868 14464
rect 17037 14427 17095 14433
rect 17862 14424 17868 14436
rect 17920 14464 17926 14476
rect 25317 14467 25375 14473
rect 25317 14464 25329 14467
rect 17920 14436 25329 14464
rect 17920 14424 17926 14436
rect 25317 14433 25329 14436
rect 25363 14433 25375 14467
rect 26970 14464 26976 14476
rect 26931 14436 26976 14464
rect 25317 14427 25375 14433
rect 26970 14424 26976 14436
rect 27028 14424 27034 14476
rect 27264 14473 27292 14504
rect 31680 14504 33508 14532
rect 27249 14467 27307 14473
rect 27249 14433 27261 14467
rect 27295 14433 27307 14467
rect 30742 14464 30748 14476
rect 27249 14427 27307 14433
rect 28184 14436 30748 14464
rect 1627 14368 6914 14396
rect 14277 14399 14335 14405
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 15105 14359 15163 14365
rect 17880 14368 18705 14396
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 15120 14260 15148 14359
rect 17880 14340 17908 14368
rect 18693 14365 18705 14368
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 28184 14405 28212 14436
rect 30742 14424 30748 14436
rect 30800 14424 30806 14476
rect 31680 14473 31708 14504
rect 33502 14492 33508 14504
rect 33560 14492 33566 14544
rect 35986 14492 35992 14544
rect 36044 14532 36050 14544
rect 37185 14535 37243 14541
rect 37185 14532 37197 14535
rect 36044 14504 37197 14532
rect 36044 14492 36050 14504
rect 37185 14501 37197 14504
rect 37231 14501 37243 14535
rect 37185 14495 37243 14501
rect 31665 14467 31723 14473
rect 31665 14433 31677 14467
rect 31711 14433 31723 14467
rect 31846 14464 31852 14476
rect 31807 14436 31852 14464
rect 31665 14427 31723 14433
rect 31846 14424 31852 14436
rect 31904 14424 31910 14476
rect 32122 14424 32128 14476
rect 32180 14464 32186 14476
rect 33597 14467 33655 14473
rect 33597 14464 33609 14467
rect 32180 14436 33609 14464
rect 32180 14424 32186 14436
rect 33597 14433 33609 14436
rect 33643 14464 33655 14467
rect 33962 14464 33968 14476
rect 33643 14436 33968 14464
rect 33643 14433 33655 14436
rect 33597 14427 33655 14433
rect 33962 14424 33968 14436
rect 34020 14424 34026 14476
rect 34238 14424 34244 14476
rect 34296 14464 34302 14476
rect 36173 14467 36231 14473
rect 36173 14464 36185 14467
rect 34296 14436 36185 14464
rect 34296 14424 34302 14436
rect 36173 14433 36185 14436
rect 36219 14433 36231 14467
rect 39298 14464 39304 14476
rect 36173 14427 36231 14433
rect 37108 14436 39304 14464
rect 22465 14399 22523 14405
rect 22465 14396 22477 14399
rect 21508 14368 22477 14396
rect 21508 14356 21514 14368
rect 22465 14365 22477 14368
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28626 14356 28632 14408
rect 28684 14396 28690 14408
rect 28813 14399 28871 14405
rect 28813 14396 28825 14399
rect 28684 14368 28825 14396
rect 28684 14356 28690 14368
rect 28813 14365 28825 14368
rect 28859 14365 28871 14399
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 28813 14359 28871 14365
rect 28920 14368 29745 14396
rect 17126 14288 17132 14340
rect 17184 14328 17190 14340
rect 17184 14300 17229 14328
rect 17184 14288 17190 14300
rect 17862 14288 17868 14340
rect 17920 14288 17926 14340
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 23658 14328 23664 14340
rect 19484 14300 23664 14328
rect 19484 14288 19490 14300
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 25041 14331 25099 14337
rect 25041 14297 25053 14331
rect 25087 14297 25099 14331
rect 25041 14291 25099 14297
rect 25133 14331 25191 14337
rect 25133 14297 25145 14331
rect 25179 14328 25191 14331
rect 25222 14328 25228 14340
rect 25179 14300 25228 14328
rect 25179 14297 25191 14300
rect 25133 14291 25191 14297
rect 17494 14260 17500 14272
rect 15120 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 18506 14260 18512 14272
rect 18467 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 22554 14260 22560 14272
rect 22515 14232 22560 14260
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 25056 14260 25084 14291
rect 25222 14288 25228 14300
rect 25280 14288 25286 14340
rect 27062 14288 27068 14340
rect 27120 14328 27126 14340
rect 27120 14300 27165 14328
rect 27120 14288 27126 14300
rect 27430 14288 27436 14340
rect 27488 14328 27494 14340
rect 28920 14328 28948 14368
rect 29733 14365 29745 14368
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30558 14396 30564 14408
rect 30423 14368 30564 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 31021 14399 31079 14405
rect 31021 14365 31033 14399
rect 31067 14396 31079 14399
rect 32306 14396 32312 14408
rect 31067 14368 32312 14396
rect 31067 14365 31079 14368
rect 31021 14359 31079 14365
rect 32306 14356 32312 14368
rect 32364 14356 32370 14408
rect 34885 14399 34943 14405
rect 34885 14365 34897 14399
rect 34931 14396 34943 14399
rect 35618 14396 35624 14408
rect 34931 14368 35624 14396
rect 34931 14365 34943 14368
rect 34885 14359 34943 14365
rect 35618 14356 35624 14368
rect 35676 14356 35682 14408
rect 35710 14356 35716 14408
rect 35768 14396 35774 14408
rect 37108 14405 37136 14436
rect 39298 14424 39304 14436
rect 39356 14424 39362 14476
rect 35989 14399 36047 14405
rect 35989 14396 36001 14399
rect 35768 14368 36001 14396
rect 35768 14356 35774 14368
rect 35989 14365 36001 14368
rect 36035 14365 36047 14399
rect 35989 14359 36047 14365
rect 37093 14399 37151 14405
rect 37093 14365 37105 14399
rect 37139 14365 37151 14399
rect 37093 14359 37151 14365
rect 37737 14399 37795 14405
rect 37737 14365 37749 14399
rect 37783 14396 37795 14399
rect 38102 14396 38108 14408
rect 37783 14368 38108 14396
rect 37783 14365 37795 14368
rect 37737 14359 37795 14365
rect 38102 14356 38108 14368
rect 38160 14356 38166 14408
rect 27488 14300 28948 14328
rect 27488 14288 27494 14300
rect 29454 14288 29460 14340
rect 29512 14328 29518 14340
rect 33318 14328 33324 14340
rect 29512 14300 31754 14328
rect 33279 14300 33324 14328
rect 29512 14288 29518 14300
rect 25498 14260 25504 14272
rect 25056 14232 25504 14260
rect 25498 14220 25504 14232
rect 25556 14260 25562 14272
rect 28905 14263 28963 14269
rect 28905 14260 28917 14263
rect 25556 14232 28917 14260
rect 25556 14220 25562 14232
rect 28905 14229 28917 14232
rect 28951 14229 28963 14263
rect 28905 14223 28963 14229
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 29825 14263 29883 14269
rect 29825 14260 29837 14263
rect 29052 14232 29837 14260
rect 29052 14220 29058 14232
rect 29825 14229 29837 14232
rect 29871 14229 29883 14263
rect 29825 14223 29883 14229
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 30469 14263 30527 14269
rect 30469 14260 30481 14263
rect 30432 14232 30481 14260
rect 30432 14220 30438 14232
rect 30469 14229 30481 14232
rect 30515 14229 30527 14263
rect 31726 14260 31754 14300
rect 33318 14288 33324 14300
rect 33376 14288 33382 14340
rect 33410 14288 33416 14340
rect 33468 14328 33474 14340
rect 33468 14300 33513 14328
rect 33468 14288 33474 14300
rect 34146 14260 34152 14272
rect 31726 14232 34152 14260
rect 30469 14223 30527 14229
rect 34146 14220 34152 14232
rect 34204 14220 34210 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 8478 14056 8484 14068
rect 1627 14028 8484 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14025 14427 14059
rect 19242 14056 19248 14068
rect 19203 14028 19248 14056
rect 14369 14019 14427 14025
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 14384 13988 14412 14019
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 22189 14059 22247 14065
rect 20680 14028 21680 14056
rect 20680 14016 20686 14028
rect 13403 13960 14228 13988
rect 14384 13960 15240 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10870 13920 10876 13932
rect 10735 13892 10876 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 8352 13824 10793 13852
rect 8352 13812 8358 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 10781 13815 10839 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13722 13852 13728 13864
rect 13683 13824 13728 13852
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14200 13852 14228 13960
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 15212 13929 15240 13960
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17126 13988 17132 14000
rect 17000 13960 17132 13988
rect 17000 13948 17006 13960
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 17221 13991 17279 13997
rect 17221 13957 17233 13991
rect 17267 13988 17279 13991
rect 18230 13988 18236 14000
rect 17267 13960 18236 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 18230 13948 18236 13960
rect 18288 13948 18294 14000
rect 20714 13948 20720 14000
rect 20772 13948 20778 14000
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14516 13892 14565 13920
rect 14516 13880 14522 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20732 13920 20760 13948
rect 19935 13892 20760 13920
rect 20809 13923 20867 13929
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20809 13889 20821 13923
rect 20855 13920 20867 13923
rect 21542 13920 21548 13932
rect 20855 13892 21548 13920
rect 20855 13889 20867 13892
rect 20809 13883 20867 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 21652 13920 21680 14028
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 25222 14056 25228 14068
rect 22235 14028 25228 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 32766 14056 32772 14068
rect 29748 14028 32772 14056
rect 22554 13948 22560 14000
rect 22612 13988 22618 14000
rect 23385 13991 23443 13997
rect 23385 13988 23397 13991
rect 22612 13960 23397 13988
rect 22612 13948 22618 13960
rect 23385 13957 23397 13960
rect 23431 13957 23443 13991
rect 23385 13951 23443 13957
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 23532 13960 23577 13988
rect 23532 13948 23538 13960
rect 25314 13948 25320 14000
rect 25372 13988 25378 14000
rect 25682 13988 25688 14000
rect 25372 13960 25688 13988
rect 25372 13948 25378 13960
rect 25682 13948 25688 13960
rect 25740 13948 25746 14000
rect 25777 13991 25835 13997
rect 25777 13957 25789 13991
rect 25823 13988 25835 13991
rect 26326 13988 26332 14000
rect 25823 13960 26332 13988
rect 25823 13957 25835 13960
rect 25777 13951 25835 13957
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 27801 13991 27859 13997
rect 27801 13957 27813 13991
rect 27847 13988 27859 13991
rect 28902 13988 28908 14000
rect 27847 13960 28908 13988
rect 27847 13957 27859 13960
rect 27801 13951 27859 13957
rect 28902 13948 28908 13960
rect 28960 13988 28966 14000
rect 29181 13991 29239 13997
rect 29181 13988 29193 13991
rect 28960 13960 29193 13988
rect 28960 13948 28966 13960
rect 29181 13957 29193 13960
rect 29227 13957 29239 13991
rect 29181 13951 29239 13957
rect 22097 13923 22155 13929
rect 21652 13918 22048 13920
rect 22097 13918 22109 13923
rect 21652 13892 22109 13918
rect 22020 13890 22109 13892
rect 22097 13889 22109 13890
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 28534 13920 28540 13932
rect 28495 13892 28540 13920
rect 27157 13883 27215 13889
rect 14200 13824 15056 13852
rect 15028 13793 15056 13824
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17770 13852 17776 13864
rect 17644 13824 17776 13852
rect 17644 13812 17650 13824
rect 17770 13812 17776 13824
rect 17828 13852 17834 13864
rect 17957 13855 18015 13861
rect 17957 13852 17969 13855
rect 17828 13824 17969 13852
rect 17828 13812 17834 13824
rect 17957 13821 17969 13824
rect 18003 13821 18015 13855
rect 18598 13852 18604 13864
rect 18559 13824 18604 13852
rect 17957 13815 18015 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19426 13852 19432 13864
rect 18831 13824 19432 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 23658 13852 23664 13864
rect 20772 13824 23520 13852
rect 23619 13824 23664 13852
rect 20772 13812 20778 13824
rect 15013 13787 15071 13793
rect 15013 13753 15025 13787
rect 15059 13753 15071 13787
rect 23492 13784 23520 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 26142 13852 26148 13864
rect 23768 13824 26004 13852
rect 26103 13824 26148 13852
rect 23768 13784 23796 13824
rect 23492 13756 23796 13784
rect 25976 13784 26004 13824
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 27172 13852 27200 13883
rect 28534 13880 28540 13892
rect 28592 13880 28598 13932
rect 28721 13923 28779 13929
rect 28721 13889 28733 13923
rect 28767 13920 28779 13923
rect 28994 13920 29000 13932
rect 28767 13892 29000 13920
rect 28767 13889 28779 13892
rect 28721 13883 28779 13889
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 29748 13929 29776 14028
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 34330 14016 34336 14068
rect 34388 14056 34394 14068
rect 38197 14059 38255 14065
rect 34388 14028 36492 14056
rect 34388 14016 34394 14028
rect 36464 14000 36492 14028
rect 38197 14025 38209 14059
rect 38243 14056 38255 14059
rect 38562 14056 38568 14068
rect 38243 14028 38568 14056
rect 38243 14025 38255 14028
rect 38197 14019 38255 14025
rect 38562 14016 38568 14028
rect 38620 14016 38626 14068
rect 30834 13988 30840 14000
rect 30795 13960 30840 13988
rect 30834 13948 30840 13960
rect 30892 13948 30898 14000
rect 33962 13988 33968 14000
rect 33923 13960 33968 13988
rect 33962 13948 33968 13960
rect 34020 13948 34026 14000
rect 35526 13988 35532 14000
rect 35487 13960 35532 13988
rect 35526 13948 35532 13960
rect 35584 13948 35590 14000
rect 36446 13988 36452 14000
rect 36359 13960 36452 13988
rect 36446 13948 36452 13960
rect 36504 13948 36510 14000
rect 37553 13991 37611 13997
rect 37553 13957 37565 13991
rect 37599 13988 37611 13991
rect 38654 13988 38660 14000
rect 37599 13960 38660 13988
rect 37599 13957 37611 13960
rect 37553 13951 37611 13957
rect 38654 13948 38660 13960
rect 38712 13948 38718 14000
rect 29733 13923 29791 13929
rect 29733 13889 29745 13923
rect 29779 13889 29791 13923
rect 29733 13883 29791 13889
rect 32309 13923 32367 13929
rect 32309 13889 32321 13923
rect 32355 13920 32367 13923
rect 33226 13920 33232 13932
rect 32355 13892 33232 13920
rect 32355 13889 32367 13892
rect 32309 13883 32367 13889
rect 33226 13880 33232 13892
rect 33284 13880 33290 13932
rect 36630 13880 36636 13932
rect 36688 13920 36694 13932
rect 37461 13923 37519 13929
rect 37461 13920 37473 13923
rect 36688 13892 37473 13920
rect 36688 13880 36694 13892
rect 37461 13889 37473 13892
rect 37507 13920 37519 13923
rect 38102 13920 38108 13932
rect 37507 13892 38108 13920
rect 37507 13889 37519 13892
rect 37461 13883 37519 13889
rect 38102 13880 38108 13892
rect 38160 13880 38166 13932
rect 27338 13852 27344 13864
rect 26252 13824 27200 13852
rect 27299 13824 27344 13852
rect 26252 13784 26280 13824
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 29825 13855 29883 13861
rect 29825 13821 29837 13855
rect 29871 13852 29883 13855
rect 30745 13855 30803 13861
rect 30745 13852 30757 13855
rect 29871 13824 30757 13852
rect 29871 13821 29883 13824
rect 29825 13815 29883 13821
rect 30745 13821 30757 13824
rect 30791 13821 30803 13855
rect 31662 13852 31668 13864
rect 31623 13824 31668 13852
rect 30745 13815 30803 13821
rect 31662 13812 31668 13824
rect 31720 13812 31726 13864
rect 31846 13812 31852 13864
rect 31904 13852 31910 13864
rect 32401 13855 32459 13861
rect 32401 13852 32413 13855
rect 31904 13824 32413 13852
rect 31904 13812 31910 13824
rect 32401 13821 32413 13824
rect 32447 13821 32459 13855
rect 32401 13815 32459 13821
rect 33137 13855 33195 13861
rect 33137 13821 33149 13855
rect 33183 13852 33195 13855
rect 33873 13855 33931 13861
rect 33873 13852 33885 13855
rect 33183 13824 33885 13852
rect 33183 13821 33195 13824
rect 33137 13815 33195 13821
rect 33873 13821 33885 13824
rect 33919 13821 33931 13855
rect 34146 13852 34152 13864
rect 34107 13824 34152 13852
rect 33873 13815 33931 13821
rect 34146 13812 34152 13824
rect 34204 13812 34210 13864
rect 35434 13852 35440 13864
rect 35395 13824 35440 13852
rect 35434 13812 35440 13824
rect 35492 13812 35498 13864
rect 25976 13756 26280 13784
rect 15013 13747 15071 13753
rect 33502 13744 33508 13796
rect 33560 13784 33566 13796
rect 33686 13784 33692 13796
rect 33560 13756 33692 13784
rect 33560 13744 33566 13756
rect 33686 13744 33692 13756
rect 33744 13744 33750 13796
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 19705 13719 19763 13725
rect 19705 13716 19717 13719
rect 19668 13688 19717 13716
rect 19668 13676 19674 13688
rect 19705 13685 19717 13688
rect 19751 13685 19763 13719
rect 20898 13716 20904 13728
rect 20859 13688 20904 13716
rect 19705 13679 19763 13685
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 13228 13484 14933 13512
rect 13228 13472 13234 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 17865 13515 17923 13521
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 18322 13512 18328 13524
rect 17911 13484 18328 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 18322 13472 18328 13484
rect 18380 13512 18386 13524
rect 18598 13512 18604 13524
rect 18380 13484 18604 13512
rect 18380 13472 18386 13484
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 20714 13472 20720 13484
rect 20772 13512 20778 13524
rect 20990 13512 20996 13524
rect 20772 13484 20996 13512
rect 20772 13472 20778 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 26789 13515 26847 13521
rect 26789 13481 26801 13515
rect 26835 13512 26847 13515
rect 27338 13512 27344 13524
rect 26835 13484 27344 13512
rect 26835 13481 26847 13484
rect 26789 13475 26847 13481
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 32858 13512 32864 13524
rect 32819 13484 32864 13512
rect 32858 13472 32864 13484
rect 32916 13472 32922 13524
rect 33962 13472 33968 13524
rect 34020 13512 34026 13524
rect 34149 13515 34207 13521
rect 34149 13512 34161 13515
rect 34020 13484 34161 13512
rect 34020 13472 34026 13484
rect 34149 13481 34161 13484
rect 34195 13481 34207 13515
rect 34149 13475 34207 13481
rect 34977 13515 35035 13521
rect 34977 13481 34989 13515
rect 35023 13512 35035 13515
rect 35526 13512 35532 13524
rect 35023 13484 35532 13512
rect 35023 13481 35035 13484
rect 34977 13475 35035 13481
rect 35526 13472 35532 13484
rect 35584 13472 35590 13524
rect 36354 13472 36360 13524
rect 36412 13512 36418 13524
rect 36449 13515 36507 13521
rect 36449 13512 36461 13515
rect 36412 13484 36461 13512
rect 36412 13472 36418 13484
rect 36449 13481 36461 13484
rect 36495 13481 36507 13515
rect 36449 13475 36507 13481
rect 37277 13515 37335 13521
rect 37277 13481 37289 13515
rect 37323 13512 37335 13515
rect 39206 13512 39212 13524
rect 37323 13484 39212 13512
rect 37323 13481 37335 13484
rect 37277 13475 37335 13481
rect 39206 13472 39212 13484
rect 39264 13472 39270 13524
rect 13630 13404 13636 13456
rect 13688 13444 13694 13456
rect 13814 13444 13820 13456
rect 13688 13416 13820 13444
rect 13688 13404 13694 13416
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 24854 13404 24860 13456
rect 24912 13444 24918 13456
rect 25593 13447 25651 13453
rect 25593 13444 25605 13447
rect 24912 13416 25605 13444
rect 24912 13404 24918 13416
rect 25593 13413 25605 13416
rect 25639 13444 25651 13447
rect 26142 13444 26148 13456
rect 25639 13416 26148 13444
rect 25639 13413 25651 13416
rect 25593 13407 25651 13413
rect 26142 13404 26148 13416
rect 26200 13404 26206 13456
rect 26237 13447 26295 13453
rect 26237 13413 26249 13447
rect 26283 13444 26295 13447
rect 27062 13444 27068 13456
rect 26283 13416 27068 13444
rect 26283 13413 26295 13416
rect 26237 13407 26295 13413
rect 27062 13404 27068 13416
rect 27120 13404 27126 13456
rect 32125 13447 32183 13453
rect 32125 13413 32137 13447
rect 32171 13444 32183 13447
rect 33134 13444 33140 13456
rect 32171 13416 33140 13444
rect 32171 13413 32183 13416
rect 32125 13407 32183 13413
rect 33134 13404 33140 13416
rect 33192 13404 33198 13456
rect 33413 13447 33471 13453
rect 33413 13413 33425 13447
rect 33459 13444 33471 13447
rect 33459 13416 36400 13444
rect 33459 13413 33471 13416
rect 33413 13407 33471 13413
rect 36372 13388 36400 13416
rect 13262 13376 13268 13388
rect 13223 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15654 13376 15660 13388
rect 14599 13348 15660 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 20073 13379 20131 13385
rect 20073 13345 20085 13379
rect 20119 13376 20131 13379
rect 20162 13376 20168 13388
rect 20119 13348 20168 13376
rect 20119 13345 20131 13348
rect 20073 13339 20131 13345
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 20898 13376 20904 13388
rect 20303 13348 20904 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 32950 13376 32956 13388
rect 26160 13348 27476 13376
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 15010 13308 15016 13320
rect 14783 13280 15016 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 17862 13308 17868 13320
rect 17819 13280 17868 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 17862 13268 17868 13280
rect 17920 13268 17926 13320
rect 19610 13308 19616 13320
rect 19571 13280 19616 13308
rect 19610 13268 19616 13280
rect 19668 13268 19674 13320
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23474 13308 23480 13320
rect 22879 13280 23480 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 23474 13268 23480 13280
rect 23532 13308 23538 13320
rect 24026 13308 24032 13320
rect 23532 13280 24032 13308
rect 23532 13268 23538 13280
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 26050 13268 26056 13320
rect 26108 13308 26114 13320
rect 26160 13317 26188 13348
rect 26145 13311 26203 13317
rect 26145 13308 26157 13311
rect 26108 13280 26157 13308
rect 26108 13268 26114 13280
rect 26145 13277 26157 13280
rect 26191 13277 26203 13311
rect 26145 13271 26203 13277
rect 26418 13268 26424 13320
rect 26476 13308 26482 13320
rect 27448 13317 27476 13348
rect 32324 13348 32956 13376
rect 32324 13317 32352 13348
rect 32950 13336 32956 13348
rect 33008 13336 33014 13388
rect 35526 13376 35532 13388
rect 33612 13348 35532 13376
rect 33612 13317 33640 13348
rect 35526 13336 35532 13348
rect 35584 13336 35590 13388
rect 35986 13336 35992 13388
rect 36044 13376 36050 13388
rect 36265 13379 36323 13385
rect 36265 13376 36277 13379
rect 36044 13348 36277 13376
rect 36044 13336 36050 13348
rect 36265 13345 36277 13348
rect 36311 13345 36323 13379
rect 36265 13339 36323 13345
rect 36354 13336 36360 13388
rect 36412 13336 36418 13388
rect 26973 13311 27031 13317
rect 26973 13308 26985 13311
rect 26476 13280 26985 13308
rect 26476 13268 26482 13280
rect 26973 13277 26985 13280
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27433 13311 27491 13317
rect 27433 13277 27445 13311
rect 27479 13277 27491 13311
rect 27433 13271 27491 13277
rect 32309 13311 32367 13317
rect 32309 13277 32321 13311
rect 32355 13277 32367 13311
rect 32309 13271 32367 13277
rect 32769 13311 32827 13317
rect 32769 13277 32781 13311
rect 32815 13277 32827 13311
rect 32769 13271 32827 13277
rect 33597 13311 33655 13317
rect 33597 13277 33609 13311
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 25041 13243 25099 13249
rect 25041 13240 25053 13243
rect 24964 13212 25053 13240
rect 24964 13184 24992 13212
rect 25041 13209 25053 13212
rect 25087 13209 25099 13243
rect 25041 13203 25099 13209
rect 25130 13200 25136 13252
rect 25188 13240 25194 13252
rect 25188 13212 25233 13240
rect 25188 13200 25194 13212
rect 27890 13200 27896 13252
rect 27948 13240 27954 13252
rect 32784 13240 32812 13271
rect 33686 13268 33692 13320
rect 33744 13308 33750 13320
rect 34057 13311 34115 13317
rect 34057 13308 34069 13311
rect 33744 13280 34069 13308
rect 33744 13268 33750 13280
rect 34057 13277 34069 13280
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 34885 13311 34943 13317
rect 34885 13277 34897 13311
rect 34931 13308 34943 13311
rect 35802 13308 35808 13320
rect 34931 13280 35808 13308
rect 34931 13277 34943 13280
rect 34885 13271 34943 13277
rect 35802 13268 35808 13280
rect 35860 13268 35866 13320
rect 36081 13311 36139 13317
rect 36081 13277 36093 13311
rect 36127 13277 36139 13311
rect 36081 13271 36139 13277
rect 27948 13212 32812 13240
rect 27948 13200 27954 13212
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 12216 13144 12265 13172
rect 12216 13132 12222 13144
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 22922 13172 22928 13184
rect 22883 13144 22928 13172
rect 12253 13135 12311 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 24946 13132 24952 13184
rect 25004 13132 25010 13184
rect 26878 13132 26884 13184
rect 26936 13172 26942 13184
rect 27525 13175 27583 13181
rect 27525 13172 27537 13175
rect 26936 13144 27537 13172
rect 26936 13132 26942 13144
rect 27525 13141 27537 13144
rect 27571 13141 27583 13175
rect 32784 13172 32812 13212
rect 32858 13200 32864 13252
rect 32916 13240 32922 13252
rect 36094 13240 36122 13271
rect 37182 13268 37188 13320
rect 37240 13308 37246 13320
rect 37240 13280 37285 13308
rect 37240 13268 37246 13280
rect 37826 13268 37832 13320
rect 37884 13308 37890 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 37884 13280 38025 13308
rect 37884 13268 37890 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 32916 13212 36122 13240
rect 37200 13212 38056 13240
rect 32916 13200 32922 13212
rect 34790 13172 34796 13184
rect 32784 13144 34796 13172
rect 27525 13135 27583 13141
rect 34790 13132 34796 13144
rect 34848 13132 34854 13184
rect 34882 13132 34888 13184
rect 34940 13172 34946 13184
rect 37200 13172 37228 13212
rect 38028 13184 38056 13212
rect 34940 13144 37228 13172
rect 34940 13132 34946 13144
rect 38010 13132 38016 13184
rect 38068 13132 38074 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12937 6975 12971
rect 6917 12931 6975 12937
rect 9309 12971 9367 12977
rect 9309 12937 9321 12971
rect 9355 12968 9367 12971
rect 10502 12968 10508 12980
rect 9355 12940 10508 12968
rect 9355 12937 9367 12940
rect 9309 12931 9367 12937
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 6932 12832 6960 12931
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 12805 12971 12863 12977
rect 12805 12937 12817 12971
rect 12851 12968 12863 12971
rect 13170 12968 13176 12980
rect 12851 12940 13176 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 15010 12968 15016 12980
rect 14971 12940 15016 12968
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 20257 12971 20315 12977
rect 20257 12968 20269 12971
rect 19208 12940 20269 12968
rect 19208 12928 19214 12940
rect 20257 12937 20269 12940
rect 20303 12937 20315 12971
rect 26418 12968 26424 12980
rect 26379 12940 26424 12968
rect 20257 12931 20315 12937
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 29362 12968 29368 12980
rect 29323 12940 29368 12968
rect 29362 12928 29368 12940
rect 29420 12928 29426 12980
rect 32306 12968 32312 12980
rect 32267 12940 32312 12968
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 32953 12971 33011 12977
rect 32953 12937 32965 12971
rect 32999 12968 33011 12971
rect 34882 12968 34888 12980
rect 32999 12940 34888 12968
rect 32999 12937 33011 12940
rect 32953 12931 33011 12937
rect 34882 12928 34888 12940
rect 34940 12928 34946 12980
rect 34977 12971 35035 12977
rect 34977 12937 34989 12971
rect 35023 12968 35035 12971
rect 35342 12968 35348 12980
rect 35023 12940 35348 12968
rect 35023 12937 35035 12940
rect 34977 12931 35035 12937
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 35621 12971 35679 12977
rect 35621 12937 35633 12971
rect 35667 12968 35679 12971
rect 35894 12968 35900 12980
rect 35667 12940 35900 12968
rect 35667 12937 35679 12940
rect 35621 12931 35679 12937
rect 35894 12928 35900 12940
rect 35952 12928 35958 12980
rect 36262 12968 36268 12980
rect 36223 12940 36268 12968
rect 36262 12928 36268 12940
rect 36320 12928 36326 12980
rect 37274 12928 37280 12980
rect 37332 12968 37338 12980
rect 37918 12968 37924 12980
rect 37332 12940 37924 12968
rect 37332 12928 37338 12940
rect 37918 12928 37924 12940
rect 37976 12928 37982 12980
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 18322 12900 18328 12912
rect 11664 12872 12434 12900
rect 18283 12872 18328 12900
rect 11664 12860 11670 12872
rect 1627 12804 6960 12832
rect 7101 12835 7159 12841
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 8294 12832 8300 12844
rect 7147 12804 8300 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 9214 12832 9220 12844
rect 9175 12804 9220 12832
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 12158 12832 12164 12844
rect 12119 12804 12164 12832
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12406 12832 12434 12872
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 18417 12903 18475 12909
rect 18417 12869 18429 12903
rect 18463 12900 18475 12903
rect 20070 12900 20076 12912
rect 18463 12872 20076 12900
rect 18463 12869 18475 12872
rect 18417 12863 18475 12869
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 33778 12900 33784 12912
rect 31726 12872 33784 12900
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 12406 12804 14933 12832
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20162 12832 20168 12844
rect 20027 12804 20168 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12832 22983 12835
rect 23474 12832 23480 12844
rect 22971 12804 23480 12832
rect 22971 12801 22983 12804
rect 22925 12795 22983 12801
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 27430 12832 27436 12844
rect 26651 12804 27436 12832
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 29270 12832 29276 12844
rect 29231 12804 29276 12832
rect 29270 12792 29276 12804
rect 29328 12792 29334 12844
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12832 31079 12835
rect 31726 12832 31754 12872
rect 33778 12860 33784 12872
rect 33836 12860 33842 12912
rect 34514 12900 34520 12912
rect 33980 12872 34520 12900
rect 32490 12832 32496 12844
rect 31067 12804 31754 12832
rect 32451 12804 32496 12832
rect 31067 12801 31079 12804
rect 31021 12795 31079 12801
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 33134 12832 33140 12844
rect 33095 12804 33140 12832
rect 33134 12792 33140 12804
rect 33192 12792 33198 12844
rect 33597 12835 33655 12841
rect 33597 12801 33609 12835
rect 33643 12832 33655 12835
rect 33980 12832 34008 12872
rect 34514 12860 34520 12872
rect 34572 12860 34578 12912
rect 34698 12860 34704 12912
rect 34756 12900 34762 12912
rect 37737 12903 37795 12909
rect 37737 12900 37749 12903
rect 34756 12872 37749 12900
rect 34756 12860 34762 12872
rect 37737 12869 37749 12872
rect 37783 12869 37795 12903
rect 37737 12863 37795 12869
rect 33643 12804 34008 12832
rect 33643 12801 33655 12804
rect 33597 12795 33655 12801
rect 34146 12792 34152 12844
rect 34204 12832 34210 12844
rect 34241 12835 34299 12841
rect 34241 12832 34253 12835
rect 34204 12804 34253 12832
rect 34204 12792 34210 12804
rect 34241 12801 34253 12804
rect 34287 12801 34299 12835
rect 34241 12795 34299 12801
rect 34885 12835 34943 12841
rect 34885 12801 34897 12835
rect 34931 12801 34943 12835
rect 34885 12795 34943 12801
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 12434 12764 12440 12776
rect 12391 12736 12440 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 18601 12767 18659 12773
rect 18601 12764 18613 12767
rect 16264 12736 18613 12764
rect 16264 12724 16270 12736
rect 18601 12733 18613 12736
rect 18647 12764 18659 12767
rect 28810 12764 28816 12776
rect 18647 12736 28816 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 28810 12724 28816 12736
rect 28868 12724 28874 12776
rect 34900 12764 34928 12795
rect 34974 12792 34980 12844
rect 35032 12832 35038 12844
rect 35529 12835 35587 12841
rect 35529 12832 35541 12835
rect 35032 12804 35541 12832
rect 35032 12792 35038 12804
rect 35529 12801 35541 12804
rect 35575 12801 35587 12835
rect 35529 12795 35587 12801
rect 36173 12835 36231 12841
rect 36173 12801 36185 12835
rect 36219 12832 36231 12835
rect 36219 12804 37228 12832
rect 36219 12801 36231 12804
rect 36173 12795 36231 12801
rect 36814 12764 36820 12776
rect 34900 12736 36820 12764
rect 36814 12724 36820 12736
rect 36872 12724 36878 12776
rect 31113 12699 31171 12705
rect 31113 12665 31125 12699
rect 31159 12696 31171 12699
rect 33502 12696 33508 12708
rect 31159 12668 33508 12696
rect 31159 12665 31171 12668
rect 31113 12659 31171 12665
rect 33502 12656 33508 12668
rect 33560 12656 33566 12708
rect 33686 12696 33692 12708
rect 33647 12668 33692 12696
rect 33686 12656 33692 12668
rect 33744 12656 33750 12708
rect 37200 12696 37228 12804
rect 37274 12724 37280 12776
rect 37332 12764 37338 12776
rect 37645 12767 37703 12773
rect 37645 12764 37657 12767
rect 37332 12736 37657 12764
rect 37332 12724 37338 12736
rect 37645 12733 37657 12736
rect 37691 12733 37703 12767
rect 37918 12764 37924 12776
rect 37879 12736 37924 12764
rect 37645 12727 37703 12733
rect 37918 12724 37924 12736
rect 37976 12724 37982 12776
rect 38102 12696 38108 12708
rect 37200 12668 38108 12696
rect 38102 12656 38108 12668
rect 38160 12656 38166 12708
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 22741 12631 22799 12637
rect 22741 12597 22753 12631
rect 22787 12628 22799 12631
rect 23014 12628 23020 12640
rect 22787 12600 23020 12628
rect 22787 12597 22799 12600
rect 22741 12591 22799 12597
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 33134 12588 33140 12640
rect 33192 12628 33198 12640
rect 34333 12631 34391 12637
rect 34333 12628 34345 12631
rect 33192 12600 34345 12628
rect 33192 12588 33198 12600
rect 34333 12597 34345 12600
rect 34379 12597 34391 12631
rect 34333 12591 34391 12597
rect 34790 12588 34796 12640
rect 34848 12628 34854 12640
rect 36538 12628 36544 12640
rect 34848 12600 36544 12628
rect 34848 12588 34854 12600
rect 36538 12588 36544 12600
rect 36596 12588 36602 12640
rect 36722 12588 36728 12640
rect 36780 12628 36786 12640
rect 37458 12628 37464 12640
rect 36780 12600 37464 12628
rect 36780 12588 36786 12600
rect 37458 12588 37464 12600
rect 37516 12588 37522 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 20070 12424 20076 12436
rect 20031 12396 20076 12424
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 28261 12427 28319 12433
rect 28261 12393 28273 12427
rect 28307 12424 28319 12427
rect 32858 12424 32864 12436
rect 28307 12396 32864 12424
rect 28307 12393 28319 12396
rect 28261 12387 28319 12393
rect 24946 12316 24952 12368
rect 25004 12356 25010 12368
rect 25004 12328 26234 12356
rect 25004 12316 25010 12328
rect 17586 12288 17592 12300
rect 6886 12260 13492 12288
rect 17547 12260 17592 12288
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 6886 12220 6914 12260
rect 4672 12192 6914 12220
rect 4672 12180 4678 12192
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 13464 12229 13492 12260
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 22554 12248 22560 12300
rect 22612 12288 22618 12300
rect 22649 12291 22707 12297
rect 22649 12288 22661 12291
rect 22612 12260 22661 12288
rect 22612 12248 22618 12260
rect 22649 12257 22661 12260
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 22833 12291 22891 12297
rect 22833 12257 22845 12291
rect 22879 12288 22891 12291
rect 22922 12288 22928 12300
rect 22879 12260 22928 12288
rect 22879 12257 22891 12260
rect 22833 12251 22891 12257
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11664 12192 11989 12220
rect 11664 12180 11670 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 19978 12220 19984 12232
rect 19939 12192 19984 12220
rect 13449 12183 13507 12189
rect 12636 12152 12664 12183
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 16942 12152 16948 12164
rect 11808 12124 12664 12152
rect 16903 12124 16948 12152
rect 11808 12093 11836 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17034 12112 17040 12164
rect 17092 12152 17098 12164
rect 17092 12124 17137 12152
rect 17092 12112 17098 12124
rect 11793 12087 11851 12093
rect 11793 12053 11805 12087
rect 11839 12053 11851 12087
rect 11793 12047 11851 12053
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 22830 12084 22836 12096
rect 13587 12056 22836 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 23293 12087 23351 12093
rect 23293 12084 23305 12087
rect 23164 12056 23305 12084
rect 23164 12044 23170 12056
rect 23293 12053 23305 12056
rect 23339 12053 23351 12087
rect 26206 12084 26234 12328
rect 26789 12291 26847 12297
rect 26789 12257 26801 12291
rect 26835 12288 26847 12291
rect 28276 12288 28304 12387
rect 32858 12384 32864 12396
rect 32916 12384 32922 12436
rect 33410 12424 33416 12436
rect 33371 12396 33416 12424
rect 33410 12384 33416 12396
rect 33468 12384 33474 12436
rect 34238 12424 34244 12436
rect 34199 12396 34244 12424
rect 34238 12384 34244 12396
rect 34296 12384 34302 12436
rect 35345 12427 35403 12433
rect 35345 12393 35357 12427
rect 35391 12424 35403 12427
rect 35710 12424 35716 12436
rect 35391 12396 35716 12424
rect 35391 12393 35403 12396
rect 35345 12387 35403 12393
rect 35710 12384 35716 12396
rect 35768 12384 35774 12436
rect 36633 12427 36691 12433
rect 36633 12393 36645 12427
rect 36679 12424 36691 12427
rect 37090 12424 37096 12436
rect 36679 12396 37096 12424
rect 36679 12393 36691 12396
rect 36633 12387 36691 12393
rect 37090 12384 37096 12396
rect 37148 12384 37154 12436
rect 39114 12424 39120 12436
rect 37200 12396 39120 12424
rect 35897 12359 35955 12365
rect 35897 12325 35909 12359
rect 35943 12356 35955 12359
rect 37200 12356 37228 12396
rect 39114 12384 39120 12396
rect 39172 12384 39178 12436
rect 38378 12356 38384 12368
rect 35943 12328 37228 12356
rect 37292 12328 38384 12356
rect 35943 12325 35955 12328
rect 35897 12319 35955 12325
rect 37292 12297 37320 12328
rect 38378 12316 38384 12328
rect 38436 12356 38442 12368
rect 38838 12356 38844 12368
rect 38436 12328 38844 12356
rect 38436 12316 38442 12328
rect 38838 12316 38844 12328
rect 38896 12316 38902 12368
rect 26835 12260 28304 12288
rect 37277 12291 37335 12297
rect 26835 12257 26847 12260
rect 26789 12251 26847 12257
rect 37277 12257 37289 12291
rect 37323 12257 37335 12291
rect 37550 12288 37556 12300
rect 37511 12260 37556 12288
rect 37277 12251 37335 12257
rect 37550 12248 37556 12260
rect 37608 12248 37614 12300
rect 28169 12223 28227 12229
rect 28169 12189 28181 12223
rect 28215 12220 28227 12223
rect 29822 12220 29828 12232
rect 28215 12192 29828 12220
rect 28215 12189 28227 12192
rect 28169 12183 28227 12189
rect 29822 12180 29828 12192
rect 29880 12180 29886 12232
rect 32306 12180 32312 12232
rect 32364 12220 32370 12232
rect 33321 12223 33379 12229
rect 33321 12220 33333 12223
rect 32364 12192 33333 12220
rect 32364 12180 32370 12192
rect 33321 12189 33333 12192
rect 33367 12189 33379 12223
rect 33321 12183 33379 12189
rect 33594 12180 33600 12232
rect 33652 12220 33658 12232
rect 34149 12223 34207 12229
rect 34149 12220 34161 12223
rect 33652 12192 34161 12220
rect 33652 12180 33658 12192
rect 34149 12189 34161 12192
rect 34195 12220 34207 12223
rect 34422 12220 34428 12232
rect 34195 12192 34428 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 34422 12180 34428 12192
rect 34480 12180 34486 12232
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12220 35311 12223
rect 36078 12220 36084 12232
rect 35299 12192 35894 12220
rect 36039 12192 36084 12220
rect 35299 12189 35311 12192
rect 35253 12183 35311 12189
rect 26878 12112 26884 12164
rect 26936 12152 26942 12164
rect 27433 12155 27491 12161
rect 26936 12124 26981 12152
rect 26936 12112 26942 12124
rect 27433 12121 27445 12155
rect 27479 12121 27491 12155
rect 27433 12115 27491 12121
rect 27448 12084 27476 12115
rect 26206 12056 27476 12084
rect 35866 12084 35894 12192
rect 36078 12180 36084 12192
rect 36136 12180 36142 12232
rect 36538 12220 36544 12232
rect 36499 12192 36544 12220
rect 36538 12180 36544 12192
rect 36596 12180 36602 12232
rect 37090 12112 37096 12164
rect 37148 12152 37154 12164
rect 37369 12155 37427 12161
rect 37369 12152 37381 12155
rect 37148 12124 37381 12152
rect 37148 12112 37154 12124
rect 37369 12121 37381 12124
rect 37415 12121 37427 12155
rect 37369 12115 37427 12121
rect 38746 12084 38752 12096
rect 35866 12056 38752 12084
rect 23293 12047 23351 12053
rect 38746 12044 38752 12056
rect 38804 12044 38810 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 10410 11880 10416 11892
rect 9631 11852 10416 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 16666 11880 16672 11892
rect 14783 11852 16672 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 16816 11852 16957 11880
rect 16816 11840 16822 11852
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 16945 11843 17003 11849
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 19521 11883 19579 11889
rect 19521 11880 19533 11883
rect 17092 11852 19533 11880
rect 17092 11840 17098 11852
rect 19521 11849 19533 11852
rect 19567 11849 19579 11883
rect 19521 11843 19579 11849
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 21048 11852 21465 11880
rect 21048 11840 21054 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 23934 11880 23940 11892
rect 23895 11852 23940 11880
rect 21453 11843 21511 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 34606 11840 34612 11892
rect 34664 11880 34670 11892
rect 34885 11883 34943 11889
rect 34885 11880 34897 11883
rect 34664 11852 34897 11880
rect 34664 11840 34670 11852
rect 34885 11849 34897 11852
rect 34931 11849 34943 11883
rect 35434 11880 35440 11892
rect 35395 11852 35440 11880
rect 34885 11843 34943 11849
rect 35434 11840 35440 11852
rect 35492 11840 35498 11892
rect 37182 11880 37188 11892
rect 35866 11852 37188 11880
rect 25225 11815 25283 11821
rect 25225 11781 25237 11815
rect 25271 11812 25283 11815
rect 26329 11815 26387 11821
rect 26329 11812 26341 11815
rect 25271 11784 26341 11812
rect 25271 11781 25283 11784
rect 25225 11775 25283 11781
rect 26329 11781 26341 11784
rect 26375 11781 26387 11815
rect 35866 11812 35894 11852
rect 37182 11840 37188 11852
rect 37240 11840 37246 11892
rect 37550 11880 37556 11892
rect 37511 11852 37556 11880
rect 37550 11840 37556 11852
rect 37608 11840 37614 11892
rect 36262 11812 36268 11824
rect 26329 11775 26387 11781
rect 33520 11784 35894 11812
rect 36223 11784 36268 11812
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 7616 11716 9505 11744
rect 7616 11704 7622 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14240 11716 14657 11744
rect 14240 11704 14246 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16724 11716 16865 11744
rect 16724 11704 16730 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 16853 11707 16911 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11744 19487 11747
rect 20622 11744 20628 11756
rect 19475 11716 20628 11744
rect 19475 11713 19487 11716
rect 19429 11707 19487 11713
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 17586 11676 17592 11688
rect 15712 11648 17592 11676
rect 15712 11636 15718 11648
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 16390 11568 16396 11620
rect 16448 11608 16454 11620
rect 18800 11608 18828 11707
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 23842 11744 23848 11756
rect 23803 11716 23848 11744
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 26234 11704 26240 11756
rect 26292 11744 26298 11756
rect 26694 11744 26700 11756
rect 26292 11716 26700 11744
rect 26292 11704 26298 11716
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 33520 11753 33548 11784
rect 36262 11772 36268 11784
rect 36320 11772 36326 11824
rect 36354 11772 36360 11824
rect 36412 11812 36418 11824
rect 36412 11784 36457 11812
rect 36412 11772 36418 11784
rect 36538 11772 36544 11824
rect 36596 11812 36602 11824
rect 36596 11784 37504 11812
rect 36596 11772 36602 11784
rect 33505 11747 33563 11753
rect 33505 11713 33517 11747
rect 33551 11713 33563 11747
rect 33505 11707 33563 11713
rect 34054 11704 34060 11756
rect 34112 11744 34118 11756
rect 37476 11753 37504 11784
rect 34333 11747 34391 11753
rect 34333 11744 34345 11747
rect 34112 11716 34345 11744
rect 34112 11704 34118 11716
rect 34333 11713 34345 11716
rect 34379 11744 34391 11747
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 34379 11716 34805 11744
rect 34379 11713 34391 11716
rect 34333 11707 34391 11713
rect 34793 11713 34805 11716
rect 34839 11713 34851 11747
rect 34793 11707 34851 11713
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 37550 11704 37556 11756
rect 37608 11744 37614 11756
rect 38194 11744 38200 11756
rect 37608 11716 38200 11744
rect 37608 11704 37614 11716
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 38289 11747 38347 11753
rect 38289 11713 38301 11747
rect 38335 11713 38347 11747
rect 38289 11707 38347 11713
rect 20806 11676 20812 11688
rect 20767 11648 20812 11676
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20956 11648 21005 11676
rect 20956 11636 20962 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 22738 11676 22744 11688
rect 22699 11648 22744 11676
rect 20993 11639 21051 11645
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 22830 11636 22836 11688
rect 22888 11676 22894 11688
rect 22925 11679 22983 11685
rect 22925 11676 22937 11679
rect 22888 11648 22937 11676
rect 22888 11636 22894 11648
rect 22925 11645 22937 11648
rect 22971 11645 22983 11679
rect 25130 11676 25136 11688
rect 25091 11648 25136 11676
rect 22925 11639 22983 11645
rect 25130 11636 25136 11648
rect 25188 11636 25194 11688
rect 25314 11636 25320 11688
rect 25372 11676 25378 11688
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 25372 11648 25421 11676
rect 25372 11636 25378 11648
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 36740 11648 38148 11676
rect 16448 11580 18828 11608
rect 18877 11611 18935 11617
rect 16448 11568 16454 11580
rect 18877 11577 18889 11611
rect 18923 11608 18935 11611
rect 19610 11608 19616 11620
rect 18923 11580 19616 11608
rect 18923 11577 18935 11580
rect 18877 11571 18935 11577
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 33597 11611 33655 11617
rect 33597 11577 33609 11611
rect 33643 11608 33655 11611
rect 33643 11580 35020 11608
rect 33643 11577 33655 11580
rect 33597 11571 33655 11577
rect 17586 11540 17592 11552
rect 17547 11512 17592 11540
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 23106 11540 23112 11552
rect 23067 11512 23112 11540
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 34149 11543 34207 11549
rect 34149 11509 34161 11543
rect 34195 11540 34207 11543
rect 34330 11540 34336 11552
rect 34195 11512 34336 11540
rect 34195 11509 34207 11512
rect 34149 11503 34207 11509
rect 34330 11500 34336 11512
rect 34388 11500 34394 11552
rect 34992 11540 35020 11580
rect 35618 11568 35624 11620
rect 35676 11608 35682 11620
rect 36740 11608 36768 11648
rect 35676 11580 36768 11608
rect 36817 11611 36875 11617
rect 35676 11568 35682 11580
rect 36817 11577 36829 11611
rect 36863 11608 36875 11611
rect 37550 11608 37556 11620
rect 36863 11580 37556 11608
rect 36863 11577 36875 11580
rect 36817 11571 36875 11577
rect 37550 11568 37556 11580
rect 37608 11568 37614 11620
rect 38120 11617 38148 11648
rect 38105 11611 38163 11617
rect 38105 11577 38117 11611
rect 38151 11577 38163 11611
rect 38105 11571 38163 11577
rect 36722 11540 36728 11552
rect 34992 11512 36728 11540
rect 36722 11500 36728 11512
rect 36780 11500 36786 11552
rect 36906 11500 36912 11552
rect 36964 11540 36970 11552
rect 38304 11540 38332 11707
rect 36964 11512 38332 11540
rect 36964 11500 36970 11512
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17184 11308 17417 11336
rect 17184 11296 17190 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 17405 11299 17463 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 34149 11339 34207 11345
rect 34149 11305 34161 11339
rect 34195 11336 34207 11339
rect 34698 11336 34704 11348
rect 34195 11308 34704 11336
rect 34195 11305 34207 11308
rect 34149 11299 34207 11305
rect 34698 11296 34704 11308
rect 34756 11296 34762 11348
rect 36262 11296 36268 11348
rect 36320 11336 36326 11348
rect 36725 11339 36783 11345
rect 36725 11336 36737 11339
rect 36320 11308 36737 11336
rect 36320 11296 36326 11308
rect 36725 11305 36737 11308
rect 36771 11305 36783 11339
rect 36725 11299 36783 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 9490 11268 9496 11280
rect 1627 11240 9496 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 35345 11271 35403 11277
rect 35345 11237 35357 11271
rect 35391 11268 35403 11271
rect 36078 11268 36084 11280
rect 35391 11240 36084 11268
rect 35391 11237 35403 11240
rect 35345 11231 35403 11237
rect 36078 11228 36084 11240
rect 36136 11228 36142 11280
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 16942 11200 16948 11212
rect 9263 11172 16948 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 17644 11172 19533 11200
rect 17644 11160 17650 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 21085 11203 21143 11209
rect 21085 11200 21097 11203
rect 20864 11172 21097 11200
rect 20864 11160 20870 11172
rect 21085 11169 21097 11172
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 28810 11160 28816 11212
rect 28868 11200 28874 11212
rect 29181 11203 29239 11209
rect 29181 11200 29193 11203
rect 28868 11172 29193 11200
rect 28868 11160 28874 11172
rect 29181 11169 29193 11172
rect 29227 11200 29239 11203
rect 31662 11200 31668 11212
rect 29227 11172 31668 11200
rect 29227 11169 29239 11172
rect 29181 11163 29239 11169
rect 31662 11160 31668 11172
rect 31720 11160 31726 11212
rect 33870 11160 33876 11212
rect 33928 11200 33934 11212
rect 33928 11172 35894 11200
rect 33928 11160 33934 11172
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 7708 11104 9137 11132
rect 7708 11092 7714 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 16390 11132 16396 11144
rect 16351 11104 16396 11132
rect 9125 11095 9183 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 21913 11135 21971 11141
rect 21913 11132 21925 11135
rect 21600 11104 21925 11132
rect 21600 11092 21606 11104
rect 21913 11101 21925 11104
rect 21959 11101 21971 11135
rect 23014 11132 23020 11144
rect 22975 11104 23020 11132
rect 21913 11095 21971 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 31846 11132 31852 11144
rect 29104 11104 31852 11132
rect 16485 11067 16543 11073
rect 16485 11033 16497 11067
rect 16531 11064 16543 11067
rect 17034 11064 17040 11076
rect 16531 11036 17040 11064
rect 16531 11033 16543 11036
rect 16485 11027 16543 11033
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 20165 11067 20223 11073
rect 19668 11036 19713 11064
rect 19668 11024 19674 11036
rect 20165 11033 20177 11067
rect 20211 11064 20223 11067
rect 24946 11064 24952 11076
rect 20211 11036 24952 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 24946 11024 24952 11036
rect 25004 11024 25010 11076
rect 25406 11024 25412 11076
rect 25464 11064 25470 11076
rect 28169 11067 28227 11073
rect 28169 11064 28181 11067
rect 25464 11036 28181 11064
rect 25464 11024 25470 11036
rect 28169 11033 28181 11036
rect 28215 11033 28227 11067
rect 28169 11027 28227 11033
rect 28261 11067 28319 11073
rect 28261 11033 28273 11067
rect 28307 11064 28319 11067
rect 29104 11064 29132 11104
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 32030 11132 32036 11144
rect 31991 11104 32036 11132
rect 32030 11092 32036 11104
rect 32088 11092 32094 11144
rect 34330 11132 34336 11144
rect 34291 11104 34336 11132
rect 34330 11092 34336 11104
rect 34388 11092 34394 11144
rect 34422 11092 34428 11144
rect 34480 11132 34486 11144
rect 35529 11135 35587 11141
rect 35529 11132 35541 11135
rect 34480 11104 35541 11132
rect 34480 11092 34486 11104
rect 35529 11101 35541 11104
rect 35575 11101 35587 11135
rect 35866 11132 35894 11172
rect 37642 11160 37648 11212
rect 37700 11200 37706 11212
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37700 11172 37749 11200
rect 37700 11160 37706 11172
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 35989 11135 36047 11141
rect 35989 11132 36001 11135
rect 35866 11104 36001 11132
rect 35529 11095 35587 11101
rect 35989 11101 36001 11104
rect 36035 11101 36047 11135
rect 35989 11095 36047 11101
rect 36538 11092 36544 11144
rect 36596 11132 36602 11144
rect 36633 11135 36691 11141
rect 36633 11132 36645 11135
rect 36596 11104 36645 11132
rect 36596 11092 36602 11104
rect 36633 11101 36645 11104
rect 36679 11101 36691 11135
rect 36633 11095 36691 11101
rect 28307 11036 29132 11064
rect 32125 11067 32183 11073
rect 28307 11033 28319 11036
rect 28261 11027 28319 11033
rect 32125 11033 32137 11067
rect 32171 11064 32183 11067
rect 32490 11064 32496 11076
rect 32171 11036 32496 11064
rect 32171 11033 32183 11036
rect 32125 11027 32183 11033
rect 32490 11024 32496 11036
rect 32548 11024 32554 11076
rect 36081 11067 36139 11073
rect 36081 11033 36093 11067
rect 36127 11064 36139 11067
rect 37734 11064 37740 11076
rect 36127 11036 37740 11064
rect 36127 11033 36139 11036
rect 36081 11027 36139 11033
rect 37734 11024 37740 11036
rect 37792 11024 37798 11076
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 21729 10999 21787 11005
rect 21729 10996 21741 10999
rect 21048 10968 21741 10996
rect 21048 10956 21054 10968
rect 21729 10965 21741 10968
rect 21775 10965 21787 10999
rect 21729 10959 21787 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 8754 10792 8760 10804
rect 1627 10764 8760 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 20809 10795 20867 10801
rect 20809 10761 20821 10795
rect 20855 10792 20867 10795
rect 20898 10792 20904 10804
rect 20855 10764 20904 10792
rect 20855 10761 20867 10764
rect 20809 10755 20867 10761
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 32398 10752 32404 10804
rect 32456 10792 32462 10804
rect 32585 10795 32643 10801
rect 32585 10792 32597 10795
rect 32456 10764 32597 10792
rect 32456 10752 32462 10764
rect 32585 10761 32597 10764
rect 32631 10761 32643 10795
rect 32585 10755 32643 10761
rect 35897 10795 35955 10801
rect 35897 10761 35909 10795
rect 35943 10792 35955 10795
rect 35986 10792 35992 10804
rect 35943 10764 35992 10792
rect 35943 10761 35955 10764
rect 35897 10755 35955 10761
rect 35986 10752 35992 10764
rect 36044 10752 36050 10804
rect 36633 10795 36691 10801
rect 36633 10761 36645 10795
rect 36679 10792 36691 10795
rect 37366 10792 37372 10804
rect 36679 10764 37372 10792
rect 36679 10761 36691 10764
rect 36633 10755 36691 10761
rect 37366 10752 37372 10764
rect 37424 10752 37430 10804
rect 12989 10727 13047 10733
rect 12989 10693 13001 10727
rect 13035 10724 13047 10727
rect 13722 10724 13728 10736
rect 13035 10696 13728 10724
rect 13035 10693 13047 10696
rect 12989 10687 13047 10693
rect 13722 10684 13728 10696
rect 13780 10684 13786 10736
rect 17034 10724 17040 10736
rect 16995 10696 17040 10724
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 17589 10727 17647 10733
rect 17589 10693 17601 10727
rect 17635 10724 17647 10727
rect 25314 10724 25320 10736
rect 17635 10696 25320 10724
rect 17635 10693 17647 10696
rect 17589 10687 17647 10693
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 34517 10727 34575 10733
rect 34517 10693 34529 10727
rect 34563 10724 34575 10727
rect 36354 10724 36360 10736
rect 34563 10696 36360 10724
rect 34563 10693 34575 10696
rect 34517 10687 34575 10693
rect 36354 10684 36360 10696
rect 36412 10684 36418 10736
rect 38470 10724 38476 10736
rect 36556 10696 38476 10724
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10656 25099 10659
rect 26234 10656 26240 10668
rect 25087 10628 26240 10656
rect 25087 10625 25099 10628
rect 25041 10619 25099 10625
rect 26234 10616 26240 10628
rect 26292 10616 26298 10668
rect 28813 10659 28871 10665
rect 28813 10625 28825 10659
rect 28859 10656 28871 10659
rect 28902 10656 28908 10668
rect 28859 10628 28908 10656
rect 28859 10625 28871 10628
rect 28813 10619 28871 10625
rect 28902 10616 28908 10628
rect 28960 10616 28966 10668
rect 32493 10659 32551 10665
rect 32493 10625 32505 10659
rect 32539 10625 32551 10659
rect 34422 10656 34428 10668
rect 34383 10628 34428 10656
rect 32493 10619 32551 10625
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 11020 10560 12909 10588
rect 11020 10548 11026 10560
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 13446 10588 13452 10600
rect 13407 10560 13452 10588
rect 12897 10551 12955 10557
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 13722 10588 13728 10600
rect 13504 10560 13728 10588
rect 13504 10548 13510 10560
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 16942 10588 16948 10600
rect 16903 10560 16948 10588
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 24397 10591 24455 10597
rect 24397 10557 24409 10591
rect 24443 10588 24455 10591
rect 24670 10588 24676 10600
rect 24443 10560 24676 10588
rect 24443 10557 24455 10560
rect 24397 10551 24455 10557
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 27798 10548 27804 10600
rect 27856 10588 27862 10600
rect 32508 10588 32536 10619
rect 34422 10616 34428 10628
rect 34480 10616 34486 10668
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10625 35311 10659
rect 36078 10656 36084 10668
rect 36039 10628 36084 10656
rect 35253 10619 35311 10625
rect 27856 10560 32536 10588
rect 27856 10548 27862 10560
rect 35268 10520 35296 10619
rect 36078 10616 36084 10628
rect 36136 10616 36142 10668
rect 36556 10665 36584 10696
rect 38470 10684 38476 10696
rect 38528 10684 38534 10736
rect 36541 10659 36599 10665
rect 36541 10625 36553 10659
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 37458 10616 37464 10668
rect 37516 10656 37522 10668
rect 38013 10659 38071 10665
rect 38013 10656 38025 10659
rect 37516 10628 38025 10656
rect 37516 10616 37522 10628
rect 38013 10625 38025 10628
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 35345 10591 35403 10597
rect 35345 10557 35357 10591
rect 35391 10588 35403 10591
rect 38378 10588 38384 10600
rect 35391 10560 38384 10588
rect 35391 10557 35403 10560
rect 35345 10551 35403 10557
rect 38378 10548 38384 10560
rect 38436 10548 38442 10600
rect 37734 10520 37740 10532
rect 35268 10492 37740 10520
rect 37734 10480 37740 10492
rect 37792 10480 37798 10532
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 25133 10455 25191 10461
rect 25133 10452 25145 10455
rect 24820 10424 25145 10452
rect 24820 10412 24826 10424
rect 25133 10421 25145 10424
rect 25179 10421 25191 10455
rect 25133 10415 25191 10421
rect 28905 10455 28963 10461
rect 28905 10421 28917 10455
rect 28951 10452 28963 10455
rect 28994 10452 29000 10464
rect 28951 10424 29000 10452
rect 28951 10421 28963 10424
rect 28905 10415 28963 10421
rect 28994 10412 29000 10424
rect 29052 10412 29058 10464
rect 38194 10452 38200 10464
rect 38155 10424 38200 10452
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 10134 10248 10140 10260
rect 7975 10220 10140 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 25866 10248 25872 10260
rect 25827 10220 25872 10248
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 36722 10248 36728 10260
rect 36683 10220 36728 10248
rect 36722 10208 36728 10220
rect 36780 10208 36786 10260
rect 24854 10180 24860 10192
rect 19720 10152 24860 10180
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7248 10016 7849 10044
rect 7248 10004 7254 10016
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 7837 10007 7895 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 19720 10053 19748 10152
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 35526 10140 35532 10192
rect 35584 10180 35590 10192
rect 37829 10183 37887 10189
rect 37829 10180 37841 10183
rect 35584 10152 37841 10180
rect 35584 10140 35590 10152
rect 37829 10149 37841 10152
rect 37875 10149 37887 10183
rect 37829 10143 37887 10149
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 23106 10112 23112 10124
rect 21775 10084 23112 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 24670 10112 24676 10124
rect 24631 10084 24676 10112
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 24946 10112 24952 10124
rect 24907 10084 24952 10112
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22094 10044 22100 10056
rect 21959 10016 22100 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10013 25835 10047
rect 36170 10044 36176 10056
rect 36131 10016 36176 10044
rect 25777 10007 25835 10013
rect 24762 9976 24768 9988
rect 24723 9948 24768 9976
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 9585 9911 9643 9917
rect 9585 9877 9597 9911
rect 9631 9908 9643 9911
rect 16942 9908 16948 9920
rect 9631 9880 16948 9908
rect 9631 9877 9643 9880
rect 9585 9871 9643 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19484 9880 19809 9908
rect 19484 9868 19490 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 20806 9868 20812 9920
rect 20864 9908 20870 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20864 9880 21005 9908
rect 20864 9868 20870 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 22370 9908 22376 9920
rect 22331 9880 22376 9908
rect 20993 9871 21051 9877
rect 22370 9868 22376 9880
rect 22428 9868 22434 9920
rect 24578 9868 24584 9920
rect 24636 9908 24642 9920
rect 25792 9908 25820 10007
rect 36170 10004 36176 10016
rect 36228 10004 36234 10056
rect 36630 10044 36636 10056
rect 36591 10016 36636 10044
rect 36630 10004 36636 10016
rect 36688 10004 36694 10056
rect 37550 10004 37556 10056
rect 37608 10044 37614 10056
rect 37737 10047 37795 10053
rect 37737 10044 37749 10047
rect 37608 10016 37749 10044
rect 37608 10004 37614 10016
rect 37737 10013 37749 10016
rect 37783 10013 37795 10047
rect 37737 10007 37795 10013
rect 35986 9908 35992 9920
rect 24636 9880 25820 9908
rect 35947 9880 35992 9908
rect 24636 9868 24642 9880
rect 35986 9868 35992 9880
rect 36044 9868 36050 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 9048 9676 9444 9704
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 8846 9636 8852 9648
rect 4847 9608 8852 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 9048 9636 9076 9676
rect 8956 9608 9076 9636
rect 9125 9639 9183 9645
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 8956 9568 8984 9608
rect 9125 9605 9137 9639
rect 9171 9636 9183 9639
rect 9306 9636 9312 9648
rect 9171 9608 9312 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 9416 9636 9444 9676
rect 13354 9636 13360 9648
rect 9416 9608 13360 9636
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 22094 9636 22100 9648
rect 19392 9608 20944 9636
rect 22055 9608 22100 9636
rect 19392 9596 19398 9608
rect 6963 9540 8984 9568
rect 9033 9571 9091 9577
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 9048 9500 9076 9531
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 18969 9571 19027 9577
rect 18969 9568 18981 9571
rect 17092 9540 18981 9568
rect 17092 9528 17098 9540
rect 18969 9537 18981 9540
rect 19015 9537 19027 9571
rect 20806 9568 20812 9580
rect 20767 9540 20812 9568
rect 18969 9531 19027 9537
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20916 9568 20944 9608
rect 22094 9596 22100 9608
rect 22152 9596 22158 9648
rect 25406 9636 25412 9648
rect 25367 9608 25412 9636
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 30374 9636 30380 9648
rect 30335 9608 30380 9636
rect 30374 9596 30380 9608
rect 30432 9596 30438 9648
rect 31297 9639 31355 9645
rect 31297 9605 31309 9639
rect 31343 9636 31355 9639
rect 36446 9636 36452 9648
rect 31343 9608 36452 9636
rect 31343 9605 31355 9608
rect 31297 9599 31355 9605
rect 36446 9596 36452 9608
rect 36504 9596 36510 9648
rect 36725 9639 36783 9645
rect 36725 9605 36737 9639
rect 36771 9636 36783 9639
rect 37274 9636 37280 9648
rect 36771 9608 37280 9636
rect 36771 9605 36783 9608
rect 36725 9599 36783 9605
rect 37274 9596 37280 9608
rect 37332 9596 37338 9648
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 20916 9540 22017 9568
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 23474 9528 23480 9580
rect 23532 9568 23538 9580
rect 25317 9571 25375 9577
rect 25317 9568 25329 9571
rect 23532 9540 25329 9568
rect 23532 9528 23538 9540
rect 25317 9537 25329 9540
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27212 9540 27445 9568
rect 27212 9528 27218 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 37734 9528 37740 9580
rect 37792 9568 37798 9580
rect 38013 9571 38071 9577
rect 38013 9568 38025 9571
rect 37792 9540 38025 9568
rect 37792 9528 37798 9540
rect 38013 9537 38025 9540
rect 38059 9568 38071 9571
rect 39666 9568 39672 9580
rect 38059 9540 39672 9568
rect 38059 9537 38071 9540
rect 38013 9531 38071 9537
rect 39666 9528 39672 9540
rect 39724 9528 39730 9580
rect 5868 9472 9076 9500
rect 5868 9460 5874 9472
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20496 9472 21005 9500
rect 20496 9460 20502 9472
rect 20993 9469 21005 9472
rect 21039 9469 21051 9503
rect 30285 9503 30343 9509
rect 30285 9500 30297 9503
rect 20993 9463 21051 9469
rect 26206 9472 30297 9500
rect 19061 9435 19119 9441
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 22738 9432 22744 9444
rect 19107 9404 22744 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 22738 9392 22744 9404
rect 22796 9432 22802 9444
rect 26206 9432 26234 9472
rect 30285 9469 30297 9472
rect 30331 9469 30343 9503
rect 30285 9463 30343 9469
rect 37826 9432 37832 9444
rect 22796 9404 26234 9432
rect 37787 9404 37832 9432
rect 22796 9392 22802 9404
rect 37826 9392 37832 9404
rect 37884 9392 37890 9444
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7098 9364 7104 9376
rect 7055 9336 7104 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 19944 9336 21189 9364
rect 19944 9324 19950 9336
rect 21177 9333 21189 9336
rect 21223 9364 21235 9367
rect 22370 9364 22376 9376
rect 21223 9336 22376 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 27525 9367 27583 9373
rect 27525 9333 27537 9367
rect 27571 9364 27583 9367
rect 28074 9364 28080 9376
rect 27571 9336 28080 9364
rect 27571 9333 27583 9336
rect 27525 9327 27583 9333
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 20438 9160 20444 9172
rect 20399 9132 20444 9160
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19392 8996 20024 9024
rect 19392 8984 19398 8996
rect 1762 8956 1768 8968
rect 1723 8928 1768 8956
rect 1762 8916 1768 8928
rect 1820 8916 1826 8968
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 19886 8956 19892 8968
rect 18739 8928 19892 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 19996 8965 20024 8996
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8925 20039 8959
rect 19981 8919 20039 8925
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8925 20683 8959
rect 28074 8956 28080 8968
rect 28035 8928 28080 8956
rect 20625 8919 20683 8925
rect 20640 8888 20668 8919
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 19812 8860 20668 8888
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19812 8829 19840 8860
rect 19797 8823 19855 8829
rect 19797 8789 19809 8823
rect 19843 8789 19855 8823
rect 19797 8783 19855 8789
rect 27893 8823 27951 8829
rect 27893 8789 27905 8823
rect 27939 8820 27951 8823
rect 30374 8820 30380 8832
rect 27939 8792 30380 8820
rect 27939 8789 27951 8792
rect 27893 8783 27951 8789
rect 30374 8780 30380 8792
rect 30432 8780 30438 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 18046 8576 18052 8628
rect 18104 8616 18110 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 18104 8588 19257 8616
rect 18104 8576 18110 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 19245 8579 19303 8585
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25188 8588 25237 8616
rect 25188 8576 25194 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 38102 8616 38108 8628
rect 38063 8588 38108 8616
rect 25225 8579 25283 8585
rect 38102 8576 38108 8588
rect 38160 8576 38166 8628
rect 38746 8548 38752 8560
rect 37660 8520 38752 8548
rect 7098 8480 7104 8492
rect 7059 8452 7104 8480
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 19426 8480 19432 8492
rect 19387 8452 19432 8480
rect 9217 8443 9275 8449
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 9232 8412 9260 8443
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 25130 8480 25136 8492
rect 25091 8452 25136 8480
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 37660 8489 37688 8520
rect 38746 8508 38752 8520
rect 38804 8508 38810 8560
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 38286 8480 38292 8492
rect 38247 8452 38292 8480
rect 37645 8443 37703 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 5684 8384 9260 8412
rect 5684 8372 5690 8384
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 5776 8316 6929 8344
rect 5776 8304 5782 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 9309 8347 9367 8353
rect 9309 8313 9321 8347
rect 9355 8344 9367 8347
rect 27246 8344 27252 8356
rect 9355 8316 27252 8344
rect 9355 8313 9367 8316
rect 9309 8307 9367 8313
rect 27246 8304 27252 8316
rect 27304 8304 27310 8356
rect 36630 8304 36636 8356
rect 36688 8344 36694 8356
rect 37461 8347 37519 8353
rect 37461 8344 37473 8347
rect 36688 8316 37473 8344
rect 36688 8304 36694 8316
rect 37461 8313 37473 8316
rect 37507 8313 37519 8347
rect 37461 8307 37519 8313
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 10962 8072 10968 8084
rect 10923 8044 10968 8072
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 1596 7908 2237 7936
rect 1596 7877 1624 7908
rect 2225 7905 2237 7908
rect 2271 7936 2283 7939
rect 20346 7936 20352 7948
rect 2271 7908 20352 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 20346 7896 20352 7908
rect 20404 7896 20410 7948
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 6972 7840 10885 7868
rect 6972 7828 6978 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 25038 7828 25044 7880
rect 25096 7868 25102 7880
rect 28994 7868 29000 7880
rect 25096 7840 26234 7868
rect 28955 7840 29000 7868
rect 25096 7828 25102 7840
rect 26206 7800 26234 7840
rect 28994 7828 29000 7840
rect 29052 7828 29058 7880
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 35866 7840 38025 7868
rect 35866 7800 35894 7840
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 26206 7772 35894 7800
rect 1762 7732 1768 7744
rect 1723 7704 1768 7732
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 28813 7735 28871 7741
rect 28813 7701 28825 7735
rect 28859 7732 28871 7735
rect 30006 7732 30012 7744
rect 28859 7704 30012 7732
rect 28859 7701 28871 7704
rect 28813 7695 28871 7701
rect 30006 7692 30012 7704
rect 30064 7692 30070 7744
rect 38194 7732 38200 7744
rect 38155 7704 38200 7732
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 32766 7488 32772 7540
rect 32824 7528 32830 7540
rect 38105 7531 38163 7537
rect 38105 7528 38117 7531
rect 32824 7500 38117 7528
rect 32824 7488 32830 7500
rect 38105 7497 38117 7500
rect 38151 7497 38163 7531
rect 38105 7491 38163 7497
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1728 7364 1869 7392
rect 1728 7352 1734 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 18782 7392 18788 7404
rect 17819 7364 18788 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 33134 7392 33140 7404
rect 33095 7364 33140 7392
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 14918 7148 14924 7200
rect 14976 7188 14982 7200
rect 17589 7191 17647 7197
rect 17589 7188 17601 7191
rect 14976 7160 17601 7188
rect 14976 7148 14982 7160
rect 17589 7157 17601 7160
rect 17635 7157 17647 7191
rect 17589 7151 17647 7157
rect 32953 7191 33011 7197
rect 32953 7157 32965 7191
rect 32999 7188 33011 7191
rect 34422 7188 34428 7200
rect 32999 7160 34428 7188
rect 32999 7157 33011 7160
rect 32953 7151 33011 7157
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8386 6304 8392 6316
rect 7975 6276 8392 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 5592 6072 7757 6100
rect 5592 6060 5598 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 8386 5896 8392 5908
rect 8347 5868 8392 5896
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 1946 5760 1952 5772
rect 1903 5732 1952 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 13630 5692 13636 5704
rect 8343 5664 13636 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 29822 5652 29828 5704
rect 29880 5692 29886 5704
rect 29917 5695 29975 5701
rect 29917 5692 29929 5695
rect 29880 5664 29929 5692
rect 29880 5652 29886 5664
rect 29917 5661 29929 5664
rect 29963 5661 29975 5695
rect 38013 5695 38071 5701
rect 38013 5692 38025 5695
rect 29917 5655 29975 5661
rect 35866 5664 38025 5692
rect 29733 5559 29791 5565
rect 29733 5525 29745 5559
rect 29779 5556 29791 5559
rect 35866 5556 35894 5664
rect 38013 5661 38025 5664
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 38194 5556 38200 5568
rect 29779 5528 35894 5556
rect 38155 5528 38200 5556
rect 29779 5525 29791 5528
rect 29733 5519 29791 5525
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 7650 4808 7656 4820
rect 1627 4780 7656 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 1762 4604 1768 4616
rect 1723 4576 1768 4604
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 32490 4564 32496 4616
rect 32548 4604 32554 4616
rect 32585 4607 32643 4613
rect 32585 4604 32597 4607
rect 32548 4576 32597 4604
rect 32548 4564 32554 4576
rect 32585 4573 32597 4576
rect 32631 4573 32643 4607
rect 38286 4604 38292 4616
rect 38247 4576 38292 4604
rect 32585 4567 32643 4573
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 32401 4471 32459 4477
rect 32401 4437 32413 4471
rect 32447 4468 32459 4471
rect 35342 4468 35348 4480
rect 32447 4440 35348 4468
rect 32447 4437 32459 4440
rect 32401 4431 32459 4437
rect 35342 4428 35348 4440
rect 35400 4428 35406 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 658 4088 664 4140
rect 716 4128 722 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 716 4100 1777 4128
rect 716 4088 722 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 36446 4088 36452 4140
rect 36504 4128 36510 4140
rect 36725 4131 36783 4137
rect 36725 4128 36737 4131
rect 36504 4100 36737 4128
rect 36504 4088 36510 4100
rect 36725 4097 36737 4100
rect 36771 4097 36783 4131
rect 38010 4128 38016 4140
rect 37971 4100 38016 4128
rect 36725 4091 36783 4097
rect 38010 4088 38016 4100
rect 38068 4088 38074 4140
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 7558 3992 7564 4004
rect 1627 3964 7564 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 36817 3927 36875 3933
rect 36817 3893 36829 3927
rect 36863 3924 36875 3927
rect 36906 3924 36912 3936
rect 36863 3896 36912 3924
rect 36863 3893 36875 3896
rect 36817 3887 36875 3893
rect 36906 3884 36912 3896
rect 36964 3884 36970 3936
rect 38194 3924 38200 3936
rect 38155 3896 38200 3924
rect 38194 3884 38200 3896
rect 38252 3884 38258 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 5626 3720 5632 3732
rect 2363 3692 5632 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 33778 3680 33784 3732
rect 33836 3720 33842 3732
rect 36817 3723 36875 3729
rect 36817 3720 36829 3723
rect 33836 3692 36829 3720
rect 33836 3680 33842 3692
rect 36817 3689 36829 3692
rect 36863 3689 36875 3723
rect 36817 3683 36875 3689
rect 5718 3584 5724 3596
rect 1596 3556 5724 3584
rect 1596 3525 1624 3556
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 28626 3544 28632 3596
rect 28684 3584 28690 3596
rect 37737 3587 37795 3593
rect 37737 3584 37749 3587
rect 28684 3556 37749 3584
rect 28684 3544 28690 3556
rect 37737 3553 37749 3556
rect 37783 3553 37795 3587
rect 37737 3547 37795 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 37001 3519 37059 3525
rect 37001 3485 37013 3519
rect 37047 3485 37059 3519
rect 37458 3516 37464 3528
rect 37419 3488 37464 3516
rect 37001 3479 37059 3485
rect 14 3408 20 3460
rect 72 3448 78 3460
rect 2516 3448 2544 3479
rect 72 3420 2544 3448
rect 72 3408 78 3420
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 34514 3448 34520 3460
rect 17920 3420 34520 3448
rect 17920 3408 17926 3420
rect 34514 3408 34520 3420
rect 34572 3408 34578 3460
rect 37016 3448 37044 3479
rect 37458 3476 37464 3488
rect 37516 3476 37522 3528
rect 38654 3448 38660 3460
rect 37016 3420 38660 3448
rect 38654 3408 38660 3420
rect 38712 3408 38718 3460
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 35529 3179 35587 3185
rect 35529 3145 35541 3179
rect 35575 3145 35587 3179
rect 35529 3139 35587 3145
rect 36725 3179 36783 3185
rect 36725 3145 36737 3179
rect 36771 3176 36783 3179
rect 38010 3176 38016 3188
rect 36771 3148 38016 3176
rect 36771 3145 36783 3148
rect 36725 3139 36783 3145
rect 13722 3108 13728 3120
rect 2148 3080 13728 3108
rect 2148 3049 2176 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 17310 3108 17316 3120
rect 16546 3080 17316 3108
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2271 3012 2881 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3040 4031 3043
rect 5534 3040 5540 3052
rect 4019 3012 5540 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16546 3040 16574 3080
rect 17310 3068 17316 3080
rect 17368 3108 17374 3120
rect 17862 3108 17868 3120
rect 17368 3080 17868 3108
rect 17368 3068 17374 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 17034 3040 17040 3052
rect 16347 3012 16574 3040
rect 16995 3012 17040 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 33045 3043 33103 3049
rect 33045 3009 33057 3043
rect 33091 3040 33103 3043
rect 35544 3040 35572 3139
rect 38010 3136 38016 3148
rect 38068 3136 38074 3188
rect 33091 3012 35572 3040
rect 35713 3043 35771 3049
rect 33091 3009 33103 3012
rect 33045 3003 33103 3009
rect 35713 3009 35725 3043
rect 35759 3009 35771 3043
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 35713 3003 35771 3009
rect 35434 2932 35440 2984
rect 35492 2972 35498 2984
rect 35728 2972 35756 3003
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 37461 3043 37519 3049
rect 37461 3009 37473 3043
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 35492 2944 35756 2972
rect 35492 2932 35498 2944
rect 34422 2864 34428 2916
rect 34480 2904 34486 2916
rect 37476 2904 37504 3003
rect 34480 2876 37504 2904
rect 34480 2864 34486 2876
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 1636 2808 2697 2836
rect 1636 2796 1642 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 3936 2808 4169 2836
rect 3936 2796 3942 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 16114 2836 16120 2848
rect 16075 2808 16120 2836
rect 4157 2799 4215 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16816 2808 16865 2836
rect 16816 2796 16822 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 32861 2839 32919 2845
rect 32861 2836 32873 2839
rect 32364 2808 32873 2836
rect 32364 2796 32370 2808
rect 32861 2805 32873 2808
rect 32907 2805 32919 2839
rect 32861 2799 32919 2805
rect 37366 2796 37372 2848
rect 37424 2836 37430 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37424 2808 37657 2836
rect 37424 2796 37430 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 37645 2799 37703 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 4706 2632 4712 2644
rect 3007 2604 4712 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5810 2632 5816 2644
rect 4816 2604 5816 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 4816 2564 4844 2604
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6914 2632 6920 2644
rect 6595 2604 6920 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7190 2632 7196 2644
rect 7151 2604 7196 2632
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 14182 2632 14188 2644
rect 8435 2604 14188 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 16666 2632 16672 2644
rect 14323 2604 16672 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 19429 2635 19487 2641
rect 19429 2601 19441 2635
rect 19475 2632 19487 2635
rect 20162 2632 20168 2644
rect 19475 2604 20168 2632
rect 19475 2601 19487 2604
rect 19429 2595 19487 2601
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20303 2635 20361 2641
rect 20303 2601 20315 2635
rect 20349 2632 20361 2635
rect 23106 2632 23112 2644
rect 20349 2604 23112 2632
rect 20349 2601 20361 2604
rect 20303 2595 20361 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23293 2635 23351 2641
rect 23293 2601 23305 2635
rect 23339 2632 23351 2635
rect 23842 2632 23848 2644
rect 23339 2604 23848 2632
rect 23339 2601 23351 2604
rect 23293 2595 23351 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 24578 2632 24584 2644
rect 24539 2604 24584 2632
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 28776 2604 29745 2632
rect 28776 2592 28782 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 29733 2595 29791 2601
rect 34514 2592 34520 2644
rect 34572 2632 34578 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34572 2604 35081 2632
rect 34572 2592 34578 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 2363 2536 4844 2564
rect 5261 2567 5319 2573
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 5261 2533 5273 2567
rect 5307 2564 5319 2567
rect 9214 2564 9220 2576
rect 5307 2536 9220 2564
rect 5307 2533 5319 2536
rect 5261 2527 5319 2533
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 16114 2564 16120 2576
rect 9600 2536 16120 2564
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2004 2400 2513 2428
rect 2004 2388 2010 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 2501 2391 2559 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3292 2400 3985 2428
rect 3292 2388 3298 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 9600 2437 9628 2536
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 20530 2564 20536 2576
rect 16546 2536 20536 2564
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 16546 2496 16574 2536
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 22005 2567 22063 2573
rect 22005 2533 22017 2567
rect 22051 2564 22063 2567
rect 23474 2564 23480 2576
rect 22051 2536 23480 2564
rect 22051 2533 22063 2536
rect 22005 2527 22063 2533
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 27157 2567 27215 2573
rect 27157 2533 27169 2567
rect 27203 2564 27215 2567
rect 29270 2564 29276 2576
rect 27203 2536 29276 2564
rect 27203 2533 27215 2536
rect 27157 2527 27215 2533
rect 29270 2524 29276 2536
rect 29328 2524 29334 2576
rect 36081 2567 36139 2573
rect 36081 2533 36093 2567
rect 36127 2564 36139 2567
rect 37182 2564 37188 2576
rect 36127 2536 37188 2564
rect 36127 2533 36139 2536
rect 36081 2527 36139 2533
rect 37182 2524 37188 2536
rect 37240 2524 37246 2576
rect 21174 2496 21180 2508
rect 10643 2468 16574 2496
rect 18156 2468 21180 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8444 2400 8585 2428
rect 8444 2388 8450 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 9585 2391 9643 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 11992 2360 12020 2391
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12952 2400 13185 2428
rect 12952 2388 12958 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13596 2400 14473 2428
rect 13596 2388 13602 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 14461 2391 14519 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16758 2428 16764 2440
rect 16071 2400 16764 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 18046 2428 18052 2440
rect 16899 2400 18052 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18156 2437 18184 2468
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 22296 2468 26065 2496
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 17770 2360 17776 2372
rect 11992 2332 17776 2360
rect 17770 2320 17776 2332
rect 17828 2320 17834 2372
rect 17880 2332 18460 2360
rect 1394 2252 1400 2304
rect 1452 2292 1458 2304
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1452 2264 1777 2292
rect 1452 2252 1458 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9732 2264 9781 2292
rect 9732 2252 9738 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 12986 2292 12992 2304
rect 12947 2264 12992 2292
rect 9769 2255 9827 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16209 2295 16267 2301
rect 16209 2292 16221 2295
rect 16172 2264 16221 2292
rect 16172 2252 16178 2264
rect 16209 2261 16221 2264
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17494 2252 17500 2304
rect 17552 2292 17558 2304
rect 17880 2292 17908 2332
rect 17552 2264 17908 2292
rect 17552 2252 17558 2264
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18432 2292 18460 2332
rect 22296 2292 22324 2468
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26053 2459 26111 2465
rect 30006 2456 30012 2508
rect 30064 2496 30070 2508
rect 35986 2496 35992 2508
rect 30064 2468 31156 2496
rect 30064 2456 30070 2468
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22612 2400 22845 2428
rect 22612 2388 22618 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23256 2400 23489 2428
rect 23256 2388 23262 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 25774 2428 25780 2440
rect 25735 2400 25780 2428
rect 24765 2391 24823 2397
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 27764 2400 27997 2428
rect 27764 2388 27770 2400
rect 27985 2397 27997 2400
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 30374 2428 30380 2440
rect 30335 2400 30380 2428
rect 29917 2391 29975 2397
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 31128 2437 31156 2468
rect 33612 2468 35992 2496
rect 31113 2431 31171 2437
rect 31113 2397 31125 2431
rect 31159 2397 31171 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 31113 2391 31171 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33612 2437 33640 2468
rect 35986 2456 35992 2468
rect 36044 2456 36050 2508
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36630 2428 36636 2440
rect 35952 2400 35997 2428
rect 36591 2400 36636 2428
rect 35952 2388 35958 2400
rect 36630 2388 36636 2400
rect 36688 2388 36694 2440
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 29822 2360 29828 2372
rect 23164 2332 29828 2360
rect 23164 2320 23170 2332
rect 29822 2320 29828 2332
rect 29880 2320 29886 2372
rect 34146 2320 34152 2372
rect 34204 2360 34210 2372
rect 34977 2363 35035 2369
rect 34977 2360 34989 2363
rect 34204 2332 34989 2360
rect 34204 2320 34210 2332
rect 34977 2329 34989 2332
rect 35023 2329 35035 2363
rect 34977 2323 35035 2329
rect 35342 2320 35348 2372
rect 35400 2360 35406 2372
rect 37476 2360 37504 2391
rect 35400 2332 37504 2360
rect 35400 2320 35406 2332
rect 18432 2264 22324 2292
rect 22649 2295 22707 2301
rect 18325 2255 18383 2261
rect 22649 2261 22661 2295
rect 22695 2292 22707 2295
rect 25130 2292 25136 2304
rect 22695 2264 25136 2292
rect 22695 2261 22707 2264
rect 22649 2255 22707 2261
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 30561 2295 30619 2301
rect 30561 2292 30573 2295
rect 30340 2264 30573 2292
rect 30340 2252 30346 2264
rect 30561 2261 30573 2264
rect 30607 2261 30619 2295
rect 30561 2255 30619 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31297 2295 31355 2301
rect 31297 2292 31309 2295
rect 30984 2264 31309 2292
rect 30984 2252 30990 2264
rect 31297 2261 31309 2264
rect 31343 2261 31355 2295
rect 31297 2255 31355 2261
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32272 2264 32505 2292
rect 32272 2252 32278 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 36814 2292 36820 2304
rect 36775 2264 36820 2292
rect 33781 2255 33839 2261
rect 36814 2252 36820 2264
rect 36872 2252 36878 2304
rect 36998 2252 37004 2304
rect 37056 2292 37062 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37056 2264 37657 2292
rect 37056 2252 37062 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 12986 2048 12992 2100
rect 13044 2088 13050 2100
rect 17034 2088 17040 2100
rect 13044 2060 17040 2088
rect 13044 2048 13050 2060
rect 17034 2048 17040 2060
rect 17092 2048 17098 2100
<< via1 >>
rect 19340 37680 19392 37732
rect 20352 37680 20404 37732
rect 17224 37612 17276 37664
rect 27896 37612 27948 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7748 37408 7800 37460
rect 17224 37408 17276 37460
rect 20260 37408 20312 37460
rect 664 37340 716 37392
rect 4620 37340 4672 37392
rect 1584 37315 1636 37324
rect 1584 37281 1593 37315
rect 1593 37281 1627 37315
rect 1627 37281 1636 37315
rect 1584 37272 1636 37281
rect 5172 37315 5224 37324
rect 5172 37281 5181 37315
rect 5181 37281 5215 37315
rect 5215 37281 5224 37315
rect 5172 37272 5224 37281
rect 5816 37272 5868 37324
rect 1952 37204 2004 37256
rect 3792 37204 3844 37256
rect 4068 37204 4120 37256
rect 5448 37247 5500 37256
rect 5448 37213 5457 37247
rect 5457 37213 5491 37247
rect 5491 37213 5500 37247
rect 5448 37204 5500 37213
rect 6644 37204 6696 37256
rect 15200 37340 15252 37392
rect 18420 37383 18472 37392
rect 18420 37349 18429 37383
rect 18429 37349 18463 37383
rect 18463 37349 18472 37383
rect 18420 37340 18472 37349
rect 18788 37383 18840 37392
rect 18788 37349 18797 37383
rect 18797 37349 18831 37383
rect 18831 37349 18840 37383
rect 18788 37340 18840 37349
rect 8484 37204 8536 37256
rect 10232 37272 10284 37324
rect 5080 37136 5132 37188
rect 9128 37136 9180 37188
rect 10048 37204 10100 37256
rect 11612 37272 11664 37324
rect 11796 37315 11848 37324
rect 11796 37281 11805 37315
rect 11805 37281 11839 37315
rect 11839 37281 11848 37315
rect 11796 37272 11848 37281
rect 12256 37272 12308 37324
rect 16120 37272 16172 37324
rect 16488 37272 16540 37324
rect 22928 37315 22980 37324
rect 11704 37247 11756 37256
rect 11704 37213 11713 37247
rect 11713 37213 11747 37247
rect 11747 37213 11756 37247
rect 11704 37204 11756 37213
rect 12440 37204 12492 37256
rect 12900 37204 12952 37256
rect 2780 37068 2832 37120
rect 3884 37068 3936 37120
rect 5816 37068 5868 37120
rect 9680 37111 9732 37120
rect 9680 37077 9689 37111
rect 9689 37077 9723 37111
rect 9723 37077 9732 37111
rect 9680 37068 9732 37077
rect 10232 37068 10284 37120
rect 13636 37136 13688 37188
rect 11980 37068 12032 37120
rect 16672 37204 16724 37256
rect 18328 37204 18380 37256
rect 15016 37136 15068 37188
rect 14832 37068 14884 37120
rect 15108 37068 15160 37120
rect 16488 37068 16540 37120
rect 16580 37068 16632 37120
rect 17776 37136 17828 37188
rect 17224 37068 17276 37120
rect 18420 37136 18472 37188
rect 19340 37204 19392 37256
rect 20812 37204 20864 37256
rect 22928 37281 22937 37315
rect 22937 37281 22971 37315
rect 22971 37281 22980 37315
rect 22928 37272 22980 37281
rect 20996 37204 21048 37256
rect 21272 37204 21324 37256
rect 22560 37204 22612 37256
rect 25504 37272 25556 37324
rect 25780 37272 25832 37324
rect 23204 37204 23256 37256
rect 24768 37204 24820 37256
rect 26240 37204 26292 37256
rect 27068 37204 27120 37256
rect 29644 37272 29696 37324
rect 34060 37272 34112 37324
rect 35164 37315 35216 37324
rect 35164 37281 35173 37315
rect 35173 37281 35207 37315
rect 35207 37281 35216 37315
rect 35164 37272 35216 37281
rect 37464 37315 37516 37324
rect 37464 37281 37473 37315
rect 37473 37281 37507 37315
rect 37507 37281 37516 37315
rect 37464 37272 37516 37281
rect 30012 37247 30064 37256
rect 18972 37068 19024 37120
rect 19984 37068 20036 37120
rect 26424 37136 26476 37188
rect 21180 37111 21232 37120
rect 21180 37077 21189 37111
rect 21189 37077 21223 37111
rect 21223 37077 21232 37111
rect 21180 37068 21232 37077
rect 22008 37111 22060 37120
rect 22008 37077 22017 37111
rect 22017 37077 22051 37111
rect 22051 37077 22060 37111
rect 22008 37068 22060 37077
rect 22100 37068 22152 37120
rect 27712 37136 27764 37188
rect 30012 37213 30021 37247
rect 30021 37213 30055 37247
rect 30055 37213 30064 37247
rect 30012 37204 30064 37213
rect 29000 37136 29052 37188
rect 32220 37204 32272 37256
rect 34520 37204 34572 37256
rect 36176 37247 36228 37256
rect 36176 37213 36185 37247
rect 36185 37213 36219 37247
rect 36219 37213 36228 37247
rect 36176 37204 36228 37213
rect 39672 37204 39724 37256
rect 33140 37136 33192 37188
rect 27620 37068 27672 37120
rect 30288 37068 30340 37120
rect 31024 37111 31076 37120
rect 31024 37077 31033 37111
rect 31033 37077 31067 37111
rect 31067 37077 31076 37111
rect 31024 37068 31076 37077
rect 34152 37111 34204 37120
rect 34152 37077 34161 37111
rect 34161 37077 34195 37111
rect 34195 37077 34204 37111
rect 34152 37068 34204 37077
rect 36084 37068 36136 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1676 36839 1728 36848
rect 1676 36805 1685 36839
rect 1685 36805 1719 36839
rect 1719 36805 1728 36839
rect 1676 36796 1728 36805
rect 3332 36864 3384 36916
rect 5080 36864 5132 36916
rect 8668 36864 8720 36916
rect 9036 36864 9088 36916
rect 9220 36864 9272 36916
rect 11980 36864 12032 36916
rect 13452 36864 13504 36916
rect 13544 36864 13596 36916
rect 13912 36864 13964 36916
rect 22008 36864 22060 36916
rect 25872 36907 25924 36916
rect 2320 36796 2372 36848
rect 3424 36728 3476 36780
rect 7104 36796 7156 36848
rect 7012 36771 7064 36780
rect 2688 36703 2740 36712
rect 2688 36669 2697 36703
rect 2697 36669 2731 36703
rect 2731 36669 2740 36703
rect 2688 36660 2740 36669
rect 7012 36737 7021 36771
rect 7021 36737 7055 36771
rect 7055 36737 7064 36771
rect 7012 36728 7064 36737
rect 11152 36796 11204 36848
rect 15292 36796 15344 36848
rect 20076 36796 20128 36848
rect 20168 36796 20220 36848
rect 9036 36771 9088 36780
rect 5632 36592 5684 36644
rect 3148 36567 3200 36576
rect 3148 36533 3157 36567
rect 3157 36533 3191 36567
rect 3191 36533 3200 36567
rect 3148 36524 3200 36533
rect 5816 36567 5868 36576
rect 5816 36533 5825 36567
rect 5825 36533 5859 36567
rect 5859 36533 5868 36567
rect 5816 36524 5868 36533
rect 8300 36660 8352 36712
rect 9036 36737 9045 36771
rect 9045 36737 9079 36771
rect 9079 36737 9088 36771
rect 9036 36728 9088 36737
rect 10232 36728 10284 36780
rect 10876 36728 10928 36780
rect 8576 36635 8628 36644
rect 7472 36524 7524 36576
rect 7656 36567 7708 36576
rect 7656 36533 7665 36567
rect 7665 36533 7699 36567
rect 7699 36533 7708 36567
rect 7656 36524 7708 36533
rect 8576 36601 8585 36635
rect 8585 36601 8619 36635
rect 8619 36601 8628 36635
rect 8576 36592 8628 36601
rect 8852 36524 8904 36576
rect 9772 36660 9824 36712
rect 13636 36771 13688 36780
rect 11704 36703 11756 36712
rect 11704 36669 11713 36703
rect 11713 36669 11747 36703
rect 11747 36669 11756 36703
rect 11704 36660 11756 36669
rect 13636 36737 13645 36771
rect 13645 36737 13679 36771
rect 13679 36737 13688 36771
rect 13636 36728 13688 36737
rect 13728 36728 13780 36780
rect 17868 36728 17920 36780
rect 20996 36728 21048 36780
rect 22744 36728 22796 36780
rect 13912 36660 13964 36712
rect 15384 36660 15436 36712
rect 16304 36703 16356 36712
rect 16304 36669 16313 36703
rect 16313 36669 16347 36703
rect 16347 36669 16356 36703
rect 16304 36660 16356 36669
rect 10140 36524 10192 36576
rect 10324 36567 10376 36576
rect 10324 36533 10333 36567
rect 10333 36533 10367 36567
rect 10367 36533 10376 36567
rect 10324 36524 10376 36533
rect 11060 36567 11112 36576
rect 11060 36533 11069 36567
rect 11069 36533 11103 36567
rect 11103 36533 11112 36567
rect 11060 36524 11112 36533
rect 12440 36592 12492 36644
rect 12532 36524 12584 36576
rect 12624 36524 12676 36576
rect 16672 36592 16724 36644
rect 16856 36592 16908 36644
rect 17684 36660 17736 36712
rect 18144 36703 18196 36712
rect 18144 36669 18153 36703
rect 18153 36669 18187 36703
rect 18187 36669 18196 36703
rect 18144 36660 18196 36669
rect 18420 36703 18472 36712
rect 18420 36669 18429 36703
rect 18429 36669 18463 36703
rect 18463 36669 18472 36703
rect 18420 36660 18472 36669
rect 19432 36660 19484 36712
rect 20352 36703 20404 36712
rect 20352 36669 20361 36703
rect 20361 36669 20395 36703
rect 20395 36669 20404 36703
rect 20352 36660 20404 36669
rect 20444 36660 20496 36712
rect 21364 36660 21416 36712
rect 25872 36873 25881 36907
rect 25881 36873 25915 36907
rect 25915 36873 25924 36907
rect 25872 36864 25924 36873
rect 24860 36728 24912 36780
rect 17224 36592 17276 36644
rect 19708 36592 19760 36644
rect 20720 36592 20772 36644
rect 14832 36524 14884 36576
rect 17776 36524 17828 36576
rect 18236 36524 18288 36576
rect 23296 36524 23348 36576
rect 23940 36660 23992 36712
rect 25412 36660 25464 36712
rect 31024 36864 31076 36916
rect 32312 36864 32364 36916
rect 32864 36864 32916 36916
rect 26148 36592 26200 36644
rect 26240 36592 26292 36644
rect 27988 36796 28040 36848
rect 29000 36728 29052 36780
rect 27896 36703 27948 36712
rect 27896 36669 27905 36703
rect 27905 36669 27939 36703
rect 27939 36669 27948 36703
rect 27896 36660 27948 36669
rect 27988 36660 28040 36712
rect 29552 36728 29604 36780
rect 30288 36728 30340 36780
rect 33876 36796 33928 36848
rect 32312 36771 32364 36780
rect 32312 36737 32321 36771
rect 32321 36737 32355 36771
rect 32355 36737 32364 36771
rect 32312 36728 32364 36737
rect 33048 36771 33100 36780
rect 33048 36737 33057 36771
rect 33057 36737 33091 36771
rect 33091 36737 33100 36771
rect 33048 36728 33100 36737
rect 36728 36864 36780 36916
rect 37372 36864 37424 36916
rect 35716 36796 35768 36848
rect 23572 36524 23624 36576
rect 24768 36524 24820 36576
rect 26424 36567 26476 36576
rect 26424 36533 26433 36567
rect 26433 36533 26467 36567
rect 26467 36533 26476 36567
rect 26424 36524 26476 36533
rect 27712 36524 27764 36576
rect 27896 36524 27948 36576
rect 32220 36660 32272 36712
rect 34428 36703 34480 36712
rect 34428 36669 34437 36703
rect 34437 36669 34471 36703
rect 34471 36669 34480 36703
rect 34428 36660 34480 36669
rect 34704 36703 34756 36712
rect 34704 36669 34713 36703
rect 34713 36669 34747 36703
rect 34747 36669 34756 36703
rect 34704 36660 34756 36669
rect 31668 36567 31720 36576
rect 31668 36533 31677 36567
rect 31677 36533 31711 36567
rect 31711 36533 31720 36567
rect 31668 36524 31720 36533
rect 33784 36567 33836 36576
rect 33784 36533 33793 36567
rect 33793 36533 33827 36567
rect 33827 36533 33836 36567
rect 33784 36524 33836 36533
rect 35808 36592 35860 36644
rect 36176 36567 36228 36576
rect 36176 36533 36185 36567
rect 36185 36533 36219 36567
rect 36219 36533 36228 36567
rect 36820 36567 36872 36576
rect 36176 36524 36228 36533
rect 36820 36533 36829 36567
rect 36829 36533 36863 36567
rect 36863 36533 36872 36567
rect 36820 36524 36872 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3792 36320 3844 36372
rect 11704 36320 11756 36372
rect 11888 36320 11940 36372
rect 20444 36320 20496 36372
rect 20720 36320 20772 36372
rect 26424 36320 26476 36372
rect 27620 36320 27672 36372
rect 9772 36252 9824 36304
rect 10140 36295 10192 36304
rect 10140 36261 10149 36295
rect 10149 36261 10183 36295
rect 10183 36261 10192 36295
rect 10140 36252 10192 36261
rect 10324 36252 10376 36304
rect 14832 36252 14884 36304
rect 26332 36295 26384 36304
rect 2688 36227 2740 36236
rect 2688 36193 2697 36227
rect 2697 36193 2731 36227
rect 2731 36193 2740 36227
rect 2688 36184 2740 36193
rect 3424 36184 3476 36236
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 4620 36116 4672 36168
rect 7012 36184 7064 36236
rect 7472 36184 7524 36236
rect 8300 36184 8352 36236
rect 6460 36159 6512 36168
rect 6460 36125 6469 36159
rect 6469 36125 6503 36159
rect 6503 36125 6512 36159
rect 6460 36116 6512 36125
rect 7564 36116 7616 36168
rect 7748 36159 7800 36168
rect 7748 36125 7757 36159
rect 7757 36125 7791 36159
rect 7791 36125 7800 36159
rect 7748 36116 7800 36125
rect 10508 36184 10560 36236
rect 9312 36159 9364 36168
rect 9312 36125 9321 36159
rect 9321 36125 9355 36159
rect 9355 36125 9364 36159
rect 9312 36116 9364 36125
rect 10048 36159 10100 36168
rect 10048 36125 10057 36159
rect 10057 36125 10091 36159
rect 10091 36125 10100 36159
rect 10048 36116 10100 36125
rect 10324 36116 10376 36168
rect 10416 36116 10468 36168
rect 12532 36184 12584 36236
rect 13452 36227 13504 36236
rect 13452 36193 13461 36227
rect 13461 36193 13495 36227
rect 13495 36193 13504 36227
rect 13452 36184 13504 36193
rect 16948 36184 17000 36236
rect 17132 36184 17184 36236
rect 19340 36184 19392 36236
rect 26332 36261 26341 36295
rect 26341 36261 26375 36295
rect 26375 36261 26384 36295
rect 26332 36252 26384 36261
rect 20168 36184 20220 36236
rect 23572 36184 23624 36236
rect 27712 36184 27764 36236
rect 14832 36159 14884 36168
rect 2412 36091 2464 36100
rect 2412 36057 2421 36091
rect 2421 36057 2455 36091
rect 2455 36057 2464 36091
rect 2412 36048 2464 36057
rect 2504 36091 2556 36100
rect 2504 36057 2513 36091
rect 2513 36057 2547 36091
rect 2547 36057 2556 36091
rect 2504 36048 2556 36057
rect 3884 35980 3936 36032
rect 5724 35980 5776 36032
rect 9220 36048 9272 36100
rect 10600 36048 10652 36100
rect 10968 36048 11020 36100
rect 11704 36048 11756 36100
rect 12072 36048 12124 36100
rect 12164 36048 12216 36100
rect 14832 36125 14841 36159
rect 14841 36125 14875 36159
rect 14875 36125 14884 36159
rect 14832 36116 14884 36125
rect 18236 36159 18288 36168
rect 15660 36091 15712 36100
rect 15660 36057 15669 36091
rect 15669 36057 15703 36091
rect 15703 36057 15712 36091
rect 16212 36091 16264 36100
rect 15660 36048 15712 36057
rect 16212 36057 16221 36091
rect 16221 36057 16255 36091
rect 16255 36057 16264 36091
rect 16212 36048 16264 36057
rect 16304 36048 16356 36100
rect 17776 36091 17828 36100
rect 7472 35980 7524 36032
rect 7840 35980 7892 36032
rect 10416 35980 10468 36032
rect 15292 35980 15344 36032
rect 17776 36057 17785 36091
rect 17785 36057 17819 36091
rect 17819 36057 17828 36091
rect 17776 36048 17828 36057
rect 18236 36125 18245 36159
rect 18245 36125 18279 36159
rect 18279 36125 18288 36159
rect 18236 36116 18288 36125
rect 19248 36116 19300 36168
rect 33048 36320 33100 36372
rect 33784 36320 33836 36372
rect 37924 36320 37976 36372
rect 28448 36252 28500 36304
rect 29552 36252 29604 36304
rect 33876 36252 33928 36304
rect 37556 36295 37608 36304
rect 32220 36227 32272 36236
rect 32220 36193 32229 36227
rect 32229 36193 32263 36227
rect 32263 36193 32272 36227
rect 32220 36184 32272 36193
rect 34428 36184 34480 36236
rect 37556 36261 37565 36295
rect 37565 36261 37599 36295
rect 37599 36261 37608 36295
rect 37556 36252 37608 36261
rect 35808 36184 35860 36236
rect 19616 36048 19668 36100
rect 17040 35980 17092 36032
rect 20720 36048 20772 36100
rect 20536 35980 20588 36032
rect 20628 35980 20680 36032
rect 21180 36023 21232 36032
rect 21180 35989 21189 36023
rect 21189 35989 21223 36023
rect 21223 35989 21232 36023
rect 21180 35980 21232 35989
rect 21916 36048 21968 36100
rect 23296 36048 23348 36100
rect 37188 36116 37240 36168
rect 38016 36159 38068 36168
rect 38016 36125 38025 36159
rect 38025 36125 38059 36159
rect 38059 36125 38068 36159
rect 38016 36116 38068 36125
rect 23480 36023 23532 36032
rect 23480 35989 23489 36023
rect 23489 35989 23523 36023
rect 23523 35989 23532 36023
rect 23480 35980 23532 35989
rect 24768 36048 24820 36100
rect 24860 36091 24912 36100
rect 24860 36057 24869 36091
rect 24869 36057 24903 36091
rect 24903 36057 24912 36091
rect 24860 36048 24912 36057
rect 24952 35980 25004 36032
rect 25320 36048 25372 36100
rect 26148 36048 26200 36100
rect 27804 36048 27856 36100
rect 28356 36048 28408 36100
rect 27896 35980 27948 36032
rect 28080 35980 28132 36032
rect 29920 36048 29972 36100
rect 30472 36048 30524 36100
rect 31760 36091 31812 36100
rect 31760 36057 31769 36091
rect 31769 36057 31803 36091
rect 31803 36057 31812 36091
rect 31760 36048 31812 36057
rect 31392 35980 31444 36032
rect 34520 36048 34572 36100
rect 34612 36048 34664 36100
rect 33968 36023 34020 36032
rect 33968 35989 33977 36023
rect 33977 35989 34011 36023
rect 34011 35989 34020 36023
rect 33968 35980 34020 35989
rect 36820 36048 36872 36100
rect 35900 35980 35952 36032
rect 35992 35980 36044 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 3332 35819 3384 35828
rect 3332 35785 3341 35819
rect 3341 35785 3375 35819
rect 3375 35785 3384 35819
rect 3332 35776 3384 35785
rect 1676 35751 1728 35760
rect 1676 35717 1685 35751
rect 1685 35717 1719 35751
rect 1719 35717 1728 35751
rect 1676 35708 1728 35717
rect 1768 35751 1820 35760
rect 1768 35717 1777 35751
rect 1777 35717 1811 35751
rect 1811 35717 1820 35751
rect 2688 35751 2740 35760
rect 1768 35708 1820 35717
rect 2688 35717 2697 35751
rect 2697 35717 2731 35751
rect 2731 35717 2740 35751
rect 2688 35708 2740 35717
rect 8576 35708 8628 35760
rect 3240 35683 3292 35692
rect 3240 35649 3249 35683
rect 3249 35649 3283 35683
rect 3283 35649 3292 35683
rect 3240 35640 3292 35649
rect 12992 35776 13044 35828
rect 13452 35776 13504 35828
rect 13544 35776 13596 35828
rect 10324 35708 10376 35760
rect 11612 35708 11664 35760
rect 15292 35708 15344 35760
rect 11244 35640 11296 35692
rect 12072 35640 12124 35692
rect 12440 35683 12492 35692
rect 12440 35649 12449 35683
rect 12449 35649 12483 35683
rect 12483 35649 12492 35683
rect 12440 35640 12492 35649
rect 13820 35640 13872 35692
rect 14832 35640 14884 35692
rect 16212 35776 16264 35828
rect 17040 35751 17092 35760
rect 17040 35717 17049 35751
rect 17049 35717 17083 35751
rect 17083 35717 17092 35751
rect 17040 35708 17092 35717
rect 17776 35776 17828 35828
rect 27528 35776 27580 35828
rect 18512 35708 18564 35760
rect 19432 35708 19484 35760
rect 33968 35776 34020 35828
rect 34336 35776 34388 35828
rect 35716 35776 35768 35828
rect 36728 35776 36780 35828
rect 16764 35640 16816 35692
rect 18144 35683 18196 35692
rect 18144 35649 18153 35683
rect 18153 35649 18187 35683
rect 18187 35649 18196 35683
rect 18144 35640 18196 35649
rect 8852 35572 8904 35624
rect 11152 35572 11204 35624
rect 10968 35504 11020 35556
rect 11244 35504 11296 35556
rect 13912 35572 13964 35624
rect 16672 35572 16724 35624
rect 17776 35572 17828 35624
rect 31392 35708 31444 35760
rect 34704 35708 34756 35760
rect 20260 35640 20312 35692
rect 24676 35640 24728 35692
rect 27620 35640 27672 35692
rect 30288 35683 30340 35692
rect 12808 35504 12860 35556
rect 24768 35572 24820 35624
rect 25136 35615 25188 35624
rect 25136 35581 25145 35615
rect 25145 35581 25179 35615
rect 25179 35581 25188 35615
rect 25136 35572 25188 35581
rect 27436 35615 27488 35624
rect 27436 35581 27445 35615
rect 27445 35581 27479 35615
rect 27479 35581 27488 35615
rect 27436 35572 27488 35581
rect 27712 35572 27764 35624
rect 27988 35615 28040 35624
rect 27988 35581 27997 35615
rect 27997 35581 28031 35615
rect 28031 35581 28040 35615
rect 27988 35572 28040 35581
rect 30288 35649 30297 35683
rect 30297 35649 30331 35683
rect 30331 35649 30340 35683
rect 30288 35640 30340 35649
rect 30472 35640 30524 35692
rect 30840 35640 30892 35692
rect 30932 35640 30984 35692
rect 35808 35640 35860 35692
rect 11704 35436 11756 35488
rect 11888 35479 11940 35488
rect 11888 35445 11897 35479
rect 11897 35445 11931 35479
rect 11931 35445 11940 35479
rect 11888 35436 11940 35445
rect 12072 35436 12124 35488
rect 13820 35436 13872 35488
rect 14832 35479 14884 35488
rect 14832 35445 14841 35479
rect 14841 35445 14875 35479
rect 14875 35445 14884 35479
rect 14832 35436 14884 35445
rect 15476 35479 15528 35488
rect 15476 35445 15485 35479
rect 15485 35445 15519 35479
rect 15519 35445 15528 35479
rect 15476 35436 15528 35445
rect 17224 35436 17276 35488
rect 19984 35436 20036 35488
rect 20996 35436 21048 35488
rect 23848 35436 23900 35488
rect 24860 35436 24912 35488
rect 26516 35436 26568 35488
rect 27528 35436 27580 35488
rect 29368 35436 29420 35488
rect 35440 35572 35492 35624
rect 36820 35640 36872 35692
rect 38292 35572 38344 35624
rect 32864 35504 32916 35556
rect 35992 35504 36044 35556
rect 31484 35436 31536 35488
rect 34704 35436 34756 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 7840 35232 7892 35284
rect 10324 35275 10376 35284
rect 10324 35241 10333 35275
rect 10333 35241 10367 35275
rect 10367 35241 10376 35275
rect 10324 35232 10376 35241
rect 11060 35275 11112 35284
rect 11060 35241 11069 35275
rect 11069 35241 11103 35275
rect 11103 35241 11112 35275
rect 11060 35232 11112 35241
rect 2872 35028 2924 35080
rect 6644 35096 6696 35148
rect 5632 35028 5684 35080
rect 8484 35096 8536 35148
rect 8852 35096 8904 35148
rect 13452 35232 13504 35284
rect 13636 35275 13688 35284
rect 13636 35241 13645 35275
rect 13645 35241 13679 35275
rect 13679 35241 13688 35275
rect 13636 35232 13688 35241
rect 14740 35232 14792 35284
rect 16580 35232 16632 35284
rect 17960 35232 18012 35284
rect 11888 35096 11940 35148
rect 12624 35096 12676 35148
rect 8668 35028 8720 35080
rect 10784 35028 10836 35080
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 10968 35028 11020 35037
rect 11980 35028 12032 35080
rect 6828 34960 6880 35012
rect 2964 34892 3016 34944
rect 9404 34892 9456 34944
rect 9772 34935 9824 34944
rect 9772 34901 9781 34935
rect 9781 34901 9815 34935
rect 9815 34901 9824 34935
rect 9772 34892 9824 34901
rect 10876 34960 10928 35012
rect 21272 35164 21324 35216
rect 23848 35232 23900 35284
rect 24860 35164 24912 35216
rect 12164 34892 12216 34944
rect 15476 35096 15528 35148
rect 20720 35096 20772 35148
rect 24308 35096 24360 35148
rect 24768 35096 24820 35148
rect 31484 35139 31536 35148
rect 13268 35028 13320 35080
rect 13820 35028 13872 35080
rect 14648 35003 14700 35012
rect 13452 34892 13504 34944
rect 14372 34892 14424 34944
rect 14648 34969 14657 35003
rect 14657 34969 14691 35003
rect 14691 34969 14700 35003
rect 14648 34960 14700 34969
rect 14924 34960 14976 35012
rect 15568 35003 15620 35012
rect 15568 34969 15577 35003
rect 15577 34969 15611 35003
rect 15611 34969 15620 35003
rect 15568 34960 15620 34969
rect 16580 35003 16632 35012
rect 16580 34969 16589 35003
rect 16589 34969 16623 35003
rect 16623 34969 16632 35003
rect 16580 34960 16632 34969
rect 16672 34960 16724 35012
rect 20812 35028 20864 35080
rect 31484 35105 31493 35139
rect 31493 35105 31527 35139
rect 31527 35105 31536 35139
rect 31484 35096 31536 35105
rect 31852 35139 31904 35148
rect 31852 35105 31861 35139
rect 31861 35105 31895 35139
rect 31895 35105 31904 35139
rect 31852 35096 31904 35105
rect 32220 35096 32272 35148
rect 32956 35096 33008 35148
rect 34520 35232 34572 35284
rect 36820 35232 36872 35284
rect 38016 35232 38068 35284
rect 39304 35232 39356 35284
rect 34336 35164 34388 35216
rect 26792 35028 26844 35080
rect 19156 34960 19208 35012
rect 20628 34960 20680 35012
rect 22008 34960 22060 35012
rect 24952 34960 25004 35012
rect 26240 34960 26292 35012
rect 26608 34960 26660 35012
rect 36452 35028 36504 35080
rect 37556 35071 37608 35080
rect 37556 35037 37565 35071
rect 37565 35037 37599 35071
rect 37599 35037 37608 35071
rect 37556 35028 37608 35037
rect 37924 35028 37976 35080
rect 29736 35003 29788 35012
rect 29736 34969 29745 35003
rect 29745 34969 29779 35003
rect 29779 34969 29788 35003
rect 29736 34960 29788 34969
rect 30564 35003 30616 35012
rect 30564 34969 30573 35003
rect 30573 34969 30607 35003
rect 30607 34969 30616 35003
rect 30564 34960 30616 34969
rect 31576 35003 31628 35012
rect 31576 34969 31585 35003
rect 31585 34969 31619 35003
rect 31619 34969 31628 35003
rect 32864 35003 32916 35012
rect 31576 34960 31628 34969
rect 32864 34969 32873 35003
rect 32873 34969 32907 35003
rect 32907 34969 32916 35003
rect 32864 34960 32916 34969
rect 36820 34960 36872 35012
rect 22560 34892 22612 34944
rect 26700 34935 26752 34944
rect 26700 34901 26709 34935
rect 26709 34901 26743 34935
rect 26743 34901 26752 34935
rect 26700 34892 26752 34901
rect 27436 34892 27488 34944
rect 31024 34892 31076 34944
rect 34336 34935 34388 34944
rect 34336 34901 34345 34935
rect 34345 34901 34379 34935
rect 34379 34901 34388 34935
rect 34336 34892 34388 34901
rect 36176 34935 36228 34944
rect 36176 34901 36185 34935
rect 36185 34901 36219 34935
rect 36219 34901 36228 34935
rect 36176 34892 36228 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1768 34688 1820 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 8668 34688 8720 34740
rect 9772 34688 9824 34740
rect 8484 34620 8536 34672
rect 10692 34620 10744 34672
rect 11980 34688 12032 34740
rect 13268 34688 13320 34740
rect 13636 34688 13688 34740
rect 14648 34688 14700 34740
rect 14832 34688 14884 34740
rect 19616 34688 19668 34740
rect 21456 34731 21508 34740
rect 11888 34663 11940 34672
rect 11888 34629 11897 34663
rect 11897 34629 11931 34663
rect 11931 34629 11940 34663
rect 11888 34620 11940 34629
rect 8300 34595 8352 34604
rect 8300 34561 8309 34595
rect 8309 34561 8343 34595
rect 8343 34561 8352 34595
rect 8300 34552 8352 34561
rect 11612 34552 11664 34604
rect 9220 34484 9272 34536
rect 9404 34527 9456 34536
rect 9404 34493 9413 34527
rect 9413 34493 9447 34527
rect 9447 34493 9456 34527
rect 9404 34484 9456 34493
rect 11152 34484 11204 34536
rect 13912 34620 13964 34672
rect 14464 34620 14516 34672
rect 15016 34620 15068 34672
rect 17500 34620 17552 34672
rect 9772 34459 9824 34468
rect 9772 34425 9781 34459
rect 9781 34425 9815 34459
rect 9815 34425 9824 34459
rect 9772 34416 9824 34425
rect 10968 34416 11020 34468
rect 13544 34484 13596 34536
rect 14740 34552 14792 34604
rect 17224 34595 17276 34604
rect 17224 34561 17233 34595
rect 17233 34561 17267 34595
rect 17267 34561 17276 34595
rect 17224 34552 17276 34561
rect 21456 34697 21465 34731
rect 21465 34697 21499 34731
rect 21499 34697 21508 34731
rect 21456 34688 21508 34697
rect 21548 34688 21600 34740
rect 19892 34620 19944 34672
rect 21272 34620 21324 34672
rect 27988 34688 28040 34740
rect 24308 34595 24360 34604
rect 12348 34459 12400 34468
rect 12348 34425 12357 34459
rect 12357 34425 12391 34459
rect 12391 34425 12400 34459
rect 12348 34416 12400 34425
rect 13728 34416 13780 34468
rect 15936 34484 15988 34536
rect 24308 34561 24317 34595
rect 24317 34561 24351 34595
rect 24351 34561 24360 34595
rect 24308 34552 24360 34561
rect 30564 34688 30616 34740
rect 36820 34731 36872 34740
rect 31484 34620 31536 34672
rect 33416 34620 33468 34672
rect 30840 34552 30892 34604
rect 34152 34552 34204 34604
rect 16212 34459 16264 34468
rect 16212 34425 16221 34459
rect 16221 34425 16255 34459
rect 16255 34425 16264 34459
rect 16212 34416 16264 34425
rect 18144 34416 18196 34468
rect 19248 34416 19300 34468
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 10140 34348 10192 34400
rect 19616 34416 19668 34468
rect 17132 34348 17184 34400
rect 19340 34348 19392 34400
rect 19432 34348 19484 34400
rect 20720 34484 20772 34536
rect 22008 34527 22060 34536
rect 22008 34493 22017 34527
rect 22017 34493 22051 34527
rect 22051 34493 22060 34527
rect 22008 34484 22060 34493
rect 22284 34527 22336 34536
rect 22284 34493 22293 34527
rect 22293 34493 22327 34527
rect 22327 34493 22336 34527
rect 22284 34484 22336 34493
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 23940 34484 23992 34536
rect 24676 34484 24728 34536
rect 21088 34348 21140 34400
rect 26516 34416 26568 34468
rect 30748 34484 30800 34536
rect 31300 34527 31352 34536
rect 31300 34493 31309 34527
rect 31309 34493 31343 34527
rect 31343 34493 31352 34527
rect 31300 34484 31352 34493
rect 33416 34459 33468 34468
rect 33416 34425 33425 34459
rect 33425 34425 33459 34459
rect 33459 34425 33468 34459
rect 33416 34416 33468 34425
rect 34612 34484 34664 34536
rect 34796 34484 34848 34536
rect 36820 34697 36829 34731
rect 36829 34697 36863 34731
rect 36863 34697 36872 34731
rect 36820 34688 36872 34697
rect 35624 34620 35676 34672
rect 35900 34484 35952 34536
rect 39028 34552 39080 34604
rect 38660 34484 38712 34536
rect 26424 34348 26476 34400
rect 35624 34348 35676 34400
rect 36084 34391 36136 34400
rect 36084 34357 36093 34391
rect 36093 34357 36127 34391
rect 36127 34357 36136 34391
rect 36084 34348 36136 34357
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 8484 34187 8536 34196
rect 8484 34153 8493 34187
rect 8493 34153 8527 34187
rect 8527 34153 8536 34187
rect 8484 34144 8536 34153
rect 10232 34144 10284 34196
rect 11428 34144 11480 34196
rect 13452 34144 13504 34196
rect 13636 34144 13688 34196
rect 12900 34076 12952 34128
rect 12992 34076 13044 34128
rect 15568 34144 15620 34196
rect 15660 34144 15712 34196
rect 16672 34144 16724 34196
rect 19616 34144 19668 34196
rect 20260 34144 20312 34196
rect 21088 34144 21140 34196
rect 21548 34076 21600 34128
rect 9036 33940 9088 33992
rect 10048 34008 10100 34060
rect 26700 34144 26752 34196
rect 34796 34144 34848 34196
rect 10140 33983 10192 33992
rect 10140 33949 10149 33983
rect 10149 33949 10183 33983
rect 10183 33949 10192 33983
rect 10140 33940 10192 33949
rect 10232 33940 10284 33992
rect 10876 33940 10928 33992
rect 11796 33940 11848 33992
rect 13820 33940 13872 33992
rect 9404 33872 9456 33924
rect 11980 33872 12032 33924
rect 12164 33915 12216 33924
rect 12164 33881 12173 33915
rect 12173 33881 12207 33915
rect 12207 33881 12216 33915
rect 12164 33872 12216 33881
rect 12808 33915 12860 33924
rect 3240 33804 3292 33856
rect 8208 33804 8260 33856
rect 9588 33847 9640 33856
rect 9588 33813 9597 33847
rect 9597 33813 9631 33847
rect 9631 33813 9640 33847
rect 9588 33804 9640 33813
rect 9772 33804 9824 33856
rect 10324 33804 10376 33856
rect 12808 33881 12817 33915
rect 12817 33881 12851 33915
rect 12851 33881 12860 33915
rect 12808 33872 12860 33881
rect 13544 33872 13596 33924
rect 15384 33915 15436 33924
rect 15384 33881 15393 33915
rect 15393 33881 15427 33915
rect 15427 33881 15436 33915
rect 15384 33872 15436 33881
rect 16028 33872 16080 33924
rect 16488 33940 16540 33992
rect 19524 33940 19576 33992
rect 19616 33940 19668 33992
rect 25136 34076 25188 34128
rect 26608 34051 26660 34060
rect 26608 34017 26617 34051
rect 26617 34017 26651 34051
rect 26651 34017 26660 34051
rect 26608 34008 26660 34017
rect 22008 33940 22060 33992
rect 17040 33804 17092 33856
rect 19984 33804 20036 33856
rect 21456 33872 21508 33924
rect 23020 33872 23072 33924
rect 24676 33872 24728 33924
rect 25136 33872 25188 33924
rect 27160 33872 27212 33924
rect 27620 33872 27672 33924
rect 24768 33804 24820 33856
rect 24860 33804 24912 33856
rect 29736 34008 29788 34060
rect 34612 34008 34664 34060
rect 35440 34051 35492 34060
rect 35440 34017 35449 34051
rect 35449 34017 35483 34051
rect 35483 34017 35492 34051
rect 35440 34008 35492 34017
rect 34152 33983 34204 33992
rect 34152 33949 34161 33983
rect 34161 33949 34195 33983
rect 34195 33949 34204 33983
rect 34152 33940 34204 33949
rect 31024 33872 31076 33924
rect 31852 33915 31904 33924
rect 28356 33847 28408 33856
rect 28356 33813 28365 33847
rect 28365 33813 28399 33847
rect 28399 33813 28408 33847
rect 28356 33804 28408 33813
rect 31852 33881 31861 33915
rect 31861 33881 31895 33915
rect 31895 33881 31904 33915
rect 31852 33872 31904 33881
rect 32956 33872 33008 33924
rect 34796 33872 34848 33924
rect 32404 33804 32456 33856
rect 33416 33804 33468 33856
rect 36360 33804 36412 33856
rect 36912 33804 36964 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 2504 33600 2556 33652
rect 8576 33643 8628 33652
rect 8576 33609 8585 33643
rect 8585 33609 8619 33643
rect 8619 33609 8628 33643
rect 8576 33600 8628 33609
rect 9588 33600 9640 33652
rect 7472 33532 7524 33584
rect 8300 33464 8352 33516
rect 9404 33464 9456 33516
rect 10324 33532 10376 33584
rect 10416 33532 10468 33584
rect 11980 33532 12032 33584
rect 16304 33600 16356 33652
rect 16580 33600 16632 33652
rect 10140 33507 10192 33516
rect 10140 33473 10149 33507
rect 10149 33473 10183 33507
rect 10183 33473 10192 33507
rect 10140 33464 10192 33473
rect 11060 33464 11112 33516
rect 14464 33575 14516 33584
rect 14464 33541 14473 33575
rect 14473 33541 14507 33575
rect 14507 33541 14516 33575
rect 14464 33532 14516 33541
rect 16488 33532 16540 33584
rect 15016 33464 15068 33516
rect 15568 33507 15620 33516
rect 15568 33473 15577 33507
rect 15577 33473 15611 33507
rect 15611 33473 15620 33507
rect 15568 33464 15620 33473
rect 17040 33507 17092 33516
rect 17040 33473 17049 33507
rect 17049 33473 17083 33507
rect 17083 33473 17092 33507
rect 17040 33464 17092 33473
rect 13820 33439 13872 33448
rect 12532 33328 12584 33380
rect 13820 33405 13829 33439
rect 13829 33405 13863 33439
rect 13863 33405 13872 33439
rect 13820 33396 13872 33405
rect 19984 33600 20036 33652
rect 24676 33600 24728 33652
rect 24768 33600 24820 33652
rect 19800 33532 19852 33584
rect 24860 33532 24912 33584
rect 25136 33575 25188 33584
rect 25136 33541 25145 33575
rect 25145 33541 25179 33575
rect 25179 33541 25188 33575
rect 25136 33532 25188 33541
rect 25596 33532 25648 33584
rect 31576 33600 31628 33652
rect 32404 33643 32456 33652
rect 32404 33609 32413 33643
rect 32413 33609 32447 33643
rect 32447 33609 32456 33643
rect 32404 33600 32456 33609
rect 36452 33600 36504 33652
rect 32864 33532 32916 33584
rect 34704 33532 34756 33584
rect 18144 33439 18196 33448
rect 18144 33405 18153 33439
rect 18153 33405 18187 33439
rect 18187 33405 18196 33439
rect 18144 33396 18196 33405
rect 18880 33396 18932 33448
rect 18972 33396 19024 33448
rect 20168 33396 20220 33448
rect 19708 33328 19760 33380
rect 19892 33371 19944 33380
rect 19892 33337 19901 33371
rect 19901 33337 19935 33371
rect 19935 33337 19944 33371
rect 19892 33328 19944 33337
rect 20260 33328 20312 33380
rect 24400 33396 24452 33448
rect 26516 33396 26568 33448
rect 9864 33260 9916 33312
rect 11980 33260 12032 33312
rect 13820 33260 13872 33312
rect 17592 33260 17644 33312
rect 26424 33260 26476 33312
rect 26608 33303 26660 33312
rect 26608 33269 26617 33303
rect 26617 33269 26651 33303
rect 26651 33269 26660 33303
rect 26608 33260 26660 33269
rect 32956 33507 33008 33516
rect 32956 33473 32965 33507
rect 32965 33473 32999 33507
rect 32999 33473 33008 33507
rect 32956 33464 33008 33473
rect 35532 33507 35584 33516
rect 35532 33473 35541 33507
rect 35541 33473 35575 33507
rect 35575 33473 35584 33507
rect 35532 33464 35584 33473
rect 36360 33507 36412 33516
rect 36360 33473 36369 33507
rect 36369 33473 36403 33507
rect 36403 33473 36412 33507
rect 36360 33464 36412 33473
rect 38108 33507 38160 33516
rect 38108 33473 38117 33507
rect 38117 33473 38151 33507
rect 38151 33473 38160 33507
rect 38108 33464 38160 33473
rect 34520 33396 34572 33448
rect 32312 33328 32364 33380
rect 38844 33328 38896 33380
rect 34520 33260 34572 33312
rect 38016 33260 38068 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2964 32852 3016 32904
rect 5724 32852 5776 32904
rect 12164 33056 12216 33108
rect 12256 33056 12308 33108
rect 15108 33056 15160 33108
rect 15200 33056 15252 33108
rect 10968 32988 11020 33040
rect 7564 32784 7616 32836
rect 9680 32852 9732 32904
rect 10600 32852 10652 32904
rect 14004 32988 14056 33040
rect 14924 32988 14976 33040
rect 20812 33056 20864 33108
rect 21364 33056 21416 33108
rect 22928 33056 22980 33108
rect 11520 32920 11572 32972
rect 15200 32920 15252 32972
rect 17040 32920 17092 32972
rect 17500 32920 17552 32972
rect 19432 32963 19484 32972
rect 19432 32929 19441 32963
rect 19441 32929 19475 32963
rect 19475 32929 19484 32963
rect 19432 32920 19484 32929
rect 24492 32988 24544 33040
rect 13268 32852 13320 32904
rect 15016 32895 15068 32904
rect 15016 32861 15025 32895
rect 15025 32861 15059 32895
rect 15059 32861 15068 32895
rect 15016 32852 15068 32861
rect 18420 32852 18472 32904
rect 22744 32920 22796 32972
rect 26608 32920 26660 32972
rect 30564 32920 30616 32972
rect 34612 33056 34664 33108
rect 34152 32988 34204 33040
rect 37556 33056 37608 33108
rect 33968 32920 34020 32972
rect 23756 32852 23808 32904
rect 24400 32852 24452 32904
rect 34796 32920 34848 32972
rect 37832 32852 37884 32904
rect 38016 32895 38068 32904
rect 38016 32861 38025 32895
rect 38025 32861 38059 32895
rect 38059 32861 38068 32895
rect 38016 32852 38068 32861
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 7288 32759 7340 32768
rect 7288 32725 7297 32759
rect 7297 32725 7331 32759
rect 7331 32725 7340 32759
rect 7288 32716 7340 32725
rect 8392 32759 8444 32768
rect 8392 32725 8401 32759
rect 8401 32725 8435 32759
rect 8435 32725 8444 32759
rect 8392 32716 8444 32725
rect 9772 32784 9824 32836
rect 11980 32827 12032 32836
rect 11980 32793 11989 32827
rect 11989 32793 12023 32827
rect 12023 32793 12032 32827
rect 11980 32784 12032 32793
rect 12164 32784 12216 32836
rect 14464 32827 14516 32836
rect 12256 32716 12308 32768
rect 13636 32759 13688 32768
rect 13636 32725 13645 32759
rect 13645 32725 13679 32759
rect 13679 32725 13688 32759
rect 13636 32716 13688 32725
rect 14464 32793 14473 32827
rect 14473 32793 14507 32827
rect 14507 32793 14516 32827
rect 14464 32784 14516 32793
rect 15844 32784 15896 32836
rect 16120 32827 16172 32836
rect 16120 32793 16129 32827
rect 16129 32793 16163 32827
rect 16163 32793 16172 32827
rect 16120 32784 16172 32793
rect 16764 32784 16816 32836
rect 16856 32784 16908 32836
rect 14740 32716 14792 32768
rect 18972 32716 19024 32768
rect 19432 32784 19484 32836
rect 20720 32784 20772 32836
rect 22652 32784 22704 32836
rect 24308 32784 24360 32836
rect 25504 32784 25556 32836
rect 30656 32784 30708 32836
rect 31668 32784 31720 32836
rect 33140 32784 33192 32836
rect 38568 32784 38620 32836
rect 20444 32716 20496 32768
rect 23940 32716 23992 32768
rect 32312 32716 32364 32768
rect 38200 32759 38252 32768
rect 38200 32725 38209 32759
rect 38209 32725 38243 32759
rect 38243 32725 38252 32759
rect 38200 32716 38252 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 9864 32487 9916 32496
rect 9864 32453 9873 32487
rect 9873 32453 9907 32487
rect 9907 32453 9916 32487
rect 9864 32444 9916 32453
rect 5908 32376 5960 32428
rect 9220 32419 9272 32428
rect 9220 32385 9229 32419
rect 9229 32385 9263 32419
rect 9263 32385 9272 32419
rect 9220 32376 9272 32385
rect 9772 32351 9824 32360
rect 9772 32317 9781 32351
rect 9781 32317 9815 32351
rect 9815 32317 9824 32351
rect 9772 32308 9824 32317
rect 12532 32512 12584 32564
rect 13360 32444 13412 32496
rect 16120 32512 16172 32564
rect 17868 32512 17920 32564
rect 13544 32376 13596 32428
rect 11796 32351 11848 32360
rect 11796 32317 11805 32351
rect 11805 32317 11839 32351
rect 11839 32317 11848 32351
rect 11796 32308 11848 32317
rect 14004 32419 14056 32428
rect 14004 32385 14013 32419
rect 14013 32385 14047 32419
rect 14047 32385 14056 32419
rect 14004 32376 14056 32385
rect 14924 32419 14976 32428
rect 14924 32385 14933 32419
rect 14933 32385 14967 32419
rect 14967 32385 14976 32419
rect 14924 32376 14976 32385
rect 15476 32444 15528 32496
rect 16028 32444 16080 32496
rect 17408 32444 17460 32496
rect 19340 32512 19392 32564
rect 19616 32512 19668 32564
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 8668 32172 8720 32224
rect 12348 32283 12400 32292
rect 12348 32249 12357 32283
rect 12357 32249 12391 32283
rect 12391 32249 12400 32283
rect 12348 32240 12400 32249
rect 15844 32308 15896 32360
rect 17960 32308 18012 32360
rect 18236 32308 18288 32360
rect 18696 32308 18748 32360
rect 12256 32172 12308 32224
rect 12716 32172 12768 32224
rect 22652 32512 22704 32564
rect 24124 32512 24176 32564
rect 20260 32444 20312 32496
rect 23940 32444 23992 32496
rect 24308 32444 24360 32496
rect 29368 32512 29420 32564
rect 33416 32512 33468 32564
rect 24492 32444 24544 32496
rect 34244 32444 34296 32496
rect 36728 32512 36780 32564
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 22284 32376 22336 32428
rect 22744 32419 22796 32428
rect 22744 32385 22753 32419
rect 22753 32385 22787 32419
rect 22787 32385 22796 32419
rect 22744 32376 22796 32385
rect 23756 32419 23808 32428
rect 23756 32385 23765 32419
rect 23765 32385 23799 32419
rect 23799 32385 23808 32419
rect 23756 32376 23808 32385
rect 20444 32308 20496 32360
rect 31760 32376 31812 32428
rect 34796 32376 34848 32428
rect 36268 32376 36320 32428
rect 36820 32376 36872 32428
rect 25780 32351 25832 32360
rect 25780 32317 25789 32351
rect 25789 32317 25823 32351
rect 25823 32317 25832 32351
rect 25780 32308 25832 32317
rect 35900 32308 35952 32360
rect 21272 32240 21324 32292
rect 23664 32240 23716 32292
rect 36452 32308 36504 32360
rect 19984 32172 20036 32224
rect 21916 32172 21968 32224
rect 23756 32172 23808 32224
rect 24400 32172 24452 32224
rect 24584 32172 24636 32224
rect 25320 32172 25372 32224
rect 27344 32215 27396 32224
rect 27344 32181 27353 32215
rect 27353 32181 27387 32215
rect 27387 32181 27396 32215
rect 27344 32172 27396 32181
rect 37832 32215 37884 32224
rect 37832 32181 37841 32215
rect 37841 32181 37875 32215
rect 37875 32181 37884 32215
rect 37832 32172 37884 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 9772 31968 9824 32020
rect 11336 31968 11388 32020
rect 8944 31900 8996 31952
rect 6828 31764 6880 31816
rect 6920 31764 6972 31816
rect 9128 31764 9180 31816
rect 12256 31900 12308 31952
rect 14924 31900 14976 31952
rect 15384 31968 15436 32020
rect 15752 31968 15804 32020
rect 15844 31968 15896 32020
rect 16396 31968 16448 32020
rect 16948 31968 17000 32020
rect 17592 31968 17644 32020
rect 19432 31968 19484 32020
rect 23664 31968 23716 32020
rect 11704 31832 11756 31884
rect 12072 31875 12124 31884
rect 12072 31841 12081 31875
rect 12081 31841 12115 31875
rect 12115 31841 12124 31875
rect 12072 31832 12124 31841
rect 12808 31832 12860 31884
rect 11060 31764 11112 31816
rect 13176 31764 13228 31816
rect 13268 31696 13320 31748
rect 14372 31807 14424 31816
rect 14372 31773 14381 31807
rect 14381 31773 14415 31807
rect 14415 31773 14424 31807
rect 14372 31764 14424 31773
rect 16396 31807 16448 31816
rect 16396 31773 16405 31807
rect 16405 31773 16439 31807
rect 16439 31773 16448 31807
rect 16396 31764 16448 31773
rect 23756 31900 23808 31952
rect 24124 31900 24176 31952
rect 24308 31900 24360 31952
rect 24584 31968 24636 32020
rect 24584 31875 24636 31884
rect 16856 31764 16908 31816
rect 15844 31739 15896 31748
rect 15844 31705 15853 31739
rect 15853 31705 15887 31739
rect 15887 31705 15896 31739
rect 15844 31696 15896 31705
rect 16580 31696 16632 31748
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 10048 31671 10100 31680
rect 10048 31637 10057 31671
rect 10057 31637 10091 31671
rect 10091 31637 10100 31671
rect 10048 31628 10100 31637
rect 10876 31628 10928 31680
rect 10968 31628 11020 31680
rect 13912 31628 13964 31680
rect 15016 31628 15068 31680
rect 19064 31696 19116 31748
rect 18236 31628 18288 31680
rect 19616 31696 19668 31748
rect 20168 31696 20220 31748
rect 20996 31628 21048 31680
rect 22100 31739 22152 31748
rect 22100 31705 22109 31739
rect 22109 31705 22143 31739
rect 22143 31705 22152 31739
rect 22100 31696 22152 31705
rect 22560 31696 22612 31748
rect 24584 31841 24593 31875
rect 24593 31841 24627 31875
rect 24627 31841 24636 31875
rect 24584 31832 24636 31841
rect 24952 31832 25004 31884
rect 27344 31968 27396 32020
rect 37004 31968 37056 32020
rect 36912 31832 36964 31884
rect 36176 31764 36228 31816
rect 38292 31807 38344 31816
rect 25320 31696 25372 31748
rect 26792 31696 26844 31748
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 39396 31764 39448 31816
rect 25504 31628 25556 31680
rect 31300 31628 31352 31680
rect 36912 31628 36964 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 9220 31424 9272 31476
rect 10416 31467 10468 31476
rect 10416 31433 10425 31467
rect 10425 31433 10459 31467
rect 10459 31433 10468 31467
rect 10416 31424 10468 31433
rect 14832 31424 14884 31476
rect 15476 31424 15528 31476
rect 15292 31399 15344 31408
rect 15292 31365 15301 31399
rect 15301 31365 15335 31399
rect 15335 31365 15344 31399
rect 15292 31356 15344 31365
rect 19432 31424 19484 31476
rect 3884 31288 3936 31340
rect 9036 31288 9088 31340
rect 8484 31127 8536 31136
rect 8484 31093 8493 31127
rect 8493 31093 8527 31127
rect 8527 31093 8536 31127
rect 8484 31084 8536 31093
rect 9312 31288 9364 31340
rect 10968 31331 11020 31340
rect 10968 31297 10977 31331
rect 10977 31297 11011 31331
rect 11011 31297 11020 31331
rect 10968 31288 11020 31297
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 13176 31288 13228 31340
rect 13912 31288 13964 31340
rect 18972 31356 19024 31408
rect 20536 31399 20588 31408
rect 20536 31365 20545 31399
rect 20545 31365 20579 31399
rect 20579 31365 20588 31399
rect 20536 31356 20588 31365
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 14004 31220 14056 31272
rect 15200 31220 15252 31272
rect 18512 31263 18564 31272
rect 18512 31229 18521 31263
rect 18521 31229 18555 31263
rect 18555 31229 18564 31263
rect 25228 31424 25280 31476
rect 36820 31467 36872 31476
rect 36820 31433 36829 31467
rect 36829 31433 36863 31467
rect 36863 31433 36872 31467
rect 36820 31424 36872 31433
rect 21088 31288 21140 31340
rect 22468 31288 22520 31340
rect 24584 31288 24636 31340
rect 27436 31356 27488 31408
rect 30564 31356 30616 31408
rect 28632 31288 28684 31340
rect 33784 31288 33836 31340
rect 36728 31331 36780 31340
rect 36728 31297 36737 31331
rect 36737 31297 36771 31331
rect 36771 31297 36780 31331
rect 36728 31288 36780 31297
rect 18512 31220 18564 31229
rect 20996 31220 21048 31272
rect 23480 31263 23532 31272
rect 23480 31229 23489 31263
rect 23489 31229 23523 31263
rect 23523 31229 23532 31263
rect 23480 31220 23532 31229
rect 25412 31263 25464 31272
rect 25412 31229 25421 31263
rect 25421 31229 25455 31263
rect 25455 31229 25464 31263
rect 25412 31220 25464 31229
rect 25504 31220 25556 31272
rect 29828 31263 29880 31272
rect 29828 31229 29837 31263
rect 29837 31229 29871 31263
rect 29871 31229 29880 31263
rect 29828 31220 29880 31229
rect 32128 31220 32180 31272
rect 32404 31263 32456 31272
rect 32404 31229 32413 31263
rect 32413 31229 32447 31263
rect 32447 31229 32456 31263
rect 32404 31220 32456 31229
rect 32772 31220 32824 31272
rect 34336 31220 34388 31272
rect 37464 31220 37516 31272
rect 11060 31195 11112 31204
rect 11060 31161 11069 31195
rect 11069 31161 11103 31195
rect 11103 31161 11112 31195
rect 11060 31152 11112 31161
rect 17316 31152 17368 31204
rect 17500 31152 17552 31204
rect 13544 31084 13596 31136
rect 17868 31084 17920 31136
rect 21640 31152 21692 31204
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 22652 31084 22704 31136
rect 25228 31084 25280 31136
rect 30472 31084 30524 31136
rect 31208 31084 31260 31136
rect 31576 31127 31628 31136
rect 31576 31093 31585 31127
rect 31585 31093 31619 31127
rect 31619 31093 31628 31127
rect 31576 31084 31628 31093
rect 34244 31084 34296 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 10416 30880 10468 30932
rect 16856 30923 16908 30932
rect 11152 30812 11204 30864
rect 16856 30889 16865 30923
rect 16865 30889 16899 30923
rect 16899 30889 16908 30923
rect 16856 30880 16908 30889
rect 18880 30923 18932 30932
rect 15568 30812 15620 30864
rect 18880 30889 18889 30923
rect 18889 30889 18923 30923
rect 18923 30889 18932 30923
rect 18880 30880 18932 30889
rect 19156 30880 19208 30932
rect 8300 30744 8352 30796
rect 8484 30744 8536 30796
rect 10140 30744 10192 30796
rect 11244 30787 11296 30796
rect 11244 30753 11253 30787
rect 11253 30753 11287 30787
rect 11287 30753 11296 30787
rect 11244 30744 11296 30753
rect 11428 30744 11480 30796
rect 15752 30744 15804 30796
rect 18144 30744 18196 30796
rect 18420 30744 18472 30796
rect 18696 30744 18748 30796
rect 19984 30744 20036 30796
rect 20996 30787 21048 30796
rect 20996 30753 21005 30787
rect 21005 30753 21039 30787
rect 21039 30753 21048 30787
rect 20996 30744 21048 30753
rect 26332 30812 26384 30864
rect 25412 30744 25464 30796
rect 34612 30880 34664 30932
rect 37832 30923 37884 30932
rect 37832 30889 37841 30923
rect 37841 30889 37875 30923
rect 37875 30889 37884 30923
rect 37832 30880 37884 30889
rect 27252 30744 27304 30796
rect 30472 30744 30524 30796
rect 34244 30744 34296 30796
rect 38384 30812 38436 30864
rect 37464 30787 37516 30796
rect 37464 30753 37473 30787
rect 37473 30753 37507 30787
rect 37507 30753 37516 30787
rect 37464 30744 37516 30753
rect 3148 30676 3200 30728
rect 8392 30608 8444 30660
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 8208 30540 8260 30592
rect 27436 30719 27488 30728
rect 10048 30608 10100 30660
rect 10416 30608 10468 30660
rect 10876 30651 10928 30660
rect 10876 30617 10885 30651
rect 10885 30617 10919 30651
rect 10919 30617 10928 30651
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 29920 30676 29972 30728
rect 32404 30676 32456 30728
rect 34704 30676 34756 30728
rect 37556 30676 37608 30728
rect 10876 30608 10928 30617
rect 12716 30651 12768 30660
rect 12716 30617 12725 30651
rect 12725 30617 12759 30651
rect 12759 30617 12768 30651
rect 13268 30651 13320 30660
rect 12716 30608 12768 30617
rect 13268 30617 13277 30651
rect 13277 30617 13311 30651
rect 13311 30617 13320 30651
rect 13268 30608 13320 30617
rect 13360 30608 13412 30660
rect 13912 30608 13964 30660
rect 15200 30608 15252 30660
rect 15292 30608 15344 30660
rect 11888 30540 11940 30592
rect 13084 30540 13136 30592
rect 17500 30608 17552 30660
rect 17960 30608 18012 30660
rect 21272 30651 21324 30660
rect 21272 30617 21281 30651
rect 21281 30617 21315 30651
rect 21315 30617 21324 30651
rect 21272 30608 21324 30617
rect 16672 30540 16724 30592
rect 17316 30540 17368 30592
rect 22928 30608 22980 30660
rect 24308 30608 24360 30660
rect 27804 30608 27856 30660
rect 32036 30608 32088 30660
rect 33416 30651 33468 30660
rect 33416 30617 33425 30651
rect 33425 30617 33459 30651
rect 33459 30617 33468 30651
rect 33416 30608 33468 30617
rect 39212 30608 39264 30660
rect 29828 30540 29880 30592
rect 30196 30540 30248 30592
rect 36636 30583 36688 30592
rect 36636 30549 36645 30583
rect 36645 30549 36679 30583
rect 36679 30549 36688 30583
rect 36636 30540 36688 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 10600 30336 10652 30388
rect 16856 30336 16908 30388
rect 17040 30336 17092 30388
rect 21272 30336 21324 30388
rect 29552 30336 29604 30388
rect 38200 30379 38252 30388
rect 14188 30311 14240 30320
rect 14188 30277 14197 30311
rect 14197 30277 14231 30311
rect 14231 30277 14240 30311
rect 14188 30268 14240 30277
rect 14740 30311 14792 30320
rect 14740 30277 14749 30311
rect 14749 30277 14783 30311
rect 14783 30277 14792 30311
rect 14740 30268 14792 30277
rect 15292 30311 15344 30320
rect 15292 30277 15301 30311
rect 15301 30277 15335 30311
rect 15335 30277 15344 30311
rect 15292 30268 15344 30277
rect 15384 30311 15436 30320
rect 15384 30277 15393 30311
rect 15393 30277 15427 30311
rect 15427 30277 15436 30311
rect 15384 30268 15436 30277
rect 16672 30268 16724 30320
rect 10232 30200 10284 30252
rect 9956 30132 10008 30184
rect 11336 30200 11388 30252
rect 11980 30200 12032 30252
rect 12808 30200 12860 30252
rect 13176 30243 13228 30252
rect 13176 30209 13185 30243
rect 13185 30209 13219 30243
rect 13219 30209 13228 30243
rect 13176 30200 13228 30209
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 13268 30132 13320 30184
rect 14464 30132 14516 30184
rect 14924 30132 14976 30184
rect 15568 30175 15620 30184
rect 11244 30064 11296 30116
rect 13176 30064 13228 30116
rect 9496 29996 9548 30048
rect 11980 29996 12032 30048
rect 15016 30064 15068 30116
rect 15568 30141 15577 30175
rect 15577 30141 15611 30175
rect 15611 30141 15620 30175
rect 15568 30132 15620 30141
rect 19800 30268 19852 30320
rect 21180 30268 21232 30320
rect 23388 30268 23440 30320
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 18604 30132 18656 30184
rect 18236 30064 18288 30116
rect 13544 29996 13596 30048
rect 23480 30200 23532 30252
rect 24216 30243 24268 30252
rect 24216 30209 24225 30243
rect 24225 30209 24259 30243
rect 24259 30209 24268 30243
rect 24216 30200 24268 30209
rect 27528 30268 27580 30320
rect 29276 30268 29328 30320
rect 30196 30311 30248 30320
rect 30196 30277 30205 30311
rect 30205 30277 30239 30311
rect 30239 30277 30248 30311
rect 30196 30268 30248 30277
rect 31484 30268 31536 30320
rect 28540 30200 28592 30252
rect 31300 30200 31352 30252
rect 35072 30268 35124 30320
rect 38200 30345 38209 30379
rect 38209 30345 38243 30379
rect 38243 30345 38252 30379
rect 38200 30336 38252 30345
rect 34704 30243 34756 30252
rect 34704 30209 34713 30243
rect 34713 30209 34747 30243
rect 34747 30209 34756 30243
rect 34704 30200 34756 30209
rect 36084 30200 36136 30252
rect 37004 30200 37056 30252
rect 20168 30132 20220 30184
rect 20628 29996 20680 30048
rect 24216 30064 24268 30116
rect 23940 29996 23992 30048
rect 24676 29996 24728 30048
rect 24860 29996 24912 30048
rect 27528 30132 27580 30184
rect 29920 30175 29972 30184
rect 29920 30141 29929 30175
rect 29929 30141 29963 30175
rect 29963 30141 29972 30175
rect 29920 30132 29972 30141
rect 34612 30132 34664 30184
rect 35072 30132 35124 30184
rect 36360 30132 36412 30184
rect 28080 29996 28132 30048
rect 28908 30039 28960 30048
rect 28908 30005 28917 30039
rect 28917 30005 28951 30039
rect 28951 30005 28960 30039
rect 28908 29996 28960 30005
rect 31392 29996 31444 30048
rect 31668 30039 31720 30048
rect 31668 30005 31677 30039
rect 31677 30005 31711 30039
rect 31711 30005 31720 30039
rect 31668 29996 31720 30005
rect 32128 29996 32180 30048
rect 33048 29996 33100 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 8208 29835 8260 29844
rect 8208 29801 8217 29835
rect 8217 29801 8251 29835
rect 8251 29801 8260 29835
rect 8208 29792 8260 29801
rect 11796 29792 11848 29844
rect 13176 29792 13228 29844
rect 14740 29792 14792 29844
rect 15844 29792 15896 29844
rect 16856 29792 16908 29844
rect 19064 29792 19116 29844
rect 9312 29724 9364 29776
rect 13268 29724 13320 29776
rect 18972 29724 19024 29776
rect 19800 29792 19852 29844
rect 26884 29792 26936 29844
rect 20904 29724 20956 29776
rect 23572 29724 23624 29776
rect 9956 29699 10008 29708
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 11520 29699 11572 29708
rect 11520 29665 11529 29699
rect 11529 29665 11563 29699
rect 11563 29665 11572 29699
rect 11520 29656 11572 29665
rect 13084 29699 13136 29708
rect 13084 29665 13093 29699
rect 13093 29665 13127 29699
rect 13127 29665 13136 29699
rect 13084 29656 13136 29665
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 7288 29588 7340 29640
rect 7564 29631 7616 29640
rect 7564 29597 7573 29631
rect 7573 29597 7607 29631
rect 7607 29597 7616 29631
rect 7564 29588 7616 29597
rect 7748 29631 7800 29640
rect 7748 29597 7757 29631
rect 7757 29597 7791 29631
rect 7791 29597 7800 29631
rect 7748 29588 7800 29597
rect 9496 29631 9548 29640
rect 9496 29597 9505 29631
rect 9505 29597 9539 29631
rect 9539 29597 9548 29631
rect 9496 29588 9548 29597
rect 9680 29588 9732 29640
rect 22100 29656 22152 29708
rect 24860 29656 24912 29708
rect 25596 29656 25648 29708
rect 18144 29588 18196 29640
rect 11152 29563 11204 29572
rect 11152 29529 11161 29563
rect 11161 29529 11195 29563
rect 11195 29529 11204 29563
rect 11152 29520 11204 29529
rect 11244 29563 11296 29572
rect 11244 29529 11253 29563
rect 11253 29529 11287 29563
rect 11287 29529 11296 29563
rect 11244 29520 11296 29529
rect 13176 29563 13228 29572
rect 13176 29529 13185 29563
rect 13185 29529 13219 29563
rect 13219 29529 13228 29563
rect 15476 29563 15528 29572
rect 13176 29520 13228 29529
rect 15476 29529 15485 29563
rect 15485 29529 15519 29563
rect 15519 29529 15528 29563
rect 15476 29520 15528 29529
rect 15568 29563 15620 29572
rect 15568 29529 15577 29563
rect 15577 29529 15611 29563
rect 15611 29529 15620 29563
rect 15568 29520 15620 29529
rect 20168 29520 20220 29572
rect 5908 29452 5960 29504
rect 9404 29452 9456 29504
rect 12900 29452 12952 29504
rect 19340 29452 19392 29504
rect 21272 29452 21324 29504
rect 24492 29588 24544 29640
rect 22928 29520 22980 29572
rect 26608 29520 26660 29572
rect 35348 29792 35400 29844
rect 33048 29724 33100 29776
rect 29920 29656 29972 29708
rect 32404 29656 32456 29708
rect 34704 29656 34756 29708
rect 29552 29520 29604 29572
rect 36728 29588 36780 29640
rect 37832 29588 37884 29640
rect 31668 29563 31720 29572
rect 31668 29529 31677 29563
rect 31677 29529 31711 29563
rect 31711 29529 31720 29563
rect 31668 29520 31720 29529
rect 32220 29520 32272 29572
rect 23572 29452 23624 29504
rect 25136 29452 25188 29504
rect 27436 29452 27488 29504
rect 28080 29452 28132 29504
rect 29644 29452 29696 29504
rect 33140 29495 33192 29504
rect 33140 29461 33149 29495
rect 33149 29461 33183 29495
rect 33183 29461 33192 29495
rect 33140 29452 33192 29461
rect 34152 29452 34204 29504
rect 37924 29520 37976 29572
rect 37648 29452 37700 29504
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 6644 29180 6696 29232
rect 1860 29112 1912 29164
rect 7656 29112 7708 29164
rect 10048 29112 10100 29164
rect 13176 29248 13228 29300
rect 10968 29155 11020 29164
rect 10968 29121 10977 29155
rect 10977 29121 11011 29155
rect 11011 29121 11020 29155
rect 10968 29112 11020 29121
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 13544 29155 13596 29164
rect 12900 29112 12952 29121
rect 11428 29044 11480 29096
rect 12164 29087 12216 29096
rect 1768 29019 1820 29028
rect 1768 28985 1777 29019
rect 1777 28985 1811 29019
rect 1811 28985 1820 29019
rect 1768 28976 1820 28985
rect 7564 28976 7616 29028
rect 9772 28976 9824 29028
rect 12164 29053 12173 29087
rect 12173 29053 12207 29087
rect 12207 29053 12216 29087
rect 12164 29044 12216 29053
rect 11244 28908 11296 28960
rect 12072 28908 12124 28960
rect 12992 28951 13044 28960
rect 12992 28917 13001 28951
rect 13001 28917 13035 28951
rect 13035 28917 13044 28951
rect 12992 28908 13044 28917
rect 13544 29121 13553 29155
rect 13553 29121 13587 29155
rect 13587 29121 13596 29155
rect 13544 29112 13596 29121
rect 13728 29180 13780 29232
rect 15660 29223 15712 29232
rect 15660 29189 15662 29223
rect 15662 29189 15696 29223
rect 15696 29189 15712 29223
rect 15660 29180 15712 29189
rect 21272 29248 21324 29300
rect 17960 29180 18012 29232
rect 20536 29223 20588 29232
rect 20536 29189 20545 29223
rect 20545 29189 20579 29223
rect 20579 29189 20588 29223
rect 20536 29180 20588 29189
rect 22100 29180 22152 29232
rect 23296 29223 23348 29232
rect 23296 29189 23305 29223
rect 23305 29189 23339 29223
rect 23339 29189 23348 29223
rect 23296 29180 23348 29189
rect 23848 29180 23900 29232
rect 26792 29248 26844 29300
rect 28080 29248 28132 29300
rect 33600 29248 33652 29300
rect 33232 29180 33284 29232
rect 13820 29044 13872 29096
rect 14556 29044 14608 29096
rect 14832 29044 14884 29096
rect 15936 29044 15988 29096
rect 16304 29044 16356 29096
rect 18144 29044 18196 29096
rect 15292 28976 15344 29028
rect 20720 29044 20772 29096
rect 21548 29112 21600 29164
rect 22928 29112 22980 29164
rect 24584 29112 24636 29164
rect 31576 29112 31628 29164
rect 32404 29112 32456 29164
rect 39120 29112 39172 29164
rect 22560 29044 22612 29096
rect 23020 29087 23072 29096
rect 23020 29053 23029 29087
rect 23029 29053 23063 29087
rect 23063 29053 23072 29087
rect 23020 29044 23072 29053
rect 19984 29019 20036 29028
rect 16948 28951 17000 28960
rect 16948 28917 16957 28951
rect 16957 28917 16991 28951
rect 16991 28917 17000 28951
rect 16948 28908 17000 28917
rect 17776 28908 17828 28960
rect 18972 28908 19024 28960
rect 19248 28908 19300 28960
rect 19984 28985 19993 29019
rect 19993 28985 20027 29019
rect 20027 28985 20036 29019
rect 19984 28976 20036 28985
rect 20996 28976 21048 29028
rect 21088 28976 21140 29028
rect 24860 29044 24912 29096
rect 26884 29044 26936 29096
rect 32312 29044 32364 29096
rect 24952 28976 25004 29028
rect 25596 28976 25648 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 20076 28908 20128 28960
rect 26884 28908 26936 28960
rect 32588 28908 32640 28960
rect 36636 28908 36688 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1584 28704 1636 28756
rect 10508 28747 10560 28756
rect 10508 28713 10517 28747
rect 10517 28713 10551 28747
rect 10551 28713 10560 28747
rect 10508 28704 10560 28713
rect 11796 28704 11848 28756
rect 13728 28704 13780 28756
rect 14188 28704 14240 28756
rect 15384 28704 15436 28756
rect 5448 28636 5500 28688
rect 8208 28568 8260 28620
rect 7932 28543 7984 28552
rect 7932 28509 7941 28543
rect 7941 28509 7975 28543
rect 7975 28509 7984 28543
rect 7932 28500 7984 28509
rect 11336 28636 11388 28688
rect 17868 28704 17920 28756
rect 20076 28704 20128 28756
rect 20352 28704 20404 28756
rect 20812 28704 20864 28756
rect 20996 28704 21048 28756
rect 12992 28568 13044 28620
rect 11612 28500 11664 28552
rect 12256 28500 12308 28552
rect 12808 28543 12860 28552
rect 12808 28509 12817 28543
rect 12817 28509 12851 28543
rect 12851 28509 12860 28543
rect 12808 28500 12860 28509
rect 13728 28500 13780 28552
rect 15936 28568 15988 28620
rect 16948 28568 17000 28620
rect 14924 28543 14976 28552
rect 14924 28509 14933 28543
rect 14933 28509 14967 28543
rect 14967 28509 14976 28543
rect 16028 28543 16080 28552
rect 14924 28500 14976 28509
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 17500 28500 17552 28552
rect 8208 28432 8260 28484
rect 15936 28432 15988 28484
rect 20352 28568 20404 28620
rect 20720 28611 20772 28620
rect 20720 28577 20729 28611
rect 20729 28577 20763 28611
rect 20763 28577 20772 28611
rect 20720 28568 20772 28577
rect 21732 28568 21784 28620
rect 26884 28704 26936 28756
rect 17776 28500 17828 28552
rect 20444 28500 20496 28552
rect 17684 28432 17736 28484
rect 19984 28432 20036 28484
rect 20996 28475 21048 28484
rect 20996 28441 21005 28475
rect 21005 28441 21039 28475
rect 21039 28441 21048 28475
rect 20996 28432 21048 28441
rect 8392 28407 8444 28416
rect 8392 28373 8401 28407
rect 8401 28373 8435 28407
rect 8435 28373 8444 28407
rect 8392 28364 8444 28373
rect 11152 28364 11204 28416
rect 12348 28364 12400 28416
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 15200 28364 15252 28416
rect 22560 28432 22612 28484
rect 23020 28500 23072 28552
rect 24860 28568 24912 28620
rect 26148 28568 26200 28620
rect 26700 28568 26752 28620
rect 37556 28704 37608 28756
rect 27620 28500 27672 28552
rect 31116 28543 31168 28552
rect 31116 28509 31125 28543
rect 31125 28509 31159 28543
rect 31159 28509 31168 28543
rect 31116 28500 31168 28509
rect 34796 28500 34848 28552
rect 37648 28543 37700 28552
rect 37648 28509 37657 28543
rect 37657 28509 37691 28543
rect 37691 28509 37700 28543
rect 37648 28500 37700 28509
rect 25320 28432 25372 28484
rect 28080 28475 28132 28484
rect 28080 28441 28089 28475
rect 28089 28441 28123 28475
rect 28123 28441 28132 28475
rect 28080 28432 28132 28441
rect 32036 28432 32088 28484
rect 21732 28364 21784 28416
rect 31668 28364 31720 28416
rect 32864 28407 32916 28416
rect 32864 28373 32873 28407
rect 32873 28373 32907 28407
rect 32907 28373 32916 28407
rect 34060 28432 34112 28484
rect 38660 28432 38712 28484
rect 32864 28364 32916 28373
rect 38016 28364 38068 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 7932 28160 7984 28212
rect 8208 28203 8260 28212
rect 8208 28169 8217 28203
rect 8217 28169 8251 28203
rect 8251 28169 8260 28203
rect 8208 28160 8260 28169
rect 7748 28092 7800 28144
rect 23940 28160 23992 28212
rect 24032 28160 24084 28212
rect 36452 28160 36504 28212
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 7104 28024 7156 28076
rect 10048 28092 10100 28144
rect 9772 28024 9824 28076
rect 10784 28024 10836 28076
rect 10508 27956 10560 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 13912 28092 13964 28144
rect 14188 28135 14240 28144
rect 14188 28101 14197 28135
rect 14197 28101 14231 28135
rect 14231 28101 14240 28135
rect 14188 28092 14240 28101
rect 15384 28135 15436 28144
rect 15384 28101 15393 28135
rect 15393 28101 15427 28135
rect 15427 28101 15436 28135
rect 15384 28092 15436 28101
rect 19524 28092 19576 28144
rect 20444 28092 20496 28144
rect 26056 28092 26108 28144
rect 29736 28092 29788 28144
rect 33416 28092 33468 28144
rect 12440 27956 12492 27965
rect 10324 27931 10376 27940
rect 10324 27897 10333 27931
rect 10333 27897 10367 27931
rect 10367 27897 10376 27931
rect 10324 27888 10376 27897
rect 10876 27888 10928 27940
rect 20720 28024 20772 28076
rect 31300 28024 31352 28076
rect 36176 28024 36228 28076
rect 14372 27956 14424 28008
rect 14556 27999 14608 28008
rect 14556 27965 14565 27999
rect 14565 27965 14599 27999
rect 14599 27965 14608 27999
rect 14556 27956 14608 27965
rect 15752 27956 15804 28008
rect 16212 27999 16264 28008
rect 16212 27965 16221 27999
rect 16221 27965 16255 27999
rect 16255 27965 16264 27999
rect 16212 27956 16264 27965
rect 18144 27956 18196 28008
rect 15660 27888 15712 27940
rect 15844 27888 15896 27940
rect 21088 27956 21140 28008
rect 27620 27999 27672 28008
rect 27620 27965 27629 27999
rect 27629 27965 27663 27999
rect 27663 27965 27672 27999
rect 27620 27956 27672 27965
rect 28908 27956 28960 28008
rect 29644 27956 29696 28008
rect 31116 27956 31168 28008
rect 31668 27956 31720 28008
rect 34796 27956 34848 28008
rect 22836 27888 22888 27940
rect 12900 27820 12952 27872
rect 26240 27888 26292 27940
rect 24952 27820 25004 27872
rect 25044 27820 25096 27872
rect 26976 27820 27028 27872
rect 29368 27863 29420 27872
rect 29368 27829 29377 27863
rect 29377 27829 29411 27863
rect 29411 27829 29420 27863
rect 29368 27820 29420 27829
rect 33416 27820 33468 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 10416 27616 10468 27668
rect 10876 27616 10928 27668
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 14740 27616 14792 27668
rect 25320 27616 25372 27668
rect 27712 27616 27764 27668
rect 28356 27616 28408 27668
rect 31392 27616 31444 27668
rect 32864 27616 32916 27668
rect 11152 27480 11204 27532
rect 23388 27548 23440 27600
rect 26332 27548 26384 27600
rect 24400 27480 24452 27532
rect 27620 27480 27672 27532
rect 30012 27480 30064 27532
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 9220 27412 9272 27464
rect 10600 27412 10652 27464
rect 12808 27412 12860 27464
rect 14004 27412 14056 27464
rect 14280 27412 14332 27464
rect 11980 27387 12032 27396
rect 11980 27353 11989 27387
rect 11989 27353 12023 27387
rect 12023 27353 12032 27387
rect 12532 27387 12584 27396
rect 11980 27344 12032 27353
rect 12532 27353 12541 27387
rect 12541 27353 12575 27387
rect 12575 27353 12584 27387
rect 12532 27344 12584 27353
rect 15200 27455 15252 27464
rect 15200 27421 15209 27455
rect 15209 27421 15243 27455
rect 15243 27421 15252 27455
rect 15200 27412 15252 27421
rect 24584 27412 24636 27464
rect 28908 27412 28960 27464
rect 31668 27480 31720 27532
rect 34796 27480 34848 27532
rect 31760 27412 31812 27464
rect 6828 27276 6880 27328
rect 10416 27319 10468 27328
rect 10416 27285 10425 27319
rect 10425 27285 10459 27319
rect 10459 27285 10468 27319
rect 10416 27276 10468 27285
rect 12164 27276 12216 27328
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 16856 27387 16908 27396
rect 15936 27344 15988 27353
rect 16856 27353 16865 27387
rect 16865 27353 16899 27387
rect 16899 27353 16908 27387
rect 16856 27344 16908 27353
rect 20076 27344 20128 27396
rect 23296 27344 23348 27396
rect 25044 27344 25096 27396
rect 25688 27344 25740 27396
rect 27712 27344 27764 27396
rect 16764 27276 16816 27328
rect 20628 27276 20680 27328
rect 29092 27319 29144 27328
rect 29092 27285 29101 27319
rect 29101 27285 29135 27319
rect 29135 27285 29144 27319
rect 29092 27276 29144 27285
rect 30012 27387 30064 27396
rect 30012 27353 30021 27387
rect 30021 27353 30055 27387
rect 30055 27353 30064 27387
rect 30012 27344 30064 27353
rect 31484 27344 31536 27396
rect 33232 27276 33284 27328
rect 37556 27344 37608 27396
rect 35900 27276 35952 27328
rect 36636 27319 36688 27328
rect 36636 27285 36645 27319
rect 36645 27285 36679 27319
rect 36679 27285 36688 27319
rect 36636 27276 36688 27285
rect 37648 27319 37700 27328
rect 37648 27285 37657 27319
rect 37657 27285 37691 27319
rect 37691 27285 37700 27319
rect 37648 27276 37700 27285
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9220 27115 9272 27124
rect 9220 27081 9229 27115
rect 9229 27081 9263 27115
rect 9263 27081 9272 27115
rect 9220 27072 9272 27081
rect 14188 27072 14240 27124
rect 15200 27004 15252 27056
rect 9404 26979 9456 26988
rect 9404 26945 9413 26979
rect 9413 26945 9447 26979
rect 9447 26945 9456 26979
rect 9404 26936 9456 26945
rect 11152 26936 11204 26988
rect 11980 26979 12032 26988
rect 11980 26945 11989 26979
rect 11989 26945 12023 26979
rect 12023 26945 12032 26979
rect 11980 26936 12032 26945
rect 12716 26936 12768 26988
rect 13544 26936 13596 26988
rect 18144 26979 18196 26988
rect 18144 26945 18153 26979
rect 18153 26945 18187 26979
rect 18187 26945 18196 26979
rect 18144 26936 18196 26945
rect 23020 27072 23072 27124
rect 23664 27004 23716 27056
rect 24584 27072 24636 27124
rect 25136 27047 25188 27056
rect 25136 27013 25145 27047
rect 25145 27013 25179 27047
rect 25179 27013 25188 27047
rect 25136 27004 25188 27013
rect 26516 27004 26568 27056
rect 27620 27072 27672 27124
rect 28908 27072 28960 27124
rect 27896 27004 27948 27056
rect 30656 27072 30708 27124
rect 36636 27072 36688 27124
rect 31024 27004 31076 27056
rect 34428 27004 34480 27056
rect 31668 26936 31720 26988
rect 15108 26868 15160 26920
rect 19156 26868 19208 26920
rect 19432 26868 19484 26920
rect 20996 26868 21048 26920
rect 22376 26868 22428 26920
rect 23296 26868 23348 26920
rect 12072 26775 12124 26784
rect 12072 26741 12081 26775
rect 12081 26741 12115 26775
rect 12115 26741 12124 26775
rect 12072 26732 12124 26741
rect 12716 26775 12768 26784
rect 12716 26741 12725 26775
rect 12725 26741 12759 26775
rect 12759 26741 12768 26775
rect 12716 26732 12768 26741
rect 25872 26868 25924 26920
rect 26332 26868 26384 26920
rect 29000 26868 29052 26920
rect 29368 26868 29420 26920
rect 29828 26868 29880 26920
rect 31760 26868 31812 26920
rect 33600 26868 33652 26920
rect 24400 26732 24452 26784
rect 27068 26800 27120 26852
rect 26700 26732 26752 26784
rect 28908 26775 28960 26784
rect 28908 26741 28917 26775
rect 28917 26741 28951 26775
rect 28951 26741 28960 26775
rect 28908 26732 28960 26741
rect 31208 26775 31260 26784
rect 31208 26741 31217 26775
rect 31217 26741 31251 26775
rect 31251 26741 31260 26775
rect 31208 26732 31260 26741
rect 34704 26732 34756 26784
rect 35440 26732 35492 26784
rect 38200 26732 38252 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9772 26571 9824 26580
rect 9772 26537 9781 26571
rect 9781 26537 9815 26571
rect 9815 26537 9824 26571
rect 9772 26528 9824 26537
rect 13544 26571 13596 26580
rect 13544 26537 13553 26571
rect 13553 26537 13587 26571
rect 13587 26537 13596 26571
rect 13544 26528 13596 26537
rect 15568 26571 15620 26580
rect 15568 26537 15577 26571
rect 15577 26537 15611 26571
rect 15611 26537 15620 26571
rect 15568 26528 15620 26537
rect 17960 26528 18012 26580
rect 6736 26460 6788 26512
rect 11980 26460 12032 26512
rect 19340 26460 19392 26512
rect 24860 26528 24912 26580
rect 25320 26528 25372 26580
rect 29000 26528 29052 26580
rect 29184 26528 29236 26580
rect 10324 26392 10376 26444
rect 14372 26435 14424 26444
rect 1768 26367 1820 26376
rect 1768 26333 1777 26367
rect 1777 26333 1811 26367
rect 1811 26333 1820 26367
rect 1768 26324 1820 26333
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 10324 26299 10376 26308
rect 10324 26265 10333 26299
rect 10333 26265 10367 26299
rect 10367 26265 10376 26299
rect 10324 26256 10376 26265
rect 10416 26299 10468 26308
rect 10416 26265 10425 26299
rect 10425 26265 10459 26299
rect 10459 26265 10468 26299
rect 10416 26256 10468 26265
rect 12440 26256 12492 26308
rect 14372 26401 14381 26435
rect 14381 26401 14415 26435
rect 14415 26401 14424 26435
rect 14372 26392 14424 26401
rect 14464 26392 14516 26444
rect 25872 26460 25924 26512
rect 30380 26460 30432 26512
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 19340 26324 19392 26376
rect 23020 26392 23072 26444
rect 24584 26435 24636 26444
rect 24584 26401 24593 26435
rect 24593 26401 24627 26435
rect 24627 26401 24636 26435
rect 24584 26392 24636 26401
rect 25596 26392 25648 26444
rect 29092 26392 29144 26444
rect 30932 26392 30984 26444
rect 21272 26324 21324 26376
rect 30564 26367 30616 26376
rect 30564 26333 30573 26367
rect 30573 26333 30607 26367
rect 30607 26333 30616 26367
rect 30564 26324 30616 26333
rect 34796 26392 34848 26444
rect 38936 26460 38988 26512
rect 38476 26392 38528 26444
rect 13912 26256 13964 26308
rect 20260 26256 20312 26308
rect 22192 26188 22244 26240
rect 26240 26256 26292 26308
rect 26424 26256 26476 26308
rect 30104 26256 30156 26308
rect 30932 26256 30984 26308
rect 32128 26256 32180 26308
rect 36544 26256 36596 26308
rect 38200 26299 38252 26308
rect 26884 26188 26936 26240
rect 37004 26188 37056 26240
rect 38200 26265 38209 26299
rect 38209 26265 38243 26299
rect 38243 26265 38252 26299
rect 38200 26256 38252 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9312 25984 9364 26036
rect 12256 25984 12308 26036
rect 14464 25984 14516 26036
rect 12072 25916 12124 25968
rect 14188 25916 14240 25968
rect 15660 25916 15712 25968
rect 5448 25848 5500 25900
rect 7748 25848 7800 25900
rect 11152 25848 11204 25900
rect 11980 25848 12032 25900
rect 13820 25848 13872 25900
rect 15108 25848 15160 25900
rect 10508 25823 10560 25832
rect 10508 25789 10517 25823
rect 10517 25789 10551 25823
rect 10551 25789 10560 25823
rect 10508 25780 10560 25789
rect 8944 25712 8996 25764
rect 13268 25823 13320 25832
rect 13268 25789 13277 25823
rect 13277 25789 13311 25823
rect 13311 25789 13320 25823
rect 13268 25780 13320 25789
rect 11060 25755 11112 25764
rect 11060 25721 11069 25755
rect 11069 25721 11103 25755
rect 11103 25721 11112 25755
rect 11060 25712 11112 25721
rect 12164 25712 12216 25764
rect 4988 25687 5040 25696
rect 4988 25653 4997 25687
rect 4997 25653 5031 25687
rect 5031 25653 5040 25687
rect 4988 25644 5040 25653
rect 16764 25712 16816 25764
rect 14648 25644 14700 25696
rect 21732 25984 21784 26036
rect 21180 25916 21232 25968
rect 30012 25916 30064 25968
rect 33876 25984 33928 26036
rect 34704 25916 34756 25968
rect 37096 25916 37148 25968
rect 22100 25848 22152 25900
rect 24400 25848 24452 25900
rect 30564 25848 30616 25900
rect 31668 25848 31720 25900
rect 33692 25848 33744 25900
rect 38292 25891 38344 25900
rect 38292 25857 38301 25891
rect 38301 25857 38335 25891
rect 38335 25857 38344 25891
rect 38292 25848 38344 25857
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 19064 25780 19116 25832
rect 19340 25823 19392 25832
rect 19340 25789 19349 25823
rect 19349 25789 19383 25823
rect 19383 25789 19392 25823
rect 19340 25780 19392 25789
rect 20168 25780 20220 25832
rect 22284 25780 22336 25832
rect 24032 25712 24084 25764
rect 29092 25780 29144 25832
rect 30748 25823 30800 25832
rect 30748 25789 30757 25823
rect 30757 25789 30791 25823
rect 30791 25789 30800 25823
rect 30748 25780 30800 25789
rect 34612 25712 34664 25764
rect 32312 25644 32364 25696
rect 33876 25644 33928 25696
rect 36820 25644 36872 25696
rect 39304 25644 39356 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7748 25483 7800 25492
rect 7748 25449 7757 25483
rect 7757 25449 7791 25483
rect 7791 25449 7800 25483
rect 7748 25440 7800 25449
rect 9772 25483 9824 25492
rect 9772 25449 9781 25483
rect 9781 25449 9815 25483
rect 9815 25449 9824 25483
rect 9772 25440 9824 25449
rect 14372 25483 14424 25492
rect 14372 25449 14381 25483
rect 14381 25449 14415 25483
rect 14415 25449 14424 25483
rect 14372 25440 14424 25449
rect 15384 25440 15436 25492
rect 16764 25440 16816 25492
rect 20904 25440 20956 25492
rect 8668 25372 8720 25424
rect 7104 25279 7156 25288
rect 7104 25245 7113 25279
rect 7113 25245 7147 25279
rect 7147 25245 7156 25279
rect 7104 25236 7156 25245
rect 10232 25372 10284 25424
rect 20720 25372 20772 25424
rect 37004 25483 37056 25492
rect 37004 25449 37013 25483
rect 37013 25449 37047 25483
rect 37047 25449 37056 25483
rect 37004 25440 37056 25449
rect 26884 25372 26936 25424
rect 19340 25304 19392 25356
rect 22284 25347 22336 25356
rect 22284 25313 22293 25347
rect 22293 25313 22327 25347
rect 22327 25313 22336 25347
rect 22284 25304 22336 25313
rect 25228 25304 25280 25356
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 17868 25236 17920 25288
rect 22192 25236 22244 25288
rect 32312 25236 32364 25288
rect 36912 25279 36964 25288
rect 36912 25245 36921 25279
rect 36921 25245 36955 25279
rect 36955 25245 36964 25279
rect 36912 25236 36964 25245
rect 10416 25168 10468 25220
rect 11612 25211 11664 25220
rect 11612 25177 11621 25211
rect 11621 25177 11655 25211
rect 11655 25177 11664 25211
rect 11612 25168 11664 25177
rect 11704 25211 11756 25220
rect 11704 25177 11713 25211
rect 11713 25177 11747 25211
rect 11747 25177 11756 25211
rect 12256 25211 12308 25220
rect 11704 25168 11756 25177
rect 12256 25177 12265 25211
rect 12265 25177 12299 25211
rect 12299 25177 12308 25211
rect 12256 25168 12308 25177
rect 6644 25100 6696 25152
rect 13636 25100 13688 25152
rect 13728 25100 13780 25152
rect 15108 25211 15160 25220
rect 15108 25177 15117 25211
rect 15117 25177 15151 25211
rect 15151 25177 15160 25211
rect 15108 25168 15160 25177
rect 16396 25168 16448 25220
rect 19708 25211 19760 25220
rect 19708 25177 19717 25211
rect 19717 25177 19751 25211
rect 19751 25177 19760 25211
rect 19708 25168 19760 25177
rect 20996 25168 21048 25220
rect 21456 25211 21508 25220
rect 21456 25177 21465 25211
rect 21465 25177 21499 25211
rect 21499 25177 21508 25211
rect 21456 25168 21508 25177
rect 21824 25168 21876 25220
rect 24584 25168 24636 25220
rect 24952 25168 25004 25220
rect 25872 25168 25924 25220
rect 29736 25168 29788 25220
rect 16028 25100 16080 25152
rect 16488 25100 16540 25152
rect 20536 25100 20588 25152
rect 22192 25100 22244 25152
rect 22652 25100 22704 25152
rect 24032 25100 24084 25152
rect 26332 25143 26384 25152
rect 26332 25109 26341 25143
rect 26341 25109 26375 25143
rect 26375 25109 26384 25143
rect 26332 25100 26384 25109
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 10416 24896 10468 24948
rect 22376 24896 22428 24948
rect 12348 24871 12400 24880
rect 4988 24760 5040 24812
rect 8392 24760 8444 24812
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 8668 24760 8720 24769
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10416 24692 10468 24701
rect 10968 24667 11020 24676
rect 10968 24633 10977 24667
rect 10977 24633 11011 24667
rect 11011 24633 11020 24667
rect 10968 24624 11020 24633
rect 12348 24837 12357 24871
rect 12357 24837 12391 24871
rect 12391 24837 12400 24871
rect 12348 24828 12400 24837
rect 14648 24871 14700 24880
rect 14648 24837 14657 24871
rect 14657 24837 14691 24871
rect 14691 24837 14700 24871
rect 14648 24828 14700 24837
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 16488 24828 16540 24880
rect 13912 24760 13964 24769
rect 15936 24760 15988 24812
rect 17132 24760 17184 24812
rect 19340 24828 19392 24880
rect 19708 24828 19760 24880
rect 22284 24760 22336 24812
rect 23204 24828 23256 24880
rect 24400 24828 24452 24880
rect 11888 24692 11940 24744
rect 12348 24692 12400 24744
rect 12808 24735 12860 24744
rect 12808 24701 12817 24735
rect 12817 24701 12851 24735
rect 12851 24701 12860 24735
rect 12808 24692 12860 24701
rect 14832 24692 14884 24744
rect 19984 24692 20036 24744
rect 12716 24624 12768 24676
rect 16580 24624 16632 24676
rect 20812 24624 20864 24676
rect 28816 24760 28868 24812
rect 30840 24760 30892 24812
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 38292 24760 38344 24812
rect 23480 24692 23532 24744
rect 25228 24692 25280 24744
rect 27160 24735 27212 24744
rect 27160 24701 27169 24735
rect 27169 24701 27203 24735
rect 27203 24701 27212 24735
rect 27160 24692 27212 24701
rect 27436 24735 27488 24744
rect 27436 24701 27445 24735
rect 27445 24701 27479 24735
rect 27479 24701 27488 24735
rect 27436 24692 27488 24701
rect 29460 24735 29512 24744
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 7288 24556 7340 24608
rect 9312 24556 9364 24608
rect 19432 24556 19484 24608
rect 22100 24556 22152 24608
rect 26700 24556 26752 24608
rect 27160 24556 27212 24608
rect 29460 24701 29469 24735
rect 29469 24701 29503 24735
rect 29503 24701 29512 24735
rect 29460 24692 29512 24701
rect 28540 24624 28592 24676
rect 28724 24624 28776 24676
rect 30196 24692 30248 24744
rect 29000 24556 29052 24608
rect 33876 24692 33928 24744
rect 34060 24735 34112 24744
rect 34060 24701 34069 24735
rect 34069 24701 34103 24735
rect 34103 24701 34112 24735
rect 34060 24692 34112 24701
rect 36452 24556 36504 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8392 24352 8444 24404
rect 11612 24352 11664 24404
rect 11704 24352 11756 24404
rect 13728 24284 13780 24336
rect 9312 24259 9364 24268
rect 9312 24225 9321 24259
rect 9321 24225 9355 24259
rect 9355 24225 9364 24259
rect 9312 24216 9364 24225
rect 11336 24216 11388 24268
rect 7288 24191 7340 24200
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 7288 24157 7297 24191
rect 7297 24157 7331 24191
rect 7331 24157 7340 24191
rect 7288 24148 7340 24157
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 13176 24080 13228 24132
rect 22100 24352 22152 24404
rect 22284 24352 22336 24404
rect 24400 24352 24452 24404
rect 32128 24352 32180 24404
rect 32404 24352 32456 24404
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 14188 24284 14240 24336
rect 19064 24284 19116 24336
rect 16304 24216 16356 24268
rect 19616 24216 19668 24268
rect 19708 24216 19760 24268
rect 20812 24216 20864 24268
rect 24860 24216 24912 24268
rect 32312 24216 32364 24268
rect 34244 24216 34296 24268
rect 36176 24216 36228 24268
rect 14004 24148 14056 24200
rect 14188 24148 14240 24200
rect 19248 24080 19300 24132
rect 14004 24012 14056 24064
rect 16488 24012 16540 24064
rect 19432 24012 19484 24064
rect 29460 24148 29512 24200
rect 31576 24148 31628 24200
rect 34796 24148 34848 24200
rect 37464 24191 37516 24200
rect 37464 24157 37473 24191
rect 37473 24157 37507 24191
rect 37507 24157 37516 24191
rect 37464 24148 37516 24157
rect 38108 24148 38160 24200
rect 20352 24123 20404 24132
rect 20352 24089 20361 24123
rect 20361 24089 20395 24123
rect 20395 24089 20404 24123
rect 20352 24080 20404 24089
rect 23296 24080 23348 24132
rect 24676 24123 24728 24132
rect 24676 24089 24685 24123
rect 24685 24089 24719 24123
rect 24719 24089 24728 24123
rect 24676 24080 24728 24089
rect 20996 24012 21048 24064
rect 21088 24012 21140 24064
rect 21824 24055 21876 24064
rect 21824 24021 21833 24055
rect 21833 24021 21867 24055
rect 21867 24021 21876 24055
rect 21824 24012 21876 24021
rect 21916 24012 21968 24064
rect 31116 24012 31168 24064
rect 34428 24080 34480 24132
rect 39488 24080 39540 24132
rect 35440 24012 35492 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 12440 23740 12492 23792
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 12256 23647 12308 23656
rect 12256 23613 12265 23647
rect 12265 23613 12299 23647
rect 12299 23613 12308 23647
rect 12256 23604 12308 23613
rect 17960 23604 18012 23656
rect 13176 23536 13228 23588
rect 19340 23808 19392 23860
rect 23388 23808 23440 23860
rect 25228 23808 25280 23860
rect 26976 23808 27028 23860
rect 19432 23740 19484 23792
rect 20996 23740 21048 23792
rect 28172 23740 28224 23792
rect 30380 23740 30432 23792
rect 36912 23808 36964 23860
rect 37556 23851 37608 23860
rect 37556 23817 37565 23851
rect 37565 23817 37599 23851
rect 37599 23817 37608 23851
rect 37556 23808 37608 23817
rect 22468 23672 22520 23724
rect 23388 23715 23440 23724
rect 23388 23681 23397 23715
rect 23397 23681 23431 23715
rect 23431 23681 23440 23715
rect 23388 23672 23440 23681
rect 27160 23672 27212 23724
rect 29460 23672 29512 23724
rect 32312 23672 32364 23724
rect 34796 23740 34848 23792
rect 37648 23740 37700 23792
rect 36452 23715 36504 23724
rect 36452 23681 36461 23715
rect 36461 23681 36495 23715
rect 36495 23681 36504 23715
rect 36452 23672 36504 23681
rect 39764 23672 39816 23724
rect 21640 23604 21692 23656
rect 21824 23604 21876 23656
rect 25136 23604 25188 23656
rect 26332 23604 26384 23656
rect 28264 23604 28316 23656
rect 28908 23604 28960 23656
rect 30104 23647 30156 23656
rect 30104 23613 30113 23647
rect 30113 23613 30147 23647
rect 30147 23613 30156 23647
rect 30104 23604 30156 23613
rect 34336 23604 34388 23656
rect 12716 23468 12768 23520
rect 18604 23468 18656 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 25596 23536 25648 23588
rect 27620 23536 27672 23588
rect 29276 23536 29328 23588
rect 21456 23468 21508 23520
rect 23756 23468 23808 23520
rect 28540 23468 28592 23520
rect 31392 23468 31444 23520
rect 32956 23468 33008 23520
rect 34520 23468 34572 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 9128 23264 9180 23316
rect 12440 23307 12492 23316
rect 12440 23273 12449 23307
rect 12449 23273 12483 23307
rect 12483 23273 12492 23307
rect 12440 23264 12492 23273
rect 15108 23264 15160 23316
rect 19432 23264 19484 23316
rect 20076 23264 20128 23316
rect 19892 23196 19944 23248
rect 8852 23060 8904 23112
rect 9312 23103 9364 23112
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 14924 23128 14976 23180
rect 19340 23128 19392 23180
rect 20720 23171 20772 23180
rect 12992 23060 13044 23112
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 17408 23060 17460 23112
rect 19892 23060 19944 23112
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 20720 23128 20772 23137
rect 22836 23264 22888 23316
rect 23756 23264 23808 23316
rect 24216 23264 24268 23316
rect 31116 23264 31168 23316
rect 27620 23196 27672 23248
rect 29368 23128 29420 23180
rect 29460 23128 29512 23180
rect 32312 23128 32364 23180
rect 34796 23128 34848 23180
rect 24768 23060 24820 23112
rect 25228 23103 25280 23112
rect 25228 23069 25237 23103
rect 25237 23069 25271 23103
rect 25271 23069 25280 23103
rect 25228 23060 25280 23069
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 37464 23060 37516 23112
rect 19984 22992 20036 23044
rect 11888 22924 11940 22976
rect 17868 22924 17920 22976
rect 20536 22924 20588 22976
rect 23480 23035 23532 23044
rect 23480 23001 23489 23035
rect 23489 23001 23523 23035
rect 23523 23001 23532 23035
rect 25504 23035 25556 23044
rect 23480 22992 23532 23001
rect 25504 23001 25513 23035
rect 25513 23001 25547 23035
rect 25547 23001 25556 23035
rect 25504 22992 25556 23001
rect 27528 22992 27580 23044
rect 31852 22992 31904 23044
rect 35072 22992 35124 23044
rect 25044 22924 25096 22976
rect 26424 22924 26476 22976
rect 26792 22924 26844 22976
rect 32680 22924 32732 22976
rect 37004 22992 37056 23044
rect 36636 22967 36688 22976
rect 36636 22933 36645 22967
rect 36645 22933 36679 22967
rect 36679 22933 36688 22967
rect 36636 22924 36688 22933
rect 37280 22924 37332 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 12348 22695 12400 22704
rect 12348 22661 12357 22695
rect 12357 22661 12391 22695
rect 12391 22661 12400 22695
rect 12348 22652 12400 22661
rect 14740 22720 14792 22772
rect 15016 22720 15068 22772
rect 20076 22720 20128 22772
rect 20536 22720 20588 22772
rect 24124 22720 24176 22772
rect 25596 22720 25648 22772
rect 14004 22695 14056 22704
rect 14004 22661 14013 22695
rect 14013 22661 14047 22695
rect 14047 22661 14056 22695
rect 14004 22652 14056 22661
rect 18236 22652 18288 22704
rect 18788 22695 18840 22704
rect 18788 22661 18797 22695
rect 18797 22661 18831 22695
rect 18831 22661 18840 22695
rect 18788 22652 18840 22661
rect 22008 22652 22060 22704
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 7288 22584 7340 22636
rect 9220 22584 9272 22636
rect 11704 22584 11756 22636
rect 15292 22584 15344 22636
rect 21364 22584 21416 22636
rect 24860 22652 24912 22704
rect 26148 22720 26200 22772
rect 31116 22720 31168 22772
rect 30472 22652 30524 22704
rect 31852 22652 31904 22704
rect 36084 22720 36136 22772
rect 36452 22720 36504 22772
rect 37188 22652 37240 22704
rect 25780 22584 25832 22636
rect 27160 22627 27212 22636
rect 11060 22516 11112 22568
rect 11612 22516 11664 22568
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 14372 22516 14424 22568
rect 14924 22559 14976 22568
rect 14924 22525 14933 22559
rect 14933 22525 14967 22559
rect 14967 22525 14976 22559
rect 14924 22516 14976 22525
rect 19340 22516 19392 22568
rect 23572 22516 23624 22568
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 29460 22584 29512 22636
rect 34244 22584 34296 22636
rect 34796 22627 34848 22636
rect 34796 22593 34805 22627
rect 34805 22593 34839 22627
rect 34839 22593 34848 22627
rect 34796 22584 34848 22593
rect 37556 22584 37608 22636
rect 9128 22448 9180 22500
rect 14832 22448 14884 22500
rect 20260 22491 20312 22500
rect 20260 22457 20269 22491
rect 20269 22457 20303 22491
rect 20303 22457 20312 22491
rect 20260 22448 20312 22457
rect 21272 22448 21324 22500
rect 26608 22516 26660 22568
rect 30196 22559 30248 22568
rect 29828 22448 29880 22500
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 17316 22380 17368 22432
rect 18604 22380 18656 22432
rect 20720 22380 20772 22432
rect 24124 22380 24176 22432
rect 30196 22525 30205 22559
rect 30205 22525 30239 22559
rect 30239 22525 30248 22559
rect 30196 22516 30248 22525
rect 30564 22516 30616 22568
rect 32312 22559 32364 22568
rect 32312 22525 32321 22559
rect 32321 22525 32355 22559
rect 32355 22525 32364 22559
rect 32312 22516 32364 22525
rect 32680 22516 32732 22568
rect 35440 22516 35492 22568
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 34336 22380 34388 22432
rect 35624 22380 35676 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 9312 22176 9364 22228
rect 14832 22176 14884 22228
rect 15016 22176 15068 22228
rect 15752 22176 15804 22228
rect 15936 22176 15988 22228
rect 25504 22176 25556 22228
rect 26792 22176 26844 22228
rect 32220 22176 32272 22228
rect 32404 22176 32456 22228
rect 21456 22108 21508 22160
rect 25136 22108 25188 22160
rect 7748 22040 7800 22092
rect 11244 22040 11296 22092
rect 12072 22083 12124 22092
rect 12072 22049 12081 22083
rect 12081 22049 12115 22083
rect 12115 22049 12124 22083
rect 12072 22040 12124 22049
rect 18880 22040 18932 22092
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 6828 21972 6880 22024
rect 6644 21904 6696 21956
rect 11428 21972 11480 22024
rect 14372 21947 14424 21956
rect 1584 21836 1636 21888
rect 6828 21836 6880 21888
rect 10876 21836 10928 21888
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 15292 21904 15344 21956
rect 16580 21972 16632 22024
rect 17408 21972 17460 22024
rect 21732 21972 21784 22024
rect 31300 22108 31352 22160
rect 22836 21904 22888 21956
rect 24768 21904 24820 21956
rect 26608 22040 26660 22092
rect 32312 22040 32364 22092
rect 36636 22176 36688 22228
rect 37004 22176 37056 22228
rect 39856 22108 39908 22160
rect 27988 21972 28040 22024
rect 29920 21972 29972 22024
rect 27436 21904 27488 21956
rect 32956 21904 33008 21956
rect 34796 22040 34848 22092
rect 35624 22040 35676 22092
rect 37464 21972 37516 22024
rect 11980 21836 12032 21888
rect 17224 21836 17276 21888
rect 17408 21836 17460 21888
rect 23940 21836 23992 21888
rect 24308 21836 24360 21888
rect 25872 21836 25924 21888
rect 28724 21836 28776 21888
rect 29920 21836 29972 21888
rect 33784 21836 33836 21888
rect 37004 21904 37056 21956
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 37832 21836 37884 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 14740 21675 14792 21684
rect 14740 21641 14749 21675
rect 14749 21641 14783 21675
rect 14783 21641 14792 21675
rect 14740 21632 14792 21641
rect 15292 21632 15344 21684
rect 20536 21632 20588 21684
rect 20904 21632 20956 21684
rect 22468 21632 22520 21684
rect 24400 21632 24452 21684
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 25872 21632 25924 21684
rect 11060 21564 11112 21616
rect 17224 21564 17276 21616
rect 1584 21539 1636 21548
rect 1584 21505 1593 21539
rect 1593 21505 1627 21539
rect 1627 21505 1636 21539
rect 1584 21496 1636 21505
rect 6736 21496 6788 21548
rect 12532 21496 12584 21548
rect 20352 21496 20404 21548
rect 23296 21564 23348 21616
rect 33968 21632 34020 21684
rect 28080 21564 28132 21616
rect 28908 21607 28960 21616
rect 28908 21573 28917 21607
rect 28917 21573 28951 21607
rect 28951 21573 28960 21607
rect 28908 21564 28960 21573
rect 34244 21564 34296 21616
rect 35440 21564 35492 21616
rect 37280 21564 37332 21616
rect 24308 21496 24360 21548
rect 24860 21496 24912 21548
rect 25596 21496 25648 21548
rect 27068 21496 27120 21548
rect 10140 21428 10192 21480
rect 10876 21428 10928 21480
rect 17868 21428 17920 21480
rect 22008 21428 22060 21480
rect 34336 21496 34388 21548
rect 34612 21496 34664 21548
rect 34796 21496 34848 21548
rect 27988 21428 28040 21480
rect 23112 21360 23164 21412
rect 23572 21360 23624 21412
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 16948 21292 17000 21344
rect 21180 21292 21232 21344
rect 26424 21292 26476 21344
rect 27620 21360 27672 21412
rect 29828 21428 29880 21480
rect 31392 21428 31444 21480
rect 37280 21428 37332 21480
rect 29368 21403 29420 21412
rect 29368 21369 29377 21403
rect 29377 21369 29411 21403
rect 29411 21369 29420 21403
rect 29368 21360 29420 21369
rect 29736 21360 29788 21412
rect 30656 21360 30708 21412
rect 31852 21360 31904 21412
rect 34336 21360 34388 21412
rect 37004 21360 37056 21412
rect 37740 21360 37792 21412
rect 33968 21292 34020 21344
rect 36176 21292 36228 21344
rect 36636 21335 36688 21344
rect 36636 21301 36645 21335
rect 36645 21301 36679 21335
rect 36679 21301 36688 21335
rect 36636 21292 36688 21301
rect 38292 21292 38344 21344
rect 39672 21292 39724 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 39672 21156 39724 21208
rect 9220 21088 9272 21140
rect 11428 21088 11480 21140
rect 19432 21088 19484 21140
rect 21916 21088 21968 21140
rect 23388 21088 23440 21140
rect 25044 21088 25096 21140
rect 26148 21088 26200 21140
rect 26424 21088 26476 21140
rect 30840 21088 30892 21140
rect 33968 21131 34020 21140
rect 33968 21097 33977 21131
rect 33977 21097 34011 21131
rect 34011 21097 34020 21131
rect 33968 21088 34020 21097
rect 35900 21131 35952 21140
rect 35900 21097 35909 21131
rect 35909 21097 35943 21131
rect 35943 21097 35952 21131
rect 35900 21088 35952 21097
rect 37280 21088 37332 21140
rect 37464 21088 37516 21140
rect 39580 21088 39632 21140
rect 3424 21020 3476 21072
rect 23940 21063 23992 21072
rect 21272 20952 21324 21004
rect 23940 21029 23949 21063
rect 23949 21029 23983 21063
rect 23983 21029 23992 21063
rect 23940 21020 23992 21029
rect 25412 21020 25464 21072
rect 27344 21020 27396 21072
rect 28448 20995 28500 21004
rect 28448 20961 28457 20995
rect 28457 20961 28491 20995
rect 28491 20961 28500 20995
rect 28448 20952 28500 20961
rect 30748 20952 30800 21004
rect 33140 21020 33192 21072
rect 33876 21020 33928 21072
rect 34244 21020 34296 21072
rect 34428 21020 34480 21072
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 16488 20927 16540 20936
rect 16488 20893 16497 20927
rect 16497 20893 16531 20927
rect 16531 20893 16540 20927
rect 16488 20884 16540 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 15200 20748 15252 20800
rect 17132 20748 17184 20800
rect 17316 20859 17368 20868
rect 17316 20825 17325 20859
rect 17325 20825 17359 20859
rect 17359 20825 17368 20859
rect 17316 20816 17368 20825
rect 19248 20816 19300 20868
rect 22192 20884 22244 20936
rect 22652 20816 22704 20868
rect 23112 20816 23164 20868
rect 23664 20816 23716 20868
rect 24124 20816 24176 20868
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 19432 20748 19484 20800
rect 20352 20748 20404 20800
rect 22928 20748 22980 20800
rect 24860 20816 24912 20868
rect 25872 20884 25924 20936
rect 26332 20884 26384 20936
rect 26608 20884 26660 20936
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 29000 20816 29052 20868
rect 29552 20816 29604 20868
rect 28448 20748 28500 20800
rect 30840 20748 30892 20800
rect 31668 20952 31720 21004
rect 37464 20952 37516 21004
rect 38108 20952 38160 21004
rect 38752 20952 38804 21004
rect 32128 20927 32180 20936
rect 32128 20893 32137 20927
rect 32137 20893 32171 20927
rect 32171 20893 32180 20927
rect 32128 20884 32180 20893
rect 32496 20884 32548 20936
rect 33508 20884 33560 20936
rect 33784 20884 33836 20936
rect 33876 20927 33928 20936
rect 33876 20893 33885 20927
rect 33885 20893 33919 20927
rect 33919 20893 33928 20927
rect 33876 20884 33928 20893
rect 34152 20884 34204 20936
rect 35992 20884 36044 20936
rect 36452 20927 36504 20936
rect 36452 20893 36461 20927
rect 36461 20893 36495 20927
rect 36495 20893 36504 20927
rect 36452 20884 36504 20893
rect 34796 20816 34848 20868
rect 37372 20859 37424 20868
rect 37372 20825 37381 20859
rect 37381 20825 37415 20859
rect 37415 20825 37424 20859
rect 37372 20816 37424 20825
rect 35164 20748 35216 20800
rect 35808 20748 35860 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 16948 20519 17000 20528
rect 16948 20485 16957 20519
rect 16957 20485 16991 20519
rect 16991 20485 17000 20519
rect 16948 20476 17000 20485
rect 18328 20476 18380 20528
rect 20996 20544 21048 20596
rect 23664 20544 23716 20596
rect 23848 20587 23900 20596
rect 23848 20553 23857 20587
rect 23857 20553 23891 20587
rect 23891 20553 23900 20587
rect 23848 20544 23900 20553
rect 24584 20544 24636 20596
rect 28908 20587 28960 20596
rect 14556 20340 14608 20392
rect 17592 20340 17644 20392
rect 26148 20519 26200 20528
rect 26148 20485 26157 20519
rect 26157 20485 26191 20519
rect 26191 20485 26200 20519
rect 26148 20476 26200 20485
rect 26424 20476 26476 20528
rect 22560 20408 22612 20460
rect 22652 20451 22704 20460
rect 22652 20417 22661 20451
rect 22661 20417 22695 20451
rect 22695 20417 22704 20451
rect 22652 20408 22704 20417
rect 22836 20408 22888 20460
rect 21824 20340 21876 20392
rect 7288 20315 7340 20324
rect 7288 20281 7297 20315
rect 7297 20281 7331 20315
rect 7331 20281 7340 20315
rect 7288 20272 7340 20281
rect 13268 20272 13320 20324
rect 13728 20272 13780 20324
rect 22100 20272 22152 20324
rect 22376 20272 22428 20324
rect 22836 20272 22888 20324
rect 23296 20340 23348 20392
rect 23572 20340 23624 20392
rect 24860 20408 24912 20460
rect 26332 20408 26384 20460
rect 25872 20340 25924 20392
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 28908 20553 28917 20587
rect 28917 20553 28951 20587
rect 28951 20553 28960 20587
rect 28908 20544 28960 20553
rect 29552 20587 29604 20596
rect 29552 20553 29561 20587
rect 29561 20553 29595 20587
rect 29595 20553 29604 20587
rect 29552 20544 29604 20553
rect 30380 20544 30432 20596
rect 33784 20544 33836 20596
rect 34152 20544 34204 20596
rect 35348 20544 35400 20596
rect 36084 20544 36136 20596
rect 38200 20587 38252 20596
rect 38200 20553 38209 20587
rect 38209 20553 38243 20587
rect 38243 20553 38252 20587
rect 38200 20544 38252 20553
rect 29184 20476 29236 20528
rect 30840 20519 30892 20528
rect 30840 20485 30849 20519
rect 30849 20485 30883 20519
rect 30883 20485 30892 20519
rect 30840 20476 30892 20485
rect 32128 20476 32180 20528
rect 29092 20408 29144 20460
rect 32404 20408 32456 20460
rect 35624 20476 35676 20528
rect 29736 20340 29788 20392
rect 30748 20383 30800 20392
rect 30748 20349 30757 20383
rect 30757 20349 30791 20383
rect 30791 20349 30800 20383
rect 30748 20340 30800 20349
rect 31852 20340 31904 20392
rect 33968 20383 34020 20392
rect 33968 20349 33977 20383
rect 33977 20349 34011 20383
rect 34011 20349 34020 20383
rect 33968 20340 34020 20349
rect 34152 20340 34204 20392
rect 36452 20408 36504 20460
rect 36728 20451 36780 20460
rect 35532 20340 35584 20392
rect 36728 20417 36737 20451
rect 36737 20417 36771 20451
rect 36771 20417 36780 20451
rect 36728 20408 36780 20417
rect 38016 20451 38068 20460
rect 38016 20417 38025 20451
rect 38025 20417 38059 20451
rect 38059 20417 38068 20451
rect 38016 20408 38068 20417
rect 11704 20204 11756 20256
rect 18144 20204 18196 20256
rect 19616 20204 19668 20256
rect 20076 20204 20128 20256
rect 32312 20204 32364 20256
rect 32496 20204 32548 20256
rect 33692 20204 33744 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 14096 20000 14148 20052
rect 21732 20000 21784 20052
rect 21824 20000 21876 20052
rect 22928 20000 22980 20052
rect 23204 20000 23256 20052
rect 23756 20000 23808 20052
rect 25964 20000 26016 20052
rect 27528 20000 27580 20052
rect 28908 20000 28960 20052
rect 32128 20000 32180 20052
rect 34152 20000 34204 20052
rect 13636 19932 13688 19984
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 19432 19932 19484 19984
rect 20076 19975 20128 19984
rect 20076 19941 20085 19975
rect 20085 19941 20119 19975
rect 20119 19941 20128 19975
rect 20076 19932 20128 19941
rect 17500 19864 17552 19916
rect 23020 19864 23072 19916
rect 27160 19864 27212 19916
rect 28172 19907 28224 19916
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 20720 19796 20772 19848
rect 21824 19796 21876 19848
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 24860 19796 24912 19848
rect 26332 19796 26384 19848
rect 11796 19771 11848 19780
rect 11796 19737 11805 19771
rect 11805 19737 11839 19771
rect 11839 19737 11848 19771
rect 11796 19728 11848 19737
rect 11888 19771 11940 19780
rect 11888 19737 11897 19771
rect 11897 19737 11931 19771
rect 11931 19737 11940 19771
rect 12808 19771 12860 19780
rect 11888 19728 11940 19737
rect 12808 19737 12817 19771
rect 12817 19737 12851 19771
rect 12851 19737 12860 19771
rect 12808 19728 12860 19737
rect 15200 19728 15252 19780
rect 17868 19728 17920 19780
rect 1860 19660 1912 19712
rect 11704 19660 11756 19712
rect 13084 19660 13136 19712
rect 19616 19771 19668 19780
rect 19616 19737 19625 19771
rect 19625 19737 19659 19771
rect 19659 19737 19668 19771
rect 26700 19771 26752 19780
rect 19616 19728 19668 19737
rect 26700 19737 26709 19771
rect 26709 19737 26743 19771
rect 26743 19737 26752 19771
rect 26700 19728 26752 19737
rect 28172 19873 28181 19907
rect 28181 19873 28215 19907
rect 28215 19873 28224 19907
rect 28172 19864 28224 19873
rect 29736 19907 29788 19916
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 29920 19907 29972 19916
rect 29920 19873 29929 19907
rect 29929 19873 29963 19907
rect 29963 19873 29972 19907
rect 29920 19864 29972 19873
rect 31852 19932 31904 19984
rect 35348 19932 35400 19984
rect 37464 19932 37516 19984
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 28448 19796 28500 19848
rect 28908 19796 28960 19848
rect 33876 19907 33928 19916
rect 33876 19873 33885 19907
rect 33885 19873 33919 19907
rect 33919 19873 33928 19907
rect 33876 19864 33928 19873
rect 35256 19907 35308 19916
rect 35256 19873 35265 19907
rect 35265 19873 35299 19907
rect 35299 19873 35308 19907
rect 35256 19864 35308 19873
rect 31668 19796 31720 19848
rect 32036 19839 32088 19848
rect 32036 19805 32045 19839
rect 32045 19805 32079 19839
rect 32079 19805 32088 19839
rect 32036 19796 32088 19805
rect 34796 19796 34848 19848
rect 35808 19864 35860 19916
rect 39396 19864 39448 19916
rect 36176 19796 36228 19848
rect 20076 19660 20128 19712
rect 20720 19703 20772 19712
rect 20720 19669 20729 19703
rect 20729 19669 20763 19703
rect 20763 19669 20772 19703
rect 20720 19660 20772 19669
rect 29460 19728 29512 19780
rect 32220 19771 32272 19780
rect 32220 19737 32229 19771
rect 32229 19737 32263 19771
rect 32263 19737 32272 19771
rect 32220 19728 32272 19737
rect 35164 19728 35216 19780
rect 35900 19728 35952 19780
rect 29092 19660 29144 19712
rect 30840 19660 30892 19712
rect 31576 19660 31628 19712
rect 33784 19660 33836 19712
rect 34428 19660 34480 19712
rect 34612 19660 34664 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 21364 19499 21416 19508
rect 21364 19465 21373 19499
rect 21373 19465 21407 19499
rect 21407 19465 21416 19499
rect 21364 19456 21416 19465
rect 21456 19456 21508 19508
rect 26240 19499 26292 19508
rect 13084 19431 13136 19440
rect 13084 19397 13093 19431
rect 13093 19397 13127 19431
rect 13127 19397 13136 19431
rect 13084 19388 13136 19397
rect 16488 19388 16540 19440
rect 16948 19431 17000 19440
rect 16948 19397 16957 19431
rect 16957 19397 16991 19431
rect 16991 19397 17000 19431
rect 16948 19388 17000 19397
rect 19156 19388 19208 19440
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 8300 19320 8352 19372
rect 12348 19320 12400 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 17868 19320 17920 19372
rect 13360 19184 13412 19236
rect 19432 19295 19484 19304
rect 19432 19261 19441 19295
rect 19441 19261 19475 19295
rect 19475 19261 19484 19295
rect 19432 19252 19484 19261
rect 20720 19388 20772 19440
rect 25964 19388 26016 19440
rect 26240 19465 26249 19499
rect 26249 19465 26283 19499
rect 26283 19465 26292 19499
rect 26240 19456 26292 19465
rect 27896 19388 27948 19440
rect 29000 19388 29052 19440
rect 30656 19431 30708 19440
rect 30656 19397 30665 19431
rect 30665 19397 30699 19431
rect 30699 19397 30708 19431
rect 30656 19388 30708 19397
rect 31576 19431 31628 19440
rect 31576 19397 31585 19431
rect 31585 19397 31619 19431
rect 31619 19397 31628 19431
rect 31576 19388 31628 19397
rect 31668 19388 31720 19440
rect 34152 19431 34204 19440
rect 34152 19397 34161 19431
rect 34161 19397 34195 19431
rect 34195 19397 34204 19431
rect 34152 19388 34204 19397
rect 34796 19431 34848 19440
rect 34796 19397 34805 19431
rect 34805 19397 34839 19431
rect 34839 19397 34848 19431
rect 34796 19388 34848 19397
rect 35256 19388 35308 19440
rect 35900 19388 35952 19440
rect 36084 19388 36136 19440
rect 21088 19320 21140 19372
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 25504 19363 25556 19372
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 25780 19320 25832 19372
rect 26240 19320 26292 19372
rect 26424 19320 26476 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27988 19363 28040 19372
rect 27988 19329 27997 19363
rect 27997 19329 28031 19363
rect 28031 19329 28040 19363
rect 27988 19320 28040 19329
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 22100 19252 22152 19261
rect 15108 19184 15160 19236
rect 28080 19252 28132 19304
rect 28356 19252 28408 19304
rect 29644 19320 29696 19372
rect 30380 19320 30432 19372
rect 32036 19320 32088 19372
rect 36176 19363 36228 19372
rect 36176 19329 36185 19363
rect 36185 19329 36219 19363
rect 36219 19329 36228 19363
rect 36176 19320 36228 19329
rect 32496 19295 32548 19304
rect 27344 19184 27396 19236
rect 27528 19184 27580 19236
rect 20076 19116 20128 19168
rect 23940 19116 23992 19168
rect 25688 19116 25740 19168
rect 29092 19116 29144 19168
rect 29920 19184 29972 19236
rect 32496 19261 32505 19295
rect 32505 19261 32539 19295
rect 32539 19261 32548 19295
rect 32496 19252 32548 19261
rect 32312 19184 32364 19236
rect 32772 19184 32824 19236
rect 31300 19116 31352 19168
rect 31668 19116 31720 19168
rect 34980 19295 35032 19304
rect 34980 19261 34989 19295
rect 34989 19261 35023 19295
rect 35023 19261 35032 19295
rect 34980 19252 35032 19261
rect 37464 19295 37516 19304
rect 37464 19261 37473 19295
rect 37473 19261 37507 19295
rect 37507 19261 37516 19295
rect 37464 19252 37516 19261
rect 34612 19184 34664 19236
rect 34152 19116 34204 19168
rect 35256 19184 35308 19236
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 14372 18912 14424 18964
rect 18328 18912 18380 18964
rect 19156 18912 19208 18964
rect 20076 18912 20128 18964
rect 20352 18912 20404 18964
rect 25136 18912 25188 18964
rect 27344 18912 27396 18964
rect 27436 18912 27488 18964
rect 30472 18912 30524 18964
rect 33232 18912 33284 18964
rect 33692 18955 33744 18964
rect 33692 18921 33701 18955
rect 33701 18921 33735 18955
rect 33735 18921 33744 18955
rect 33692 18912 33744 18921
rect 36912 18955 36964 18964
rect 36912 18921 36921 18955
rect 36921 18921 36955 18955
rect 36955 18921 36964 18955
rect 36912 18912 36964 18921
rect 37648 18912 37700 18964
rect 1676 18708 1728 18760
rect 12532 18844 12584 18896
rect 13176 18844 13228 18896
rect 15108 18887 15160 18896
rect 15108 18853 15117 18887
rect 15117 18853 15151 18887
rect 15151 18853 15160 18887
rect 15108 18844 15160 18853
rect 15568 18844 15620 18896
rect 32404 18887 32456 18896
rect 12348 18776 12400 18828
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 19524 18776 19576 18828
rect 20720 18776 20772 18828
rect 23940 18776 23992 18828
rect 26332 18776 26384 18828
rect 27160 18776 27212 18828
rect 32404 18853 32413 18887
rect 32413 18853 32447 18887
rect 32447 18853 32456 18887
rect 32404 18844 32456 18853
rect 32772 18844 32824 18896
rect 33048 18844 33100 18896
rect 34704 18844 34756 18896
rect 35716 18844 35768 18896
rect 38936 18844 38988 18896
rect 35900 18776 35952 18828
rect 35992 18776 36044 18828
rect 12624 18708 12676 18760
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 24768 18708 24820 18760
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 27068 18708 27120 18760
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 28908 18708 28960 18760
rect 30380 18751 30432 18760
rect 30380 18717 30389 18751
rect 30389 18717 30423 18751
rect 30423 18717 30432 18751
rect 30380 18708 30432 18717
rect 30472 18708 30524 18760
rect 9312 18640 9364 18692
rect 11060 18640 11112 18692
rect 13728 18640 13780 18692
rect 14648 18683 14700 18692
rect 14648 18649 14657 18683
rect 14657 18649 14691 18683
rect 14691 18649 14700 18683
rect 14648 18640 14700 18649
rect 17500 18640 17552 18692
rect 20168 18640 20220 18692
rect 20352 18640 20404 18692
rect 12164 18572 12216 18624
rect 14188 18572 14240 18624
rect 14372 18572 14424 18624
rect 25688 18640 25740 18692
rect 26884 18683 26936 18692
rect 26884 18649 26893 18683
rect 26893 18649 26927 18683
rect 26927 18649 26936 18683
rect 26884 18640 26936 18649
rect 27896 18683 27948 18692
rect 27896 18649 27905 18683
rect 27905 18649 27939 18683
rect 27939 18649 27948 18683
rect 27896 18640 27948 18649
rect 28448 18640 28500 18692
rect 28816 18640 28868 18692
rect 31576 18708 31628 18760
rect 32956 18751 33008 18760
rect 32956 18717 32965 18751
rect 32965 18717 32999 18751
rect 32999 18717 33008 18751
rect 32956 18708 33008 18717
rect 33232 18708 33284 18760
rect 38016 18708 38068 18760
rect 39580 18708 39632 18760
rect 27344 18572 27396 18624
rect 31116 18640 31168 18692
rect 32588 18640 32640 18692
rect 34612 18640 34664 18692
rect 36268 18640 36320 18692
rect 30840 18572 30892 18624
rect 31576 18572 31628 18624
rect 33876 18572 33928 18624
rect 36176 18572 36228 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 8300 18368 8352 18420
rect 14648 18368 14700 18420
rect 17500 18411 17552 18420
rect 17500 18377 17509 18411
rect 17509 18377 17543 18411
rect 17543 18377 17552 18411
rect 17500 18368 17552 18377
rect 18328 18368 18380 18420
rect 26424 18368 26476 18420
rect 26516 18368 26568 18420
rect 29092 18411 29144 18420
rect 29092 18377 29101 18411
rect 29101 18377 29135 18411
rect 29135 18377 29144 18411
rect 29092 18368 29144 18377
rect 11796 18300 11848 18352
rect 11980 18300 12032 18352
rect 14188 18300 14240 18352
rect 14832 18300 14884 18352
rect 18880 18300 18932 18352
rect 20168 18300 20220 18352
rect 20720 18300 20772 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 16396 18232 16448 18284
rect 19432 18232 19484 18284
rect 24860 18300 24912 18352
rect 27068 18300 27120 18352
rect 27344 18343 27396 18352
rect 27344 18309 27353 18343
rect 27353 18309 27387 18343
rect 27387 18309 27396 18343
rect 27344 18300 27396 18309
rect 29184 18300 29236 18352
rect 30196 18368 30248 18420
rect 30656 18368 30708 18420
rect 32220 18368 32272 18420
rect 34336 18411 34388 18420
rect 34336 18377 34345 18411
rect 34345 18377 34379 18411
rect 34379 18377 34388 18411
rect 34336 18368 34388 18377
rect 34796 18368 34848 18420
rect 35624 18411 35676 18420
rect 35624 18377 35633 18411
rect 35633 18377 35667 18411
rect 35667 18377 35676 18411
rect 35624 18368 35676 18377
rect 36268 18411 36320 18420
rect 36268 18377 36277 18411
rect 36277 18377 36311 18411
rect 36311 18377 36320 18411
rect 36268 18368 36320 18377
rect 37556 18368 37608 18420
rect 30472 18300 30524 18352
rect 31944 18300 31996 18352
rect 26976 18232 27028 18284
rect 28356 18275 28408 18284
rect 28356 18241 28365 18275
rect 28365 18241 28399 18275
rect 28399 18241 28408 18275
rect 28356 18232 28408 18241
rect 29000 18275 29052 18284
rect 29000 18241 29009 18275
rect 29009 18241 29043 18275
rect 29043 18241 29052 18275
rect 29000 18232 29052 18241
rect 31392 18232 31444 18284
rect 31852 18232 31904 18284
rect 32956 18275 33008 18284
rect 32956 18241 32965 18275
rect 32965 18241 32999 18275
rect 32999 18241 33008 18275
rect 32956 18232 33008 18241
rect 33876 18232 33928 18284
rect 36636 18300 36688 18352
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 16304 18164 16356 18216
rect 23572 18164 23624 18216
rect 27068 18164 27120 18216
rect 19432 18028 19484 18080
rect 20444 18028 20496 18080
rect 25136 18028 25188 18080
rect 27528 18207 27580 18216
rect 27528 18173 27537 18207
rect 27537 18173 27571 18207
rect 27571 18173 27580 18207
rect 27528 18164 27580 18173
rect 29736 18164 29788 18216
rect 31116 18164 31168 18216
rect 35716 18232 35768 18284
rect 37648 18275 37700 18284
rect 37648 18241 37657 18275
rect 37657 18241 37691 18275
rect 37691 18241 37700 18275
rect 37648 18232 37700 18241
rect 33876 18096 33928 18148
rect 31852 18028 31904 18080
rect 33232 18028 33284 18080
rect 36360 18164 36412 18216
rect 37464 18164 37516 18216
rect 38016 18164 38068 18216
rect 34244 18096 34296 18148
rect 37464 18028 37516 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4068 17867 4120 17876
rect 4068 17833 4077 17867
rect 4077 17833 4111 17867
rect 4111 17833 4120 17867
rect 4068 17824 4120 17833
rect 11060 17824 11112 17876
rect 17960 17824 18012 17876
rect 1860 17756 1912 17808
rect 14280 17756 14332 17808
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 10600 17688 10652 17740
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 12256 17688 12308 17740
rect 13544 17688 13596 17740
rect 27068 17824 27120 17876
rect 1952 17620 2004 17672
rect 9128 17620 9180 17672
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 17684 17663 17736 17672
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 19984 17688 20036 17740
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 22836 17688 22888 17740
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 25044 17688 25096 17740
rect 29644 17756 29696 17808
rect 30012 17824 30064 17876
rect 30196 17824 30248 17876
rect 37372 17824 37424 17876
rect 37740 17824 37792 17876
rect 27160 17688 27212 17740
rect 29092 17688 29144 17740
rect 22468 17620 22520 17672
rect 26608 17620 26660 17672
rect 28080 17663 28132 17672
rect 28080 17629 28089 17663
rect 28089 17629 28123 17663
rect 28123 17629 28132 17663
rect 28540 17663 28592 17672
rect 28080 17620 28132 17629
rect 28540 17629 28549 17663
rect 28549 17629 28583 17663
rect 28583 17629 28592 17663
rect 28540 17620 28592 17629
rect 29184 17620 29236 17672
rect 29460 17620 29512 17672
rect 30380 17756 30432 17808
rect 31944 17731 31996 17740
rect 31944 17697 31953 17731
rect 31953 17697 31987 17731
rect 31987 17697 31996 17731
rect 31944 17688 31996 17697
rect 32128 17688 32180 17740
rect 33968 17731 34020 17740
rect 33968 17697 33977 17731
rect 33977 17697 34011 17731
rect 34011 17697 34020 17731
rect 33968 17688 34020 17697
rect 34520 17688 34572 17740
rect 34704 17688 34756 17740
rect 37648 17756 37700 17808
rect 35716 17688 35768 17740
rect 37188 17688 37240 17740
rect 30380 17663 30432 17672
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 30380 17620 30432 17629
rect 35348 17620 35400 17672
rect 36176 17663 36228 17672
rect 9956 17595 10008 17604
rect 9956 17561 9965 17595
rect 9965 17561 9999 17595
rect 9999 17561 10008 17595
rect 9956 17552 10008 17561
rect 10968 17552 11020 17604
rect 12164 17595 12216 17604
rect 12164 17561 12173 17595
rect 12173 17561 12207 17595
rect 12207 17561 12216 17595
rect 12164 17552 12216 17561
rect 13452 17552 13504 17604
rect 16488 17552 16540 17604
rect 17960 17484 18012 17536
rect 20720 17552 20772 17604
rect 21364 17552 21416 17604
rect 21640 17552 21692 17604
rect 22744 17595 22796 17604
rect 22744 17561 22753 17595
rect 22753 17561 22787 17595
rect 22787 17561 22796 17595
rect 22744 17552 22796 17561
rect 26976 17552 27028 17604
rect 28632 17595 28684 17604
rect 28632 17561 28641 17595
rect 28641 17561 28675 17595
rect 28675 17561 28684 17595
rect 28632 17552 28684 17561
rect 22560 17484 22612 17536
rect 25320 17484 25372 17536
rect 33232 17595 33284 17604
rect 33232 17561 33241 17595
rect 33241 17561 33275 17595
rect 33275 17561 33284 17595
rect 33232 17552 33284 17561
rect 33784 17552 33836 17604
rect 34336 17552 34388 17604
rect 36176 17629 36185 17663
rect 36185 17629 36219 17663
rect 36219 17629 36228 17663
rect 36176 17620 36228 17629
rect 37280 17620 37332 17672
rect 37464 17663 37516 17672
rect 37464 17629 37473 17663
rect 37473 17629 37507 17663
rect 37507 17629 37516 17663
rect 37464 17620 37516 17629
rect 37832 17552 37884 17604
rect 35992 17484 36044 17536
rect 36268 17527 36320 17536
rect 36268 17493 36277 17527
rect 36277 17493 36311 17527
rect 36311 17493 36320 17527
rect 36268 17484 36320 17493
rect 36452 17484 36504 17536
rect 36636 17484 36688 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 11244 17280 11296 17332
rect 14188 17280 14240 17332
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 21364 17323 21416 17332
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 25044 17280 25096 17332
rect 27068 17280 27120 17332
rect 27252 17323 27304 17332
rect 27252 17289 27261 17323
rect 27261 17289 27295 17323
rect 27295 17289 27304 17323
rect 27252 17280 27304 17289
rect 9956 17212 10008 17264
rect 17684 17212 17736 17264
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 12532 17144 12584 17196
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 17960 17144 18012 17196
rect 18236 17144 18288 17196
rect 20812 17144 20864 17196
rect 20996 17144 21048 17196
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 22468 17212 22520 17264
rect 28448 17280 28500 17332
rect 29184 17212 29236 17264
rect 29460 17255 29512 17264
rect 29460 17221 29469 17255
rect 29469 17221 29503 17255
rect 29503 17221 29512 17255
rect 29460 17212 29512 17221
rect 29644 17212 29696 17264
rect 33968 17280 34020 17332
rect 25228 17144 25280 17196
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 27436 17144 27488 17196
rect 30288 17144 30340 17196
rect 17776 17076 17828 17128
rect 12992 16940 13044 16992
rect 20168 17008 20220 17060
rect 21640 17008 21692 17060
rect 27988 17076 28040 17128
rect 28448 17119 28500 17128
rect 27252 17008 27304 17060
rect 25412 16940 25464 16992
rect 25596 16940 25648 16992
rect 28448 17085 28457 17119
rect 28457 17085 28491 17119
rect 28491 17085 28500 17119
rect 28448 17076 28500 17085
rect 28540 17076 28592 17128
rect 31852 17076 31904 17128
rect 30748 17008 30800 17060
rect 30932 17008 30984 17060
rect 31944 17008 31996 17060
rect 34152 17212 34204 17264
rect 34796 17212 34848 17264
rect 35348 17212 35400 17264
rect 37372 17212 37424 17264
rect 38476 17212 38528 17264
rect 38844 17212 38896 17264
rect 34152 17119 34204 17128
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 35716 17119 35768 17128
rect 33968 17008 34020 17060
rect 35716 17085 35725 17119
rect 35725 17085 35759 17119
rect 35759 17085 35768 17119
rect 35716 17076 35768 17085
rect 35900 17076 35952 17128
rect 37556 17119 37608 17128
rect 37556 17085 37565 17119
rect 37565 17085 37599 17119
rect 37599 17085 37608 17119
rect 37556 17076 37608 17085
rect 38292 17076 38344 17128
rect 36268 16940 36320 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 12808 16736 12860 16788
rect 17040 16736 17092 16788
rect 17592 16736 17644 16788
rect 22744 16736 22796 16788
rect 26976 16736 27028 16788
rect 29184 16736 29236 16788
rect 13268 16668 13320 16720
rect 1584 16600 1636 16652
rect 16856 16600 16908 16652
rect 17040 16600 17092 16652
rect 18972 16668 19024 16720
rect 20812 16711 20864 16720
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 14004 16532 14056 16584
rect 14924 16532 14976 16584
rect 19064 16600 19116 16652
rect 20812 16677 20821 16711
rect 20821 16677 20855 16711
rect 20855 16677 20864 16711
rect 20812 16668 20864 16677
rect 19984 16600 20036 16652
rect 26148 16668 26200 16720
rect 35532 16736 35584 16788
rect 25504 16643 25556 16652
rect 25504 16609 25513 16643
rect 25513 16609 25547 16643
rect 25547 16609 25556 16643
rect 25504 16600 25556 16609
rect 26792 16600 26844 16652
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 21548 16532 21600 16541
rect 22560 16532 22612 16584
rect 27160 16600 27212 16652
rect 30380 16668 30432 16720
rect 35164 16668 35216 16720
rect 35900 16668 35952 16720
rect 30104 16600 30156 16652
rect 30472 16575 30524 16584
rect 30472 16541 30481 16575
rect 30481 16541 30515 16575
rect 30515 16541 30524 16575
rect 31024 16575 31076 16584
rect 30472 16532 30524 16541
rect 31024 16541 31033 16575
rect 31033 16541 31067 16575
rect 31067 16541 31076 16575
rect 31024 16532 31076 16541
rect 31116 16575 31168 16584
rect 31116 16541 31125 16575
rect 31125 16541 31159 16575
rect 31159 16541 31168 16575
rect 31760 16600 31812 16652
rect 32680 16600 32732 16652
rect 33048 16600 33100 16652
rect 31116 16532 31168 16541
rect 32404 16532 32456 16584
rect 32772 16532 32824 16584
rect 33508 16532 33560 16584
rect 36268 16600 36320 16652
rect 37464 16600 37516 16652
rect 10048 16464 10100 16516
rect 16764 16464 16816 16516
rect 16948 16464 17000 16516
rect 20536 16464 20588 16516
rect 20720 16464 20772 16516
rect 10784 16396 10836 16448
rect 17040 16396 17092 16448
rect 19432 16396 19484 16448
rect 20076 16396 20128 16448
rect 22284 16396 22336 16448
rect 25596 16507 25648 16516
rect 25596 16473 25605 16507
rect 25605 16473 25639 16507
rect 25639 16473 25648 16507
rect 26516 16507 26568 16516
rect 25596 16464 25648 16473
rect 26516 16473 26525 16507
rect 26525 16473 26559 16507
rect 26559 16473 26568 16507
rect 28080 16507 28132 16516
rect 26516 16464 26568 16473
rect 27620 16396 27672 16448
rect 28080 16473 28089 16507
rect 28089 16473 28123 16507
rect 28123 16473 28132 16507
rect 28080 16464 28132 16473
rect 28172 16507 28224 16516
rect 28172 16473 28181 16507
rect 28181 16473 28215 16507
rect 28215 16473 28224 16507
rect 28172 16464 28224 16473
rect 29276 16464 29328 16516
rect 30196 16464 30248 16516
rect 31300 16464 31352 16516
rect 35900 16507 35952 16516
rect 35900 16473 35909 16507
rect 35909 16473 35943 16507
rect 35943 16473 35952 16507
rect 35900 16464 35952 16473
rect 37924 16464 37976 16516
rect 29920 16396 29972 16448
rect 31760 16439 31812 16448
rect 31760 16405 31769 16439
rect 31769 16405 31803 16439
rect 31803 16405 31812 16439
rect 31760 16396 31812 16405
rect 32496 16396 32548 16448
rect 33692 16439 33744 16448
rect 33692 16405 33701 16439
rect 33701 16405 33735 16439
rect 33735 16405 33744 16439
rect 33692 16396 33744 16405
rect 34980 16439 35032 16448
rect 34980 16405 34989 16439
rect 34989 16405 35023 16439
rect 35023 16405 35032 16439
rect 34980 16396 35032 16405
rect 39488 16396 39540 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11980 16192 12032 16244
rect 12716 16124 12768 16176
rect 14004 16124 14056 16176
rect 10784 16056 10836 16108
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 8484 15920 8536 15972
rect 11428 15988 11480 16040
rect 14372 16167 14424 16176
rect 14372 16133 14381 16167
rect 14381 16133 14415 16167
rect 14415 16133 14424 16167
rect 14372 16124 14424 16133
rect 14740 16192 14792 16244
rect 16304 16124 16356 16176
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 19984 16192 20036 16244
rect 22652 16124 22704 16176
rect 28172 16192 28224 16244
rect 29460 16192 29512 16244
rect 31484 16192 31536 16244
rect 33692 16192 33744 16244
rect 35256 16192 35308 16244
rect 36452 16235 36504 16244
rect 36452 16201 36461 16235
rect 36461 16201 36495 16235
rect 36495 16201 36504 16235
rect 36452 16192 36504 16201
rect 16948 16031 17000 16040
rect 13728 15920 13780 15972
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 19800 16056 19852 16108
rect 20352 16056 20404 16108
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 28724 16056 28776 16108
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 30196 16099 30248 16108
rect 30196 16065 30205 16099
rect 30205 16065 30239 16099
rect 30239 16065 30248 16099
rect 30196 16056 30248 16065
rect 32220 16124 32272 16176
rect 32404 16124 32456 16176
rect 33784 16124 33836 16176
rect 37740 16167 37792 16176
rect 37740 16133 37749 16167
rect 37749 16133 37783 16167
rect 37783 16133 37792 16167
rect 37740 16124 37792 16133
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 35532 16056 35584 16108
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 10600 15852 10652 15904
rect 20536 15988 20588 16040
rect 22652 16031 22704 16040
rect 22652 15997 22662 16031
rect 22662 15997 22696 16031
rect 22696 15997 22704 16031
rect 22652 15988 22704 15997
rect 17316 15920 17368 15972
rect 31668 15988 31720 16040
rect 32036 15988 32088 16040
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 33324 16031 33376 16040
rect 33324 15997 33333 16031
rect 33333 15997 33367 16031
rect 33367 15997 33376 16031
rect 33324 15988 33376 15997
rect 33692 15988 33744 16040
rect 34152 15988 34204 16040
rect 34520 15920 34572 15972
rect 35440 15988 35492 16040
rect 35164 15920 35216 15972
rect 36452 16056 36504 16108
rect 37648 16031 37700 16040
rect 37648 15997 37657 16031
rect 37657 15997 37691 16031
rect 37691 15997 37700 16031
rect 37648 15988 37700 15997
rect 38292 16031 38344 16040
rect 38292 15997 38301 16031
rect 38301 15997 38335 16031
rect 38335 15997 38344 16031
rect 38292 15988 38344 15997
rect 36176 15920 36228 15972
rect 36728 15920 36780 15972
rect 17592 15852 17644 15904
rect 19984 15852 20036 15904
rect 20628 15852 20680 15904
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 26332 15852 26384 15904
rect 29184 15852 29236 15904
rect 32036 15852 32088 15904
rect 32588 15852 32640 15904
rect 38200 15852 38252 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 14464 15648 14516 15700
rect 19800 15691 19852 15700
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 12256 15580 12308 15632
rect 17316 15580 17368 15632
rect 19800 15657 19809 15691
rect 19809 15657 19843 15691
rect 19843 15657 19852 15691
rect 19800 15648 19852 15657
rect 24952 15648 25004 15700
rect 32588 15648 32640 15700
rect 19984 15580 20036 15632
rect 26516 15580 26568 15632
rect 27252 15580 27304 15632
rect 28540 15580 28592 15632
rect 30932 15623 30984 15632
rect 30932 15589 30941 15623
rect 30941 15589 30975 15623
rect 30975 15589 30984 15623
rect 30932 15580 30984 15589
rect 11704 15512 11756 15564
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 14464 15444 14516 15496
rect 18052 15444 18104 15496
rect 19432 15444 19484 15496
rect 21456 15487 21508 15496
rect 17960 15376 18012 15428
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 21548 15444 21600 15496
rect 23388 15376 23440 15428
rect 29276 15444 29328 15496
rect 29368 15444 29420 15496
rect 31576 15512 31628 15564
rect 30748 15444 30800 15496
rect 32220 15580 32272 15632
rect 33232 15623 33284 15632
rect 33232 15589 33241 15623
rect 33241 15589 33275 15623
rect 33275 15589 33284 15623
rect 33232 15580 33284 15589
rect 33784 15648 33836 15700
rect 34796 15648 34848 15700
rect 39028 15648 39080 15700
rect 35716 15580 35768 15632
rect 32864 15512 32916 15564
rect 36360 15512 36412 15564
rect 34888 15487 34940 15496
rect 34888 15453 34897 15487
rect 34897 15453 34931 15487
rect 34931 15453 34940 15487
rect 34888 15444 34940 15453
rect 37464 15444 37516 15496
rect 38016 15487 38068 15496
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 28724 15419 28776 15428
rect 28724 15385 28733 15419
rect 28733 15385 28767 15419
rect 28767 15385 28776 15419
rect 28724 15376 28776 15385
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 13268 15308 13320 15360
rect 18236 15351 18288 15360
rect 18236 15317 18245 15351
rect 18245 15317 18279 15351
rect 18279 15317 18288 15351
rect 18236 15308 18288 15317
rect 21180 15308 21232 15360
rect 25044 15351 25096 15360
rect 25044 15317 25053 15351
rect 25053 15317 25087 15351
rect 25087 15317 25096 15351
rect 25044 15308 25096 15317
rect 27344 15308 27396 15360
rect 27620 15308 27672 15360
rect 31944 15376 31996 15428
rect 31392 15308 31444 15360
rect 31760 15308 31812 15360
rect 34612 15376 34664 15428
rect 37924 15376 37976 15428
rect 32956 15308 33008 15360
rect 35440 15308 35492 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 11428 15104 11480 15156
rect 11520 15104 11572 15156
rect 10876 15036 10928 15088
rect 17776 15104 17828 15156
rect 18880 15104 18932 15156
rect 19432 15104 19484 15156
rect 19984 15104 20036 15156
rect 13268 15079 13320 15088
rect 13268 15045 13277 15079
rect 13277 15045 13311 15079
rect 13311 15045 13320 15079
rect 13268 15036 13320 15045
rect 1676 14968 1728 15020
rect 11888 15011 11940 15020
rect 8760 14900 8812 14952
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 20168 15036 20220 15088
rect 20260 15036 20312 15088
rect 20628 15036 20680 15088
rect 18052 14968 18104 15020
rect 20076 14968 20128 15020
rect 20812 14968 20864 15020
rect 24216 15104 24268 15156
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 28356 15104 28408 15156
rect 33048 15104 33100 15156
rect 36176 15104 36228 15156
rect 36544 15104 36596 15156
rect 38108 15104 38160 15156
rect 27344 15079 27396 15088
rect 27344 15045 27353 15079
rect 27353 15045 27387 15079
rect 27387 15045 27396 15079
rect 27344 15036 27396 15045
rect 29184 15079 29236 15088
rect 29184 15045 29193 15079
rect 29193 15045 29227 15079
rect 29227 15045 29236 15079
rect 29184 15036 29236 15045
rect 32496 15079 32548 15088
rect 32496 15045 32505 15079
rect 32505 15045 32539 15079
rect 32539 15045 32548 15079
rect 32496 15036 32548 15045
rect 31208 14968 31260 15020
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 34428 15036 34480 15088
rect 34520 15036 34572 15088
rect 33232 14968 33284 15020
rect 34244 14968 34296 15020
rect 34888 15011 34940 15020
rect 34888 14977 34897 15011
rect 34897 14977 34931 15011
rect 34931 14977 34940 15011
rect 34888 14968 34940 14977
rect 14372 14900 14424 14952
rect 22836 14943 22888 14952
rect 22836 14909 22845 14943
rect 22845 14909 22879 14943
rect 22879 14909 22888 14943
rect 22836 14900 22888 14909
rect 26884 14900 26936 14952
rect 27252 14943 27304 14952
rect 27252 14909 27261 14943
rect 27261 14909 27295 14943
rect 27295 14909 27304 14943
rect 27252 14900 27304 14909
rect 27620 14943 27672 14952
rect 27620 14909 27629 14943
rect 27629 14909 27663 14943
rect 27663 14909 27672 14943
rect 27620 14900 27672 14909
rect 29736 14943 29788 14952
rect 19248 14832 19300 14884
rect 13452 14764 13504 14816
rect 13636 14764 13688 14816
rect 17132 14764 17184 14816
rect 26976 14832 27028 14884
rect 29736 14909 29745 14943
rect 29745 14909 29779 14943
rect 29779 14909 29788 14943
rect 29736 14900 29788 14909
rect 32220 14900 32272 14952
rect 33324 14900 33376 14952
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 33508 14900 33560 14909
rect 35624 14900 35676 14952
rect 32128 14832 32180 14884
rect 32312 14832 32364 14884
rect 36452 15036 36504 15088
rect 36636 14968 36688 15020
rect 38108 15011 38160 15020
rect 38108 14977 38117 15011
rect 38117 14977 38151 15011
rect 38151 14977 38160 15011
rect 38108 14968 38160 14977
rect 39764 14968 39816 15020
rect 37188 14900 37240 14952
rect 30840 14764 30892 14816
rect 31852 14764 31904 14816
rect 33416 14764 33468 14816
rect 37004 14764 37056 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 27804 14560 27856 14612
rect 31760 14560 31812 14612
rect 32036 14603 32088 14612
rect 32036 14569 32045 14603
rect 32045 14569 32079 14603
rect 32079 14569 32088 14603
rect 32036 14560 32088 14569
rect 32220 14560 32272 14612
rect 36360 14603 36412 14612
rect 36360 14569 36369 14603
rect 36369 14569 36403 14603
rect 36403 14569 36412 14603
rect 36360 14560 36412 14569
rect 39856 14560 39908 14612
rect 25688 14492 25740 14544
rect 11888 14424 11940 14476
rect 15660 14424 15712 14476
rect 16856 14424 16908 14476
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 26976 14467 27028 14476
rect 26976 14433 26985 14467
rect 26985 14433 27019 14467
rect 27019 14433 27028 14467
rect 26976 14424 27028 14433
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 21456 14356 21508 14408
rect 30748 14424 30800 14476
rect 33508 14492 33560 14544
rect 35992 14492 36044 14544
rect 31852 14467 31904 14476
rect 31852 14433 31861 14467
rect 31861 14433 31895 14467
rect 31895 14433 31904 14467
rect 31852 14424 31904 14433
rect 32128 14424 32180 14476
rect 33968 14424 34020 14476
rect 34244 14424 34296 14476
rect 28632 14356 28684 14408
rect 17132 14331 17184 14340
rect 17132 14297 17141 14331
rect 17141 14297 17175 14331
rect 17175 14297 17184 14331
rect 17132 14288 17184 14297
rect 17868 14288 17920 14340
rect 19432 14288 19484 14340
rect 23664 14288 23716 14340
rect 17500 14220 17552 14272
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 22560 14263 22612 14272
rect 22560 14229 22569 14263
rect 22569 14229 22603 14263
rect 22603 14229 22612 14263
rect 22560 14220 22612 14229
rect 25228 14288 25280 14340
rect 27068 14331 27120 14340
rect 27068 14297 27077 14331
rect 27077 14297 27111 14331
rect 27111 14297 27120 14331
rect 27068 14288 27120 14297
rect 27436 14288 27488 14340
rect 30564 14356 30616 14408
rect 32312 14356 32364 14408
rect 35624 14356 35676 14408
rect 35716 14356 35768 14408
rect 39304 14424 39356 14476
rect 38108 14356 38160 14408
rect 29460 14288 29512 14340
rect 33324 14331 33376 14340
rect 25504 14220 25556 14272
rect 29000 14220 29052 14272
rect 30380 14220 30432 14272
rect 33324 14297 33333 14331
rect 33333 14297 33367 14331
rect 33367 14297 33376 14331
rect 33324 14288 33376 14297
rect 33416 14331 33468 14340
rect 33416 14297 33425 14331
rect 33425 14297 33459 14331
rect 33459 14297 33468 14331
rect 33416 14288 33468 14297
rect 34152 14220 34204 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 8484 14016 8536 14068
rect 19248 14059 19300 14068
rect 19248 14025 19257 14059
rect 19257 14025 19291 14059
rect 19291 14025 19300 14059
rect 19248 14016 19300 14025
rect 20628 14016 20680 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 10876 13880 10928 13932
rect 8300 13812 8352 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 14464 13880 14516 13932
rect 16948 13948 17000 14000
rect 17132 13991 17184 14000
rect 17132 13957 17141 13991
rect 17141 13957 17175 13991
rect 17175 13957 17184 13991
rect 17132 13948 17184 13957
rect 18236 13948 18288 14000
rect 20720 13948 20772 14000
rect 21548 13880 21600 13932
rect 25228 14016 25280 14068
rect 22560 13948 22612 14000
rect 23480 13991 23532 14000
rect 23480 13957 23489 13991
rect 23489 13957 23523 13991
rect 23523 13957 23532 13991
rect 23480 13948 23532 13957
rect 25320 13948 25372 14000
rect 25688 13991 25740 14000
rect 25688 13957 25697 13991
rect 25697 13957 25731 13991
rect 25731 13957 25740 13991
rect 25688 13948 25740 13957
rect 26332 13948 26384 14000
rect 28908 13948 28960 14000
rect 28540 13923 28592 13932
rect 17592 13812 17644 13864
rect 17776 13812 17828 13864
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19432 13812 19484 13864
rect 20720 13812 20772 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 26148 13855 26200 13864
rect 26148 13821 26157 13855
rect 26157 13821 26191 13855
rect 26191 13821 26200 13855
rect 26148 13812 26200 13821
rect 28540 13889 28549 13923
rect 28549 13889 28583 13923
rect 28583 13889 28592 13923
rect 28540 13880 28592 13889
rect 29000 13880 29052 13932
rect 32772 14016 32824 14068
rect 34336 14016 34388 14068
rect 38568 14016 38620 14068
rect 30840 13991 30892 14000
rect 30840 13957 30849 13991
rect 30849 13957 30883 13991
rect 30883 13957 30892 13991
rect 30840 13948 30892 13957
rect 33968 13991 34020 14000
rect 33968 13957 33977 13991
rect 33977 13957 34011 13991
rect 34011 13957 34020 13991
rect 33968 13948 34020 13957
rect 35532 13991 35584 14000
rect 35532 13957 35541 13991
rect 35541 13957 35575 13991
rect 35575 13957 35584 13991
rect 35532 13948 35584 13957
rect 36452 13991 36504 14000
rect 36452 13957 36461 13991
rect 36461 13957 36495 13991
rect 36495 13957 36504 13991
rect 36452 13948 36504 13957
rect 38660 13948 38712 14000
rect 33232 13880 33284 13932
rect 36636 13880 36688 13932
rect 38108 13923 38160 13932
rect 38108 13889 38117 13923
rect 38117 13889 38151 13923
rect 38151 13889 38160 13923
rect 38108 13880 38160 13889
rect 27344 13855 27396 13864
rect 27344 13821 27353 13855
rect 27353 13821 27387 13855
rect 27387 13821 27396 13855
rect 27344 13812 27396 13821
rect 31668 13855 31720 13864
rect 31668 13821 31677 13855
rect 31677 13821 31711 13855
rect 31711 13821 31720 13855
rect 31668 13812 31720 13821
rect 31852 13812 31904 13864
rect 34152 13855 34204 13864
rect 34152 13821 34161 13855
rect 34161 13821 34195 13855
rect 34195 13821 34204 13855
rect 34152 13812 34204 13821
rect 35440 13855 35492 13864
rect 35440 13821 35449 13855
rect 35449 13821 35483 13855
rect 35483 13821 35492 13855
rect 35440 13812 35492 13821
rect 33508 13744 33560 13796
rect 33692 13744 33744 13796
rect 19616 13676 19668 13728
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 13176 13472 13228 13524
rect 18328 13472 18380 13524
rect 18604 13472 18656 13524
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20996 13472 21048 13524
rect 27344 13472 27396 13524
rect 32864 13515 32916 13524
rect 32864 13481 32873 13515
rect 32873 13481 32907 13515
rect 32907 13481 32916 13515
rect 32864 13472 32916 13481
rect 33968 13472 34020 13524
rect 35532 13472 35584 13524
rect 36360 13472 36412 13524
rect 39212 13472 39264 13524
rect 13636 13404 13688 13456
rect 13820 13404 13872 13456
rect 24860 13404 24912 13456
rect 26148 13404 26200 13456
rect 27068 13404 27120 13456
rect 33140 13404 33192 13456
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 15660 13336 15712 13388
rect 20168 13336 20220 13388
rect 20904 13336 20956 13388
rect 15016 13268 15068 13320
rect 17868 13268 17920 13320
rect 19616 13311 19668 13320
rect 19616 13277 19625 13311
rect 19625 13277 19659 13311
rect 19659 13277 19668 13311
rect 19616 13268 19668 13277
rect 23480 13268 23532 13320
rect 24032 13268 24084 13320
rect 26056 13268 26108 13320
rect 26424 13268 26476 13320
rect 32956 13336 33008 13388
rect 35532 13336 35584 13388
rect 35992 13336 36044 13388
rect 36360 13336 36412 13388
rect 25136 13243 25188 13252
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 27896 13200 27948 13252
rect 33692 13268 33744 13320
rect 35808 13268 35860 13320
rect 12164 13132 12216 13184
rect 22928 13175 22980 13184
rect 22928 13141 22937 13175
rect 22937 13141 22971 13175
rect 22971 13141 22980 13175
rect 22928 13132 22980 13141
rect 24952 13132 25004 13184
rect 26884 13132 26936 13184
rect 32864 13200 32916 13252
rect 37188 13311 37240 13320
rect 37188 13277 37197 13311
rect 37197 13277 37231 13311
rect 37231 13277 37240 13311
rect 37188 13268 37240 13277
rect 37832 13268 37884 13320
rect 34796 13132 34848 13184
rect 34888 13132 34940 13184
rect 38016 13132 38068 13184
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 10508 12928 10560 12980
rect 13176 12928 13228 12980
rect 15016 12971 15068 12980
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 19156 12928 19208 12980
rect 26424 12971 26476 12980
rect 26424 12937 26433 12971
rect 26433 12937 26467 12971
rect 26467 12937 26476 12971
rect 26424 12928 26476 12937
rect 29368 12971 29420 12980
rect 29368 12937 29377 12971
rect 29377 12937 29411 12971
rect 29411 12937 29420 12971
rect 29368 12928 29420 12937
rect 32312 12971 32364 12980
rect 32312 12937 32321 12971
rect 32321 12937 32355 12971
rect 32355 12937 32364 12971
rect 32312 12928 32364 12937
rect 34888 12928 34940 12980
rect 35348 12928 35400 12980
rect 35900 12928 35952 12980
rect 36268 12971 36320 12980
rect 36268 12937 36277 12971
rect 36277 12937 36311 12971
rect 36311 12937 36320 12971
rect 36268 12928 36320 12937
rect 37280 12928 37332 12980
rect 37924 12928 37976 12980
rect 11612 12860 11664 12912
rect 18328 12903 18380 12912
rect 8300 12792 8352 12844
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 18328 12869 18337 12903
rect 18337 12869 18371 12903
rect 18371 12869 18380 12903
rect 18328 12860 18380 12869
rect 20076 12860 20128 12912
rect 20168 12792 20220 12844
rect 23480 12792 23532 12844
rect 27436 12792 27488 12844
rect 29276 12835 29328 12844
rect 29276 12801 29285 12835
rect 29285 12801 29319 12835
rect 29319 12801 29328 12835
rect 29276 12792 29328 12801
rect 33784 12860 33836 12912
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 33140 12835 33192 12844
rect 33140 12801 33149 12835
rect 33149 12801 33183 12835
rect 33183 12801 33192 12835
rect 33140 12792 33192 12801
rect 34520 12860 34572 12912
rect 34704 12860 34756 12912
rect 34152 12792 34204 12844
rect 12440 12724 12492 12776
rect 16212 12724 16264 12776
rect 28816 12724 28868 12776
rect 34980 12792 35032 12844
rect 36820 12724 36872 12776
rect 33508 12656 33560 12708
rect 33692 12699 33744 12708
rect 33692 12665 33701 12699
rect 33701 12665 33735 12699
rect 33735 12665 33744 12699
rect 33692 12656 33744 12665
rect 37280 12724 37332 12776
rect 37924 12767 37976 12776
rect 37924 12733 37933 12767
rect 37933 12733 37967 12767
rect 37967 12733 37976 12767
rect 37924 12724 37976 12733
rect 38108 12656 38160 12708
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 23020 12588 23072 12640
rect 33140 12588 33192 12640
rect 34796 12588 34848 12640
rect 36544 12588 36596 12640
rect 36728 12588 36780 12640
rect 37464 12588 37516 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 20076 12427 20128 12436
rect 20076 12393 20085 12427
rect 20085 12393 20119 12427
rect 20119 12393 20128 12427
rect 20076 12384 20128 12393
rect 24952 12316 25004 12368
rect 17592 12291 17644 12300
rect 4620 12180 4672 12232
rect 11612 12180 11664 12232
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 22560 12248 22612 12300
rect 22928 12248 22980 12300
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 16948 12155 17000 12164
rect 16948 12121 16957 12155
rect 16957 12121 16991 12155
rect 16991 12121 17000 12155
rect 16948 12112 17000 12121
rect 17040 12155 17092 12164
rect 17040 12121 17049 12155
rect 17049 12121 17083 12155
rect 17083 12121 17092 12155
rect 17040 12112 17092 12121
rect 22836 12044 22888 12096
rect 23112 12044 23164 12096
rect 32864 12384 32916 12436
rect 33416 12427 33468 12436
rect 33416 12393 33425 12427
rect 33425 12393 33459 12427
rect 33459 12393 33468 12427
rect 33416 12384 33468 12393
rect 34244 12427 34296 12436
rect 34244 12393 34253 12427
rect 34253 12393 34287 12427
rect 34287 12393 34296 12427
rect 34244 12384 34296 12393
rect 35716 12384 35768 12436
rect 37096 12384 37148 12436
rect 39120 12384 39172 12436
rect 38384 12316 38436 12368
rect 38844 12316 38896 12368
rect 37556 12291 37608 12300
rect 37556 12257 37565 12291
rect 37565 12257 37599 12291
rect 37599 12257 37608 12291
rect 37556 12248 37608 12257
rect 29828 12180 29880 12232
rect 32312 12180 32364 12232
rect 33600 12180 33652 12232
rect 34428 12180 34480 12232
rect 36084 12223 36136 12232
rect 26884 12155 26936 12164
rect 26884 12121 26893 12155
rect 26893 12121 26927 12155
rect 26927 12121 26936 12155
rect 26884 12112 26936 12121
rect 36084 12189 36093 12223
rect 36093 12189 36127 12223
rect 36127 12189 36136 12223
rect 36084 12180 36136 12189
rect 36544 12223 36596 12232
rect 36544 12189 36553 12223
rect 36553 12189 36587 12223
rect 36587 12189 36596 12223
rect 36544 12180 36596 12189
rect 37096 12112 37148 12164
rect 38752 12044 38804 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 10416 11840 10468 11892
rect 16672 11840 16724 11892
rect 16764 11840 16816 11892
rect 17040 11840 17092 11892
rect 20996 11840 21048 11892
rect 23940 11883 23992 11892
rect 23940 11849 23949 11883
rect 23949 11849 23983 11883
rect 23983 11849 23992 11883
rect 23940 11840 23992 11849
rect 34612 11840 34664 11892
rect 35440 11883 35492 11892
rect 35440 11849 35449 11883
rect 35449 11849 35483 11883
rect 35483 11849 35492 11883
rect 35440 11840 35492 11849
rect 37188 11840 37240 11892
rect 37556 11883 37608 11892
rect 37556 11849 37565 11883
rect 37565 11849 37599 11883
rect 37599 11849 37608 11883
rect 37556 11840 37608 11849
rect 36268 11815 36320 11824
rect 7564 11704 7616 11756
rect 14188 11704 14240 11756
rect 16672 11704 16724 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 15660 11636 15712 11688
rect 17592 11636 17644 11688
rect 16396 11568 16448 11620
rect 20628 11704 20680 11756
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26240 11704 26292 11713
rect 26700 11704 26752 11756
rect 36268 11781 36277 11815
rect 36277 11781 36311 11815
rect 36311 11781 36320 11815
rect 36268 11772 36320 11781
rect 36360 11815 36412 11824
rect 36360 11781 36369 11815
rect 36369 11781 36403 11815
rect 36403 11781 36412 11815
rect 36360 11772 36412 11781
rect 36544 11772 36596 11824
rect 34060 11704 34112 11756
rect 37556 11704 37608 11756
rect 38200 11704 38252 11756
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 20904 11636 20956 11688
rect 22744 11679 22796 11688
rect 22744 11645 22753 11679
rect 22753 11645 22787 11679
rect 22787 11645 22796 11679
rect 22744 11636 22796 11645
rect 22836 11636 22888 11688
rect 25136 11679 25188 11688
rect 25136 11645 25145 11679
rect 25145 11645 25179 11679
rect 25179 11645 25188 11679
rect 25136 11636 25188 11645
rect 25320 11636 25372 11688
rect 19616 11568 19668 11620
rect 17592 11543 17644 11552
rect 17592 11509 17601 11543
rect 17601 11509 17635 11543
rect 17635 11509 17644 11543
rect 17592 11500 17644 11509
rect 23112 11543 23164 11552
rect 23112 11509 23121 11543
rect 23121 11509 23155 11543
rect 23155 11509 23164 11543
rect 23112 11500 23164 11509
rect 34336 11500 34388 11552
rect 35624 11568 35676 11620
rect 37556 11568 37608 11620
rect 36728 11500 36780 11552
rect 36912 11500 36964 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 17132 11296 17184 11348
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 34704 11296 34756 11348
rect 36268 11296 36320 11348
rect 9496 11228 9548 11280
rect 36084 11228 36136 11280
rect 16948 11160 17000 11212
rect 17592 11160 17644 11212
rect 20812 11160 20864 11212
rect 28816 11160 28868 11212
rect 31668 11160 31720 11212
rect 33876 11160 33928 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 7656 11092 7708 11144
rect 16396 11135 16448 11144
rect 16396 11101 16405 11135
rect 16405 11101 16439 11135
rect 16439 11101 16448 11135
rect 16396 11092 16448 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 21548 11092 21600 11144
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 17040 11024 17092 11076
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 19616 11024 19668 11033
rect 24952 11024 25004 11076
rect 25412 11024 25464 11076
rect 31852 11092 31904 11144
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 34336 11135 34388 11144
rect 34336 11101 34345 11135
rect 34345 11101 34379 11135
rect 34379 11101 34388 11135
rect 34336 11092 34388 11101
rect 34428 11092 34480 11144
rect 37648 11160 37700 11212
rect 36544 11092 36596 11144
rect 32496 11024 32548 11076
rect 37740 11024 37792 11076
rect 20996 10956 21048 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 8760 10752 8812 10804
rect 20904 10752 20956 10804
rect 32404 10752 32456 10804
rect 35992 10752 36044 10804
rect 37372 10752 37424 10804
rect 13728 10684 13780 10736
rect 17040 10727 17092 10736
rect 17040 10693 17049 10727
rect 17049 10693 17083 10727
rect 17083 10693 17092 10727
rect 17040 10684 17092 10693
rect 25320 10684 25372 10736
rect 36360 10684 36412 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 26240 10616 26292 10668
rect 28908 10616 28960 10668
rect 34428 10659 34480 10668
rect 10968 10548 11020 10600
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 13728 10548 13780 10600
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 24676 10548 24728 10600
rect 27804 10548 27856 10600
rect 34428 10625 34437 10659
rect 34437 10625 34471 10659
rect 34471 10625 34480 10659
rect 34428 10616 34480 10625
rect 36084 10659 36136 10668
rect 36084 10625 36093 10659
rect 36093 10625 36127 10659
rect 36127 10625 36136 10659
rect 36084 10616 36136 10625
rect 38476 10684 38528 10736
rect 37464 10616 37516 10668
rect 38384 10548 38436 10600
rect 37740 10480 37792 10532
rect 24768 10412 24820 10464
rect 29000 10412 29052 10464
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10140 10208 10192 10260
rect 25872 10251 25924 10260
rect 25872 10217 25881 10251
rect 25881 10217 25915 10251
rect 25915 10217 25924 10251
rect 25872 10208 25924 10217
rect 36728 10251 36780 10260
rect 36728 10217 36737 10251
rect 36737 10217 36771 10251
rect 36771 10217 36780 10251
rect 36728 10208 36780 10217
rect 7196 10004 7248 10056
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 24860 10140 24912 10192
rect 35532 10140 35584 10192
rect 23112 10072 23164 10124
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 24952 10115 25004 10124
rect 24952 10081 24961 10115
rect 24961 10081 24995 10115
rect 24995 10081 25004 10115
rect 24952 10072 25004 10081
rect 22100 10004 22152 10056
rect 36176 10047 36228 10056
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 16948 9868 17000 9920
rect 19432 9868 19484 9920
rect 20812 9868 20864 9920
rect 22376 9911 22428 9920
rect 22376 9877 22385 9911
rect 22385 9877 22419 9911
rect 22419 9877 22428 9911
rect 22376 9868 22428 9877
rect 24584 9868 24636 9920
rect 36176 10013 36185 10047
rect 36185 10013 36219 10047
rect 36219 10013 36228 10047
rect 36176 10004 36228 10013
rect 36636 10047 36688 10056
rect 36636 10013 36645 10047
rect 36645 10013 36679 10047
rect 36679 10013 36688 10047
rect 36636 10004 36688 10013
rect 37556 10004 37608 10056
rect 35992 9911 36044 9920
rect 35992 9877 36001 9911
rect 36001 9877 36035 9911
rect 36035 9877 36044 9911
rect 35992 9868 36044 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 8852 9596 8904 9648
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 9312 9596 9364 9648
rect 13360 9596 13412 9648
rect 19340 9596 19392 9648
rect 22100 9639 22152 9648
rect 5816 9460 5868 9512
rect 17040 9528 17092 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 22100 9605 22109 9639
rect 22109 9605 22143 9639
rect 22143 9605 22152 9639
rect 22100 9596 22152 9605
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 30380 9639 30432 9648
rect 30380 9605 30389 9639
rect 30389 9605 30423 9639
rect 30423 9605 30432 9639
rect 30380 9596 30432 9605
rect 36452 9596 36504 9648
rect 37280 9596 37332 9648
rect 23480 9528 23532 9580
rect 27160 9528 27212 9580
rect 37740 9528 37792 9580
rect 39672 9528 39724 9580
rect 20444 9460 20496 9512
rect 22744 9392 22796 9444
rect 37832 9435 37884 9444
rect 37832 9401 37841 9435
rect 37841 9401 37875 9435
rect 37875 9401 37884 9435
rect 37832 9392 37884 9401
rect 7104 9324 7156 9376
rect 19892 9324 19944 9376
rect 22376 9324 22428 9376
rect 28080 9324 28132 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 20444 9163 20496 9172
rect 20444 9129 20453 9163
rect 20453 9129 20487 9163
rect 20487 9129 20496 9163
rect 20444 9120 20496 9129
rect 19340 8984 19392 9036
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 19892 8916 19944 8968
rect 28080 8959 28132 8968
rect 28080 8925 28089 8959
rect 28089 8925 28123 8959
rect 28123 8925 28132 8959
rect 28080 8916 28132 8925
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 30380 8780 30432 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 18052 8576 18104 8628
rect 25136 8576 25188 8628
rect 38108 8619 38160 8628
rect 38108 8585 38117 8619
rect 38117 8585 38151 8619
rect 38151 8585 38160 8619
rect 38108 8576 38160 8585
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 19432 8483 19484 8492
rect 5632 8372 5684 8424
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 38752 8508 38804 8560
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 5724 8304 5776 8356
rect 27252 8304 27304 8356
rect 36636 8304 36688 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 20352 7896 20404 7948
rect 6920 7828 6972 7880
rect 25044 7828 25096 7880
rect 29000 7871 29052 7880
rect 29000 7837 29009 7871
rect 29009 7837 29043 7871
rect 29043 7837 29052 7871
rect 29000 7828 29052 7837
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 30012 7692 30064 7744
rect 38200 7735 38252 7744
rect 38200 7701 38209 7735
rect 38209 7701 38243 7735
rect 38243 7701 38252 7735
rect 38200 7692 38252 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 32772 7488 32824 7540
rect 1676 7352 1728 7404
rect 18788 7352 18840 7404
rect 33140 7395 33192 7404
rect 33140 7361 33149 7395
rect 33149 7361 33183 7395
rect 33183 7361 33192 7395
rect 33140 7352 33192 7361
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 14924 7148 14976 7200
rect 34428 7148 34480 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 8392 6264 8444 6316
rect 5540 6060 5592 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 8392 5899 8444 5908
rect 8392 5865 8401 5899
rect 8401 5865 8435 5899
rect 8435 5865 8444 5899
rect 8392 5856 8444 5865
rect 1952 5720 2004 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 13636 5652 13688 5704
rect 29828 5652 29880 5704
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 7656 4768 7708 4820
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 32496 4564 32548 4616
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 35348 4428 35400 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 664 4088 716 4140
rect 36452 4088 36504 4140
rect 38016 4131 38068 4140
rect 38016 4097 38025 4131
rect 38025 4097 38059 4131
rect 38059 4097 38068 4131
rect 38016 4088 38068 4097
rect 7564 3952 7616 4004
rect 36912 3884 36964 3936
rect 38200 3927 38252 3936
rect 38200 3893 38209 3927
rect 38209 3893 38243 3927
rect 38243 3893 38252 3927
rect 38200 3884 38252 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 5632 3680 5684 3732
rect 33784 3680 33836 3732
rect 5724 3544 5776 3596
rect 28632 3544 28684 3596
rect 37464 3519 37516 3528
rect 20 3408 72 3460
rect 17868 3408 17920 3460
rect 34520 3408 34572 3460
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 38660 3408 38712 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 13728 3068 13780 3120
rect 5540 3000 5592 3052
rect 17316 3068 17368 3120
rect 17868 3068 17920 3120
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 38016 3136 38068 3188
rect 36912 3043 36964 3052
rect 35440 2932 35492 2984
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 34428 2864 34480 2916
rect 1584 2796 1636 2848
rect 3884 2796 3936 2848
rect 16120 2839 16172 2848
rect 16120 2805 16129 2839
rect 16129 2805 16163 2839
rect 16163 2805 16172 2839
rect 16120 2796 16172 2805
rect 16764 2796 16816 2848
rect 32312 2796 32364 2848
rect 37372 2796 37424 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4712 2592 4764 2644
rect 5816 2592 5868 2644
rect 6920 2592 6972 2644
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 7196 2592 7248 2601
rect 14188 2592 14240 2644
rect 16672 2592 16724 2644
rect 20168 2592 20220 2644
rect 23112 2592 23164 2644
rect 23848 2592 23900 2644
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 28724 2592 28776 2644
rect 34520 2592 34572 2644
rect 9220 2524 9272 2576
rect 4620 2456 4672 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 1952 2388 2004 2440
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 3240 2388 3292 2440
rect 5172 2388 5224 2440
rect 6460 2388 6512 2440
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 16120 2524 16172 2576
rect 20536 2524 20588 2576
rect 23480 2524 23532 2576
rect 29276 2524 29328 2576
rect 37188 2524 37240 2576
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11612 2388 11664 2440
rect 12900 2388 12952 2440
rect 13544 2388 13596 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 16764 2388 16816 2440
rect 18052 2388 18104 2440
rect 21180 2456 21232 2508
rect 19340 2388 19392 2440
rect 19984 2388 20036 2440
rect 21272 2388 21324 2440
rect 17776 2320 17828 2372
rect 1400 2252 1452 2304
rect 9680 2252 9732 2304
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 14832 2252 14884 2304
rect 16120 2252 16172 2304
rect 16764 2252 16816 2304
rect 17500 2252 17552 2304
rect 18052 2252 18104 2304
rect 30012 2456 30064 2508
rect 22560 2388 22612 2440
rect 23204 2388 23256 2440
rect 24492 2388 24544 2440
rect 25780 2431 25832 2440
rect 25780 2397 25789 2431
rect 25789 2397 25823 2431
rect 25823 2397 25832 2431
rect 25780 2388 25832 2397
rect 27068 2388 27120 2440
rect 27712 2388 27764 2440
rect 29000 2388 29052 2440
rect 30380 2431 30432 2440
rect 30380 2397 30389 2431
rect 30389 2397 30423 2431
rect 30423 2397 30432 2431
rect 30380 2388 30432 2397
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 35992 2456 36044 2508
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 36636 2431 36688 2440
rect 35900 2388 35952 2397
rect 36636 2397 36645 2431
rect 36645 2397 36679 2431
rect 36679 2397 36688 2431
rect 36636 2388 36688 2397
rect 23112 2320 23164 2372
rect 29828 2320 29880 2372
rect 34152 2320 34204 2372
rect 35348 2320 35400 2372
rect 25136 2252 25188 2304
rect 30288 2252 30340 2304
rect 30932 2252 30984 2304
rect 32220 2252 32272 2304
rect 33508 2252 33560 2304
rect 36820 2295 36872 2304
rect 36820 2261 36829 2295
rect 36829 2261 36863 2295
rect 36863 2261 36872 2295
rect 36820 2252 36872 2261
rect 37004 2252 37056 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 12992 2048 13044 2100
rect 17040 2048 17092 2100
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2056 39222 2360 39250
rect 676 37398 704 39200
rect 1964 39114 1992 39200
rect 2056 39114 2084 39222
rect 1964 39086 2084 39114
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 664 37392 716 37398
rect 664 37334 716 37340
rect 1596 37330 1624 38791
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1674 36952 1730 36961
rect 1674 36887 1730 36896
rect 1688 36854 1716 36887
rect 1676 36848 1728 36854
rect 1676 36790 1728 36796
rect 1768 36168 1820 36174
rect 1766 36136 1768 36145
rect 1820 36136 1822 36145
rect 1766 36071 1822 36080
rect 1676 35760 1728 35766
rect 1674 35728 1676 35737
rect 1768 35760 1820 35766
rect 1728 35728 1730 35737
rect 1768 35702 1820 35708
rect 1674 35663 1730 35672
rect 1780 34746 1808 35702
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 28762 1624 34546
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1768 32768 1820 32774
rect 1766 32736 1768 32745
rect 1820 32736 1822 32745
rect 1766 32671 1822 32680
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30598 1808 30631
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1780 29345 1808 29582
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1860 29164 1912 29170
rect 1860 29106 1912 29112
rect 1768 29028 1820 29034
rect 1768 28970 1820 28976
rect 1584 28756 1636 28762
rect 1584 28698 1636 28704
rect 1780 28665 1808 28970
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 27305 1808 27406
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1780 25945 1808 26318
rect 1766 25936 1822 25945
rect 1766 25871 1822 25880
rect 1768 24608 1820 24614
rect 1766 24576 1768 24585
rect 1820 24576 1822 24585
rect 1766 24511 1822 24520
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22545 1716 22578
rect 1674 22536 1730 22545
rect 1674 22471 1730 22480
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21554 1624 21830
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21185 1808 21286
rect 1766 21176 1822 21185
rect 1766 21111 1822 21120
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1872 20346 1900 29106
rect 1964 22030 1992 37198
rect 2332 36854 2360 39222
rect 2594 39200 2650 39800
rect 3422 39536 3478 39545
rect 3422 39471 3478 39480
rect 2608 37210 2636 39200
rect 2870 37496 2926 37505
rect 2870 37431 2926 37440
rect 2608 37182 2820 37210
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2320 36848 2372 36854
rect 2320 36790 2372 36796
rect 2688 36712 2740 36718
rect 2688 36654 2740 36660
rect 2700 36242 2728 36654
rect 2688 36236 2740 36242
rect 2688 36178 2740 36184
rect 2412 36100 2464 36106
rect 2412 36042 2464 36048
rect 2504 36100 2556 36106
rect 2504 36042 2556 36048
rect 2424 35601 2452 36042
rect 2410 35592 2466 35601
rect 2410 35527 2466 35536
rect 2516 33658 2544 36042
rect 2700 35766 2728 36178
rect 2688 35760 2740 35766
rect 2688 35702 2740 35708
rect 2884 35086 2912 37431
rect 3332 36916 3384 36922
rect 3332 36858 3384 36864
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 2872 35080 2924 35086
rect 2872 35022 2924 35028
rect 2964 34944 3016 34950
rect 2964 34886 3016 34892
rect 2504 33652 2556 33658
rect 2504 33594 2556 33600
rect 2976 32910 3004 34886
rect 2964 32904 3016 32910
rect 2964 32846 3016 32852
rect 3160 30734 3188 36518
rect 3344 35834 3372 36858
rect 3436 36786 3464 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 24596 39222 24808 39250
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3424 36780 3476 36786
rect 3424 36722 3476 36728
rect 3804 36378 3832 37198
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4620 37392 4672 37398
rect 4620 37334 4672 37340
rect 4068 37256 4120 37262
rect 4068 37198 4120 37204
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3792 36372 3844 36378
rect 3792 36314 3844 36320
rect 3424 36236 3476 36242
rect 3424 36178 3476 36184
rect 3332 35828 3384 35834
rect 3332 35770 3384 35776
rect 3240 35692 3292 35698
rect 3240 35634 3292 35640
rect 3252 33862 3280 35634
rect 3240 33856 3292 33862
rect 3240 33798 3292 33804
rect 3148 30728 3200 30734
rect 3148 30670 3200 30676
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 3436 21078 3464 36178
rect 3884 36032 3936 36038
rect 3884 35974 3936 35980
rect 3896 31346 3924 35974
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 1780 20318 1900 20346
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 19145 1624 19246
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1780 18970 1808 20318
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1584 17128 1636 17134
rect 1582 17096 1584 17105
rect 1636 17096 1638 17105
rect 1582 17031 1638 17040
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 9178 1624 16594
rect 1688 15026 1716 18702
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 4080 17882 4108 37198
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 37334
rect 5184 37330 5212 39200
rect 5828 37330 5856 39200
rect 5172 37324 5224 37330
rect 5172 37266 5224 37272
rect 5816 37324 5868 37330
rect 5816 37266 5868 37272
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 6644 37256 6696 37262
rect 6644 37198 6696 37204
rect 5080 37188 5132 37194
rect 5080 37130 5132 37136
rect 5092 36922 5120 37130
rect 5080 36916 5132 36922
rect 5080 36858 5132 36864
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5460 28694 5488 37198
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5632 36644 5684 36650
rect 5632 36586 5684 36592
rect 5644 35086 5672 36586
rect 5828 36582 5856 37062
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 6458 36272 6514 36281
rect 6458 36207 6514 36216
rect 6472 36174 6500 36207
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 5724 36032 5776 36038
rect 5724 35974 5776 35980
rect 5632 35080 5684 35086
rect 5632 35022 5684 35028
rect 5736 32910 5764 35974
rect 6656 35154 6684 37198
rect 7116 36854 7144 39200
rect 7748 37460 7800 37466
rect 7748 37402 7800 37408
rect 7104 36848 7156 36854
rect 7010 36816 7066 36825
rect 7104 36790 7156 36796
rect 7010 36751 7012 36760
rect 7064 36751 7066 36760
rect 7012 36722 7064 36728
rect 7024 36242 7052 36722
rect 7472 36576 7524 36582
rect 7472 36518 7524 36524
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 7484 36242 7512 36518
rect 7012 36236 7064 36242
rect 7012 36178 7064 36184
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7564 36168 7616 36174
rect 7564 36110 7616 36116
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 6644 35148 6696 35154
rect 6644 35090 6696 35096
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5908 32428 5960 32434
rect 5908 32370 5960 32376
rect 5920 29510 5948 32370
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 6656 29238 6684 35090
rect 6828 35012 6880 35018
rect 6828 34954 6880 34960
rect 6840 31906 6868 34954
rect 7484 33590 7512 35974
rect 7472 33584 7524 33590
rect 7472 33526 7524 33532
rect 7576 32842 7604 36110
rect 7564 32836 7616 32842
rect 7564 32778 7616 32784
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 6840 31878 6960 31906
rect 6932 31822 6960 31878
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 6644 29232 6696 29238
rect 6644 29174 6696 29180
rect 5448 28688 5500 28694
rect 5448 28630 5500 28636
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5460 25906 5488 28630
rect 6840 28082 6868 31758
rect 7300 29646 7328 32710
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 7576 29034 7604 29582
rect 7668 29170 7696 36518
rect 7760 36174 7788 37402
rect 8300 36712 8352 36718
rect 8404 36700 8432 39200
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8352 36672 8432 36700
rect 8300 36654 8352 36660
rect 8300 36236 8352 36242
rect 8300 36178 8352 36184
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7840 36032 7892 36038
rect 7840 35974 7892 35980
rect 7852 35290 7880 35974
rect 7840 35284 7892 35290
rect 7840 35226 7892 35232
rect 8312 34610 8340 36178
rect 8496 35154 8524 37198
rect 9048 36922 9076 39200
rect 10336 37346 10364 39200
rect 10244 37330 10364 37346
rect 10232 37324 10364 37330
rect 10284 37318 10364 37324
rect 10506 37360 10562 37369
rect 11624 37330 11652 39200
rect 12268 37330 12296 39200
rect 10506 37295 10562 37304
rect 11612 37324 11664 37330
rect 10232 37266 10284 37272
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 9128 37188 9180 37194
rect 9128 37130 9180 37136
rect 8668 36916 8720 36922
rect 8668 36858 8720 36864
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 8574 36680 8630 36689
rect 8574 36615 8576 36624
rect 8628 36615 8630 36624
rect 8576 36586 8628 36592
rect 8576 35760 8628 35766
rect 8576 35702 8628 35708
rect 8484 35148 8536 35154
rect 8484 35090 8536 35096
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 8300 34604 8352 34610
rect 8300 34546 8352 34552
rect 8496 34202 8524 34614
rect 8484 34196 8536 34202
rect 8484 34138 8536 34144
rect 8208 33856 8260 33862
rect 8208 33798 8260 33804
rect 8220 31385 8248 33798
rect 8588 33658 8616 35702
rect 8680 35086 8708 36858
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 8852 36576 8904 36582
rect 9048 36553 9076 36722
rect 8852 36518 8904 36524
rect 9034 36544 9090 36553
rect 8864 35630 8892 36518
rect 9034 36479 9090 36488
rect 8852 35624 8904 35630
rect 8852 35566 8904 35572
rect 8864 35154 8892 35566
rect 8852 35148 8904 35154
rect 8852 35090 8904 35096
rect 8668 35080 8720 35086
rect 8668 35022 8720 35028
rect 8668 34740 8720 34746
rect 8668 34682 8720 34688
rect 8576 33652 8628 33658
rect 8576 33594 8628 33600
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8312 32473 8340 33458
rect 8392 32768 8444 32774
rect 8392 32710 8444 32716
rect 8298 32464 8354 32473
rect 8298 32399 8354 32408
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8206 31376 8262 31385
rect 8206 31311 8262 31320
rect 8312 30802 8340 31622
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8404 30666 8432 32710
rect 8680 32230 8708 34682
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8944 31952 8996 31958
rect 8944 31894 8996 31900
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8496 30802 8524 31078
rect 8484 30796 8536 30802
rect 8484 30738 8536 30744
rect 8392 30660 8444 30666
rect 8392 30602 8444 30608
rect 8208 30592 8260 30598
rect 8208 30534 8260 30540
rect 8220 29850 8248 30534
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7656 29164 7708 29170
rect 7656 29106 7708 29112
rect 7564 29028 7616 29034
rect 7564 28970 7616 28976
rect 7760 28150 7788 29582
rect 8220 28626 8248 29786
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7944 28218 7972 28494
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 8220 28218 8248 28426
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 7932 28212 7984 28218
rect 7932 28154 7984 28160
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 6840 27418 6868 28018
rect 6656 27390 6868 27418
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5000 24818 5028 25638
rect 6656 25158 6684 27390
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6736 26512 6788 26518
rect 6736 26454 6788 26460
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6656 21962 6684 25094
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6748 21554 6776 26454
rect 6840 22030 6868 27270
rect 7116 25294 7144 28018
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7760 25498 7788 25842
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 8404 24818 8432 28358
rect 8956 25770 8984 31894
rect 9048 31346 9076 33934
rect 9140 31822 9168 37130
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 9220 36916 9272 36922
rect 9220 36858 9272 36864
rect 9232 36106 9260 36858
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9220 36100 9272 36106
rect 9220 36042 9272 36048
rect 9220 34536 9272 34542
rect 9324 34513 9352 36110
rect 9404 34944 9456 34950
rect 9404 34886 9456 34892
rect 9416 34542 9444 34886
rect 9404 34536 9456 34542
rect 9220 34478 9272 34484
rect 9310 34504 9366 34513
rect 9232 33402 9260 34478
rect 9404 34478 9456 34484
rect 9310 34439 9366 34448
rect 9404 33924 9456 33930
rect 9404 33866 9456 33872
rect 9416 33522 9444 33866
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9600 33658 9628 33798
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9404 33516 9456 33522
rect 9404 33458 9456 33464
rect 9232 33374 9444 33402
rect 9220 32428 9272 32434
rect 9220 32370 9272 32376
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 9232 31482 9260 32370
rect 9220 31476 9272 31482
rect 9220 31418 9272 31424
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 9324 29782 9352 31282
rect 9312 29776 9364 29782
rect 9312 29718 9364 29724
rect 9416 29510 9444 33374
rect 9692 32910 9720 37062
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9784 36310 9812 36654
rect 9772 36304 9824 36310
rect 9772 36246 9824 36252
rect 10060 36174 10088 37198
rect 10232 37120 10284 37126
rect 10232 37062 10284 37068
rect 10244 36786 10272 37062
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10140 36576 10192 36582
rect 10138 36544 10140 36553
rect 10192 36544 10194 36553
rect 10138 36479 10194 36488
rect 10140 36304 10192 36310
rect 10140 36246 10192 36252
rect 10048 36168 10100 36174
rect 10048 36110 10100 36116
rect 10152 35465 10180 36246
rect 10138 35456 10194 35465
rect 10138 35391 10194 35400
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9784 34746 9812 34886
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 9784 34474 9812 34682
rect 9772 34468 9824 34474
rect 9772 34410 9824 34416
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9784 32842 9812 33798
rect 10060 33504 10088 34002
rect 10152 33998 10180 34342
rect 10244 34202 10272 36722
rect 10324 36576 10376 36582
rect 10324 36518 10376 36524
rect 10336 36310 10364 36518
rect 10324 36304 10376 36310
rect 10324 36246 10376 36252
rect 10520 36242 10548 37295
rect 11612 37266 11664 37272
rect 11796 37324 11848 37330
rect 11796 37266 11848 37272
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 11704 37256 11756 37262
rect 11702 37224 11704 37233
rect 11756 37224 11758 37233
rect 11702 37159 11758 37168
rect 11808 36961 11836 37266
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 11980 37120 12032 37126
rect 11980 37062 12032 37068
rect 11794 36952 11850 36961
rect 11072 36910 11376 36938
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 10416 36168 10468 36174
rect 10416 36110 10468 36116
rect 10336 36009 10364 36110
rect 10428 36038 10456 36110
rect 10600 36100 10652 36106
rect 10600 36042 10652 36048
rect 10416 36032 10468 36038
rect 10322 36000 10378 36009
rect 10416 35974 10468 35980
rect 10322 35935 10378 35944
rect 10612 35873 10640 36042
rect 10598 35864 10654 35873
rect 10598 35799 10654 35808
rect 10324 35760 10376 35766
rect 10324 35702 10376 35708
rect 10336 35290 10364 35702
rect 10888 35329 10916 36722
rect 11072 36582 11100 36910
rect 11152 36848 11204 36854
rect 11152 36790 11204 36796
rect 11060 36576 11112 36582
rect 11060 36518 11112 36524
rect 11058 36136 11114 36145
rect 10968 36100 11020 36106
rect 11058 36071 11114 36080
rect 10968 36042 11020 36048
rect 10980 35562 11008 36042
rect 10968 35556 11020 35562
rect 10968 35498 11020 35504
rect 10874 35320 10930 35329
rect 10324 35284 10376 35290
rect 11072 35290 11100 36071
rect 11164 35630 11192 36790
rect 11242 36000 11298 36009
rect 11242 35935 11298 35944
rect 11256 35698 11284 35935
rect 11244 35692 11296 35698
rect 11244 35634 11296 35640
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 11244 35556 11296 35562
rect 11244 35498 11296 35504
rect 10874 35255 10930 35264
rect 11060 35284 11112 35290
rect 10324 35226 10376 35232
rect 11060 35226 11112 35232
rect 10966 35184 11022 35193
rect 10966 35119 11022 35128
rect 10980 35086 11008 35119
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10692 34672 10744 34678
rect 10690 34640 10692 34649
rect 10744 34640 10746 34649
rect 10690 34575 10746 34584
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10140 33516 10192 33522
rect 10060 33476 10140 33504
rect 10140 33458 10192 33464
rect 9864 33312 9916 33318
rect 9864 33254 9916 33260
rect 9772 32836 9824 32842
rect 9772 32778 9824 32784
rect 9876 32502 9904 33254
rect 10152 33017 10180 33458
rect 10138 33008 10194 33017
rect 10138 32943 10194 32952
rect 9864 32496 9916 32502
rect 9864 32438 9916 32444
rect 9772 32360 9824 32366
rect 9772 32302 9824 32308
rect 9784 32026 9812 32302
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9508 29646 9536 29990
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9232 27130 9260 27406
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9416 26994 9444 29446
rect 9692 27606 9720 29582
rect 9784 29034 9812 31962
rect 10048 31680 10100 31686
rect 10048 31622 10100 31628
rect 10060 30666 10088 31622
rect 10140 30796 10192 30802
rect 10140 30738 10192 30744
rect 10048 30660 10100 30666
rect 10048 30602 10100 30608
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9968 29714 9996 30126
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9772 29028 9824 29034
rect 9772 28970 9824 28976
rect 10060 28150 10088 29106
rect 10048 28144 10100 28150
rect 10048 28086 10100 28092
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9784 26586 9812 28018
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9324 26042 9352 26318
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 8944 25764 8996 25770
rect 8944 25706 8996 25712
rect 9784 25498 9812 26522
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 8668 25424 8720 25430
rect 8668 25366 8720 25372
rect 8680 24818 8708 25366
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 24206 7328 24550
rect 8404 24410 8432 24754
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 9324 24274 9352 24550
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 6840 20466 6868 21830
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 7300 20330 7328 22578
rect 7760 22098 7788 24142
rect 9140 23322 9168 24142
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 8312 18426 8340 19314
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 1860 17808 1912 17814
rect 1766 17776 1822 17785
rect 1860 17750 1912 17756
rect 1766 17711 1822 17720
rect 1872 17202 1900 17750
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 7410 1716 14962
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1780 14278 1808 14311
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1780 13705 1808 13874
rect 1766 13696 1822 13705
rect 1766 13631 1822 13640
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12345 1808 12582
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10305 1808 10610
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1768 8968 1820 8974
rect 1766 8936 1768 8945
rect 1820 8936 1822 8945
rect 1766 8871 1822 8880
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7585 1808 7686
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6905 1624 7278
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1964 5778 1992 17614
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 8496 14074 8524 15914
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8312 12850 8340 13806
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5545 1624 5646
rect 1582 5536 1638 5545
rect 1582 5471 1638 5480
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1780 4185 1808 4558
rect 1766 4176 1822 4185
rect 664 4140 716 4146
rect 1766 4111 1822 4120
rect 664 4082 716 4088
rect 20 3460 72 3466
rect 20 3402 72 3408
rect 32 800 60 3402
rect 676 800 704 4082
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1780 3398 1808 3431
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 1596 2446 1624 2790
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 1400 2304 1452 2310
rect 1400 2246 1452 2252
rect 18 200 74 800
rect 662 200 718 800
rect 1412 785 1440 2246
rect 1964 800 1992 2382
rect 3160 2145 3188 2382
rect 3146 2136 3202 2145
rect 3146 2071 3202 2080
rect 3252 800 3280 2382
rect 3896 800 3924 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 12174
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4724 2650 4752 9522
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 3058 5580 6054
rect 5644 3738 5672 8366
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5736 3602 5764 8298
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5828 2650 5856 9454
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8498 7144 9318
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 2650 6960 7822
rect 7208 2650 7236 9998
rect 7576 4010 7604 11698
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7668 4826 7696 11086
rect 8772 10810 8800 14894
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8864 9654 8892 23054
rect 9140 22506 9168 23258
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9232 21146 9260 22578
rect 9324 22234 9352 23054
rect 9312 22228 9364 22234
rect 9312 22170 9364 22176
rect 10152 22094 10180 30738
rect 10244 30258 10272 33934
rect 10324 33856 10376 33862
rect 10324 33798 10376 33804
rect 10336 33590 10364 33798
rect 10324 33584 10376 33590
rect 10324 33526 10376 33532
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10428 31482 10456 33526
rect 10796 33425 10824 35022
rect 10876 35012 10928 35018
rect 10876 34954 10928 34960
rect 10888 33998 10916 34954
rect 11152 34536 11204 34542
rect 11152 34478 11204 34484
rect 10968 34468 11020 34474
rect 10968 34410 11020 34416
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10782 33416 10838 33425
rect 10782 33351 10838 33360
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10416 31476 10468 31482
rect 10416 31418 10468 31424
rect 10416 30932 10468 30938
rect 10416 30874 10468 30880
rect 10428 30666 10456 30874
rect 10416 30660 10468 30666
rect 10416 30602 10468 30608
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10324 27940 10376 27946
rect 10324 27882 10376 27888
rect 10336 26450 10364 27882
rect 10428 27674 10456 30602
rect 10612 30394 10640 32846
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 10506 28792 10562 28801
rect 10506 28727 10508 28736
rect 10560 28727 10562 28736
rect 10508 28698 10560 28704
rect 10508 28008 10560 28014
rect 10508 27950 10560 27956
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10428 26314 10456 27270
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10060 22066 10180 22094
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 17202 9168 17614
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8404 5914 8432 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 9232 2582 9260 12786
rect 9324 9654 9352 18634
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9968 17270 9996 17546
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 10060 16522 10088 22066
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9508 10062 9536 11222
rect 10152 10266 10180 21422
rect 10244 17746 10272 25366
rect 10336 24732 10364 26250
rect 10520 25838 10548 27950
rect 10612 27470 10640 30330
rect 10796 28082 10824 33351
rect 10888 31754 10916 33934
rect 10980 33046 11008 34410
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 11072 33289 11100 33458
rect 11058 33280 11114 33289
rect 11058 33215 11114 33224
rect 10968 33040 11020 33046
rect 10968 32982 11020 32988
rect 11072 31822 11100 33215
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 10888 31726 11008 31754
rect 10980 31686 11008 31726
rect 10876 31680 10928 31686
rect 10876 31622 10928 31628
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10888 30666 10916 31622
rect 10980 31346 11008 31622
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 11058 31240 11114 31249
rect 11058 31175 11060 31184
rect 11112 31175 11114 31184
rect 11060 31146 11112 31152
rect 11164 30870 11192 34478
rect 11152 30864 11204 30870
rect 11152 30806 11204 30812
rect 11256 30802 11284 35498
rect 11348 32026 11376 36910
rect 11992 36922 12020 37062
rect 11794 36887 11850 36896
rect 11980 36916 12032 36922
rect 11980 36858 12032 36864
rect 11704 36712 11756 36718
rect 11704 36654 11756 36660
rect 11716 36378 11744 36654
rect 12452 36650 12480 37198
rect 12440 36644 12492 36650
rect 12440 36586 12492 36592
rect 12532 36576 12584 36582
rect 11886 36544 11942 36553
rect 11886 36479 11942 36488
rect 12070 36544 12126 36553
rect 12532 36518 12584 36524
rect 12624 36576 12676 36582
rect 12624 36518 12676 36524
rect 12070 36479 12126 36488
rect 11900 36378 11928 36479
rect 11704 36372 11756 36378
rect 11704 36314 11756 36320
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11612 35760 11664 35766
rect 11612 35702 11664 35708
rect 11624 34610 11652 35702
rect 11716 35494 11744 36042
rect 11900 35578 11928 36314
rect 12084 36106 12112 36479
rect 12544 36242 12572 36518
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12072 36100 12124 36106
rect 12072 36042 12124 36048
rect 12164 36100 12216 36106
rect 12164 36042 12216 36048
rect 12176 35873 12204 36042
rect 12162 35864 12218 35873
rect 12162 35799 12218 35808
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12440 35692 12492 35698
rect 12636 35680 12664 36518
rect 12492 35652 12664 35680
rect 12440 35634 12492 35640
rect 11808 35550 11928 35578
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11428 34196 11480 34202
rect 11428 34138 11480 34144
rect 11440 33674 11468 34138
rect 11808 33998 11836 35550
rect 12084 35494 12112 35634
rect 12808 35556 12860 35562
rect 12808 35498 12860 35504
rect 11888 35488 11940 35494
rect 11888 35430 11940 35436
rect 12072 35488 12124 35494
rect 12820 35442 12848 35498
rect 12072 35430 12124 35436
rect 11900 35154 11928 35430
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 11980 35080 12032 35086
rect 11980 35022 12032 35028
rect 11992 34746 12020 35022
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 11888 34672 11940 34678
rect 11886 34640 11888 34649
rect 11940 34640 11942 34649
rect 11886 34575 11942 34584
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11980 33924 12032 33930
rect 11980 33866 12032 33872
rect 11992 33833 12020 33866
rect 11978 33824 12034 33833
rect 11978 33759 12034 33768
rect 11440 33646 12020 33674
rect 11992 33590 12020 33646
rect 11980 33584 12032 33590
rect 11980 33526 12032 33532
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 11702 33144 11758 33153
rect 11702 33079 11758 33088
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11336 32020 11388 32026
rect 11336 31962 11388 31968
rect 11244 30796 11296 30802
rect 11244 30738 11296 30744
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 10874 29880 10930 29889
rect 10874 29815 10930 29824
rect 10784 28076 10836 28082
rect 10784 28018 10836 28024
rect 10888 27946 10916 29815
rect 11256 29578 11284 30058
rect 11152 29572 11204 29578
rect 11152 29514 11204 29520
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 10980 29073 11008 29106
rect 10966 29064 11022 29073
rect 10966 28999 11022 29008
rect 11164 28422 11192 29514
rect 11244 28960 11296 28966
rect 11244 28902 11296 28908
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10428 24954 10456 25162
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10416 24744 10468 24750
rect 10336 24704 10416 24732
rect 10416 24686 10468 24692
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10244 15570 10272 15982
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10428 11898 10456 24686
rect 10520 12986 10548 25774
rect 10888 22094 10916 27610
rect 11164 27538 11192 28358
rect 11152 27532 11204 27538
rect 11152 27474 11204 27480
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 11164 25906 11192 26930
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 11060 25764 11112 25770
rect 11060 25706 11112 25712
rect 10968 24676 11020 24682
rect 11072 24664 11100 25706
rect 11020 24636 11100 24664
rect 10968 24618 11020 24624
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11072 22574 11100 24142
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10888 22066 11008 22094
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10888 21486 10916 21830
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10612 15910 10640 17682
rect 10980 17610 11008 22066
rect 11072 21622 11100 22374
rect 11256 22098 11284 28902
rect 11348 28694 11376 30194
rect 11440 29102 11468 30738
rect 11532 29714 11560 32914
rect 11716 31890 11744 33079
rect 11992 32842 12020 33254
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 12084 32722 12112 35430
rect 12636 35414 12848 35442
rect 12636 35154 12664 35414
rect 12912 35170 12940 37198
rect 13556 36922 13584 39200
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 13464 36242 13492 36858
rect 13648 36786 13676 37130
rect 14844 37126 14872 39200
rect 15200 37392 15252 37398
rect 15200 37334 15252 37340
rect 15016 37188 15068 37194
rect 15016 37130 15068 37136
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 13636 36780 13688 36786
rect 13636 36722 13688 36728
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13452 36236 13504 36242
rect 13452 36178 13504 36184
rect 13464 35834 13492 36178
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 13544 35828 13596 35834
rect 13544 35770 13596 35776
rect 12624 35148 12676 35154
rect 12624 35090 12676 35096
rect 12820 35142 12940 35170
rect 12164 34944 12216 34950
rect 12164 34886 12216 34892
rect 12176 33930 12204 34886
rect 12820 34490 12848 35142
rect 12348 34468 12400 34474
rect 12348 34410 12400 34416
rect 12636 34462 12848 34490
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 12256 33108 12308 33114
rect 12256 33050 12308 33056
rect 12176 32842 12204 33050
rect 12164 32836 12216 32842
rect 12164 32778 12216 32784
rect 12268 32774 12296 33050
rect 11992 32694 12112 32722
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 11796 32360 11848 32366
rect 11796 32302 11848 32308
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11716 31346 11744 31826
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11808 29850 11836 32302
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11428 29096 11480 29102
rect 11428 29038 11480 29044
rect 11336 28688 11388 28694
rect 11336 28630 11388 28636
rect 11348 24274 11376 28630
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 11440 21146 11468 21966
rect 11532 21593 11560 29650
rect 11808 28762 11836 29786
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11624 25226 11652 28494
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11704 25220 11756 25226
rect 11704 25162 11756 25168
rect 11624 24410 11652 25162
rect 11716 24410 11744 25162
rect 11900 24750 11928 30534
rect 11992 30258 12020 32694
rect 12360 32298 12388 34410
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 12544 32570 12572 33322
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12348 32292 12400 32298
rect 12348 32234 12400 32240
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12268 31958 12296 32166
rect 12256 31952 12308 31958
rect 12256 31894 12308 31900
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11992 27402 12020 29990
rect 12084 28966 12112 31826
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 12072 28960 12124 28966
rect 12072 28902 12124 28908
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 12176 27334 12204 29038
rect 12268 28558 12296 31894
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 11992 26518 12020 26930
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 11980 26512 12032 26518
rect 11980 26454 12032 26460
rect 12084 25974 12112 26726
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11716 22642 11744 24142
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11518 21584 11574 21593
rect 11518 21519 11574 21528
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 17882 11100 18634
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10980 17134 11008 17546
rect 11256 17338 11284 17614
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 11440 16574 11468 21082
rect 11624 19530 11652 22510
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11716 19718 11744 20198
rect 11900 19786 11928 22918
rect 11992 21894 12020 25842
rect 12176 25770 12204 27270
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12164 25764 12216 25770
rect 12164 25706 12216 25712
rect 12268 25226 12296 25978
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12268 23662 12296 25162
rect 12360 24886 12388 28358
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12452 26314 12480 27950
rect 12544 27402 12572 32506
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12360 22710 12388 24686
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 12452 23322 12480 23734
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11624 19502 11744 19530
rect 11440 16546 11652 16574
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16114 10824 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 15094 10916 15302
rect 11440 15162 11468 15982
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 15162 11560 15438
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10888 13938 10916 15030
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 11624 12918 11652 16546
rect 11716 15570 11744 19502
rect 11808 18358 11836 19722
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11992 16250 12020 18294
rect 12084 17746 12112 22034
rect 12544 21554 12572 27338
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12360 18834 12388 19314
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12176 17610 12204 18566
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12268 15638 12296 17682
rect 12544 17202 12572 18838
rect 12636 18766 12664 34462
rect 13004 34134 13032 35770
rect 13556 35714 13584 35770
rect 13372 35686 13584 35714
rect 13174 35320 13230 35329
rect 13174 35255 13230 35264
rect 12900 34128 12952 34134
rect 12898 34096 12900 34105
rect 12992 34128 13044 34134
rect 12952 34096 12954 34105
rect 12992 34070 13044 34076
rect 12898 34031 12954 34040
rect 12808 33924 12860 33930
rect 12808 33866 12860 33872
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 30666 12756 32166
rect 12820 31890 12848 33866
rect 13188 33697 13216 35255
rect 13268 35080 13320 35086
rect 13372 35068 13400 35686
rect 13634 35320 13690 35329
rect 13452 35284 13504 35290
rect 13634 35255 13636 35264
rect 13452 35226 13504 35232
rect 13688 35255 13690 35264
rect 13636 35226 13688 35232
rect 13320 35040 13400 35068
rect 13268 35022 13320 35028
rect 13280 34746 13308 35022
rect 13464 34950 13492 35226
rect 13452 34944 13504 34950
rect 13452 34886 13504 34892
rect 13268 34740 13320 34746
rect 13268 34682 13320 34688
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13174 33688 13230 33697
rect 13174 33623 13230 33632
rect 12808 31884 12860 31890
rect 12808 31826 12860 31832
rect 13188 31822 13216 33623
rect 13280 32910 13308 34682
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13556 34218 13584 34478
rect 13464 34202 13584 34218
rect 13648 34202 13676 34682
rect 13740 34474 13768 36722
rect 13924 36718 13952 36858
rect 13912 36712 13964 36718
rect 13912 36654 13964 36660
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 14844 36310 14872 36518
rect 14832 36304 14884 36310
rect 14832 36246 14884 36252
rect 14832 36168 14884 36174
rect 14832 36110 14884 36116
rect 14844 35698 14872 36110
rect 13820 35692 13872 35698
rect 13820 35634 13872 35640
rect 14832 35692 14884 35698
rect 14832 35634 14884 35640
rect 13832 35494 13860 35634
rect 13912 35624 13964 35630
rect 13912 35566 13964 35572
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13832 35086 13860 35430
rect 13820 35080 13872 35086
rect 13820 35022 13872 35028
rect 13728 34468 13780 34474
rect 13728 34410 13780 34416
rect 13452 34196 13584 34202
rect 13504 34190 13584 34196
rect 13452 34138 13504 34144
rect 13556 33930 13584 34190
rect 13636 34196 13688 34202
rect 13636 34138 13688 34144
rect 13832 33998 13860 35022
rect 13924 34678 13952 35566
rect 14832 35488 14884 35494
rect 14832 35430 14884 35436
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14648 35012 14700 35018
rect 14648 34954 14700 34960
rect 14372 34944 14424 34950
rect 14372 34886 14424 34892
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 13820 33992 13872 33998
rect 14384 33969 14412 34886
rect 14660 34746 14688 34954
rect 14648 34740 14700 34746
rect 14648 34682 14700 34688
rect 14464 34672 14516 34678
rect 14464 34614 14516 34620
rect 13820 33934 13872 33940
rect 14370 33960 14426 33969
rect 13544 33924 13596 33930
rect 14370 33895 14426 33904
rect 13544 33866 13596 33872
rect 14476 33590 14504 34614
rect 14752 34610 14780 35226
rect 14844 34746 14872 35430
rect 14924 35012 14976 35018
rect 14924 34954 14976 34960
rect 14832 34740 14884 34746
rect 14832 34682 14884 34688
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14464 33584 14516 33590
rect 14464 33526 14516 33532
rect 13820 33448 13872 33454
rect 14936 33402 14964 34954
rect 15028 34678 15056 37130
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 15120 34513 15148 37062
rect 15106 34504 15162 34513
rect 15106 34439 15162 34448
rect 15120 33674 15148 34439
rect 15028 33646 15148 33674
rect 15028 33522 15056 33646
rect 15106 33552 15162 33561
rect 15016 33516 15068 33522
rect 15106 33487 15162 33496
rect 15016 33458 15068 33464
rect 13820 33390 13872 33396
rect 13832 33318 13860 33390
rect 14844 33374 14964 33402
rect 13820 33312 13872 33318
rect 13820 33254 13872 33260
rect 13268 32904 13320 32910
rect 13268 32846 13320 32852
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 13280 31754 13308 32846
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 13360 32496 13412 32502
rect 13360 32438 13412 32444
rect 13268 31748 13320 31754
rect 13268 31690 13320 31696
rect 12806 31376 12862 31385
rect 12806 31311 12862 31320
rect 13176 31340 13228 31346
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 12820 30410 12848 31311
rect 13280 31328 13308 31690
rect 13228 31300 13308 31328
rect 13176 31282 13228 31288
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 12728 30382 12848 30410
rect 12728 26994 12756 30382
rect 12808 30252 12860 30258
rect 12808 30194 12860 30200
rect 12820 29345 12848 30194
rect 13096 29714 13124 30534
rect 13188 30297 13216 31282
rect 13372 30666 13400 32438
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13556 32337 13584 32370
rect 13542 32328 13598 32337
rect 13542 32263 13598 32272
rect 13544 31136 13596 31142
rect 13542 31104 13544 31113
rect 13596 31104 13598 31113
rect 13542 31039 13598 31048
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13174 30288 13230 30297
rect 13174 30223 13176 30232
rect 13228 30223 13230 30232
rect 13176 30194 13228 30200
rect 13280 30190 13308 30602
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 13188 29850 13216 30058
rect 13176 29844 13228 29850
rect 13176 29786 13228 29792
rect 13280 29782 13308 30126
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 13268 29776 13320 29782
rect 13268 29718 13320 29724
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12806 29336 12862 29345
rect 12806 29271 12862 29280
rect 12820 28994 12848 29271
rect 12912 29170 12940 29446
rect 13188 29306 13216 29514
rect 13176 29300 13228 29306
rect 13176 29242 13228 29248
rect 13556 29170 13584 29990
rect 13648 29617 13676 32710
rect 13634 29608 13690 29617
rect 13634 29543 13690 29552
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 12820 28966 12940 28994
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12912 28506 12940 28966
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 13004 28626 13032 28902
rect 13740 28762 13768 29174
rect 13832 29102 13860 33254
rect 14004 33040 14056 33046
rect 14004 32982 14056 32988
rect 14016 32434 14044 32982
rect 14462 32872 14518 32881
rect 14462 32807 14464 32816
rect 14516 32807 14518 32816
rect 14464 32778 14516 32784
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14004 32428 14056 32434
rect 14004 32370 14056 32376
rect 14016 31754 14044 32370
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14016 31726 14136 31754
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13924 31346 13952 31622
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 14004 31272 14056 31278
rect 14004 31214 14056 31220
rect 13912 30660 13964 30666
rect 13912 30602 13964 30608
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 12992 28620 13044 28626
rect 12992 28562 13044 28568
rect 13728 28552 13780 28558
rect 12820 27470 12848 28494
rect 12912 28478 13032 28506
rect 13728 28494 13780 28500
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12912 27878 12940 28358
rect 12900 27872 12952 27878
rect 12900 27814 12952 27820
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12728 24682 12756 26726
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12716 24676 12768 24682
rect 12716 24618 12768 24624
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12636 16590 12664 18702
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12728 16182 12756 23462
rect 12820 19786 12848 24686
rect 13004 23118 13032 28478
rect 13082 27840 13138 27849
rect 13082 27775 13138 27784
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13096 22094 13124 27775
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13556 26586 13584 26930
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13740 26382 13768 28494
rect 13924 28150 13952 30602
rect 13912 28144 13964 28150
rect 13912 28086 13964 28092
rect 14016 27962 14044 31214
rect 13832 27934 14044 27962
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13832 25906 13860 27934
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13188 23594 13216 24074
rect 13176 23588 13228 23594
rect 13176 23530 13228 23536
rect 13096 22066 13216 22094
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12820 16794 12848 19722
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19446 13124 19654
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13188 18902 13216 22066
rect 13280 20330 13308 25774
rect 13634 25392 13690 25401
rect 13634 25327 13690 25336
rect 13648 25158 13676 25327
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13740 24342 13768 25094
rect 13832 24818 13860 25842
rect 13924 24818 13952 26250
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 14016 24206 14044 27406
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 22710 14044 24006
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13372 19242 13400 22510
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 13372 18222 13400 19178
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 13004 15502 13032 16934
rect 13280 16726 13308 17138
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15094 13308 15302
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14482 11928 14962
rect 13464 14958 13492 17546
rect 13176 14952 13228 14958
rect 13452 14952 13504 14958
rect 13176 14894 13228 14900
rect 13372 14900 13452 14906
rect 13372 14894 13504 14900
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 13188 13530 13216 14894
rect 13372 14878 13492 14894
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11624 12238 11652 12854
rect 12176 12850 12204 13126
rect 13188 12986 13216 13466
rect 13280 13394 13308 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 10980 8090 11008 10542
rect 13372 9654 13400 14878
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 10606 13492 14758
rect 13556 13546 13584 17682
rect 13648 14822 13676 19926
rect 13740 19310 13768 20266
rect 14108 20058 14136 31726
rect 14384 30433 14412 31758
rect 14370 30424 14426 30433
rect 14370 30359 14426 30368
rect 14752 30326 14780 32710
rect 14844 31482 14872 33374
rect 15120 33114 15148 33487
rect 15212 33114 15240 37334
rect 16132 37330 16160 39200
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 16488 37324 16540 37330
rect 16488 37266 16540 37272
rect 16500 37126 16528 37266
rect 16672 37256 16724 37262
rect 16672 37198 16724 37204
rect 16488 37120 16540 37126
rect 16488 37062 16540 37068
rect 16580 37120 16632 37126
rect 16580 37062 16632 37068
rect 15290 36952 15346 36961
rect 15290 36887 15346 36896
rect 15304 36854 15332 36887
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15384 36712 15436 36718
rect 15384 36654 15436 36660
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 15304 35766 15332 35974
rect 15292 35760 15344 35766
rect 15292 35702 15344 35708
rect 15396 34048 15424 36654
rect 16316 36553 16344 36654
rect 16302 36544 16358 36553
rect 16302 36479 16358 36488
rect 15660 36100 15712 36106
rect 15660 36042 15712 36048
rect 16212 36100 16264 36106
rect 16212 36042 16264 36048
rect 16304 36100 16356 36106
rect 16304 36042 16356 36048
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15488 35154 15516 35430
rect 15476 35148 15528 35154
rect 15476 35090 15528 35096
rect 15568 35012 15620 35018
rect 15568 34954 15620 34960
rect 15580 34649 15608 34954
rect 15566 34640 15622 34649
rect 15566 34575 15622 34584
rect 15566 34232 15622 34241
rect 15672 34202 15700 36042
rect 16224 35834 16252 36042
rect 16212 35828 16264 35834
rect 16212 35770 16264 35776
rect 15936 34536 15988 34542
rect 15936 34478 15988 34484
rect 15566 34167 15568 34176
rect 15620 34167 15622 34176
rect 15660 34196 15712 34202
rect 15568 34138 15620 34144
rect 15660 34138 15712 34144
rect 15304 34020 15424 34048
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15200 33108 15252 33114
rect 15200 33050 15252 33056
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14936 32434 14964 32982
rect 15200 32972 15252 32978
rect 15200 32914 15252 32920
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 14832 31476 14884 31482
rect 14832 31418 14884 31424
rect 14188 30320 14240 30326
rect 14188 30262 14240 30268
rect 14740 30320 14792 30326
rect 14740 30262 14792 30268
rect 14200 28762 14228 30262
rect 14936 30190 14964 31894
rect 15028 31686 15056 32846
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 15212 31278 15240 32914
rect 15304 31414 15332 34020
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15396 32026 15424 33866
rect 15566 33688 15622 33697
rect 15566 33623 15622 33632
rect 15580 33522 15608 33623
rect 15568 33516 15620 33522
rect 15568 33458 15620 33464
rect 15844 32836 15896 32842
rect 15844 32778 15896 32784
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15488 31482 15516 32438
rect 15856 32366 15884 32778
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 15856 32026 15884 32302
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 15844 32020 15896 32026
rect 15844 31962 15896 31968
rect 15764 31793 15792 31962
rect 15750 31784 15806 31793
rect 15750 31719 15806 31728
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15304 30784 15332 31350
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15212 30756 15332 30784
rect 15212 30666 15240 30756
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15304 30326 15332 30602
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15384 30320 15436 30326
rect 15384 30262 15436 30268
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14924 30184 14976 30190
rect 14924 30126 14976 30132
rect 14188 28756 14240 28762
rect 14188 28698 14240 28704
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14200 27130 14228 28086
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14200 24342 14228 25910
rect 14292 25294 14320 27406
rect 14384 26450 14412 27950
rect 14476 26450 14504 30126
rect 15028 30122 15240 30138
rect 15016 30116 15240 30122
rect 15068 30110 15240 30116
rect 15016 30058 15068 30064
rect 14740 29844 14792 29850
rect 14740 29786 14792 29792
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14568 28014 14596 29038
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14464 26444 14516 26450
rect 14464 26386 14516 26392
rect 14384 25498 14412 26386
rect 14476 26042 14504 26386
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14188 24336 14240 24342
rect 14188 24278 14240 24284
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13740 18698 13768 19246
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 14200 18630 14228 24142
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14200 17338 14228 18294
rect 14292 17814 14320 25230
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14384 21962 14412 22510
rect 14568 22094 14596 27950
rect 14752 27674 14780 29786
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 15106 29064 15162 29073
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 14660 24886 14688 25638
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14844 24750 14872 29038
rect 15106 28999 15162 29008
rect 14924 28552 14976 28558
rect 14922 28520 14924 28529
rect 14976 28520 14978 28529
rect 14922 28455 14978 28464
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14568 22066 14688 22094
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14384 18970 14412 21898
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14568 19922 14596 20334
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14660 19428 14688 22066
rect 14752 21690 14780 22714
rect 14844 22506 14872 24686
rect 14936 23186 14964 28455
rect 15120 28234 15148 28999
rect 15212 28422 15240 30110
rect 15304 29034 15332 30262
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15396 28762 15424 30262
rect 15580 30190 15608 30806
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15764 29730 15792 30738
rect 15856 29850 15884 31690
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15764 29702 15884 29730
rect 15476 29572 15528 29578
rect 15476 29514 15528 29520
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15120 28206 15332 28234
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15212 27062 15240 27406
rect 15200 27056 15252 27062
rect 15200 26998 15252 27004
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15120 25906 15148 26862
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 15120 23322 15148 25162
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14660 19400 14780 19428
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18290 14412 18566
rect 14660 18426 14688 18634
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 16182 14044 16526
rect 14752 16250 14780 19400
rect 14844 18358 14872 22170
rect 14936 20505 14964 22510
rect 15028 22234 15056 22714
rect 15304 22642 15332 28206
rect 15384 28144 15436 28150
rect 15384 28086 15436 28092
rect 15396 25498 15424 28086
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15488 22094 15516 29514
rect 15580 26586 15608 29514
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15672 27946 15700 29174
rect 15856 29084 15884 29702
rect 15948 29102 15976 34478
rect 16224 34474 16252 35770
rect 16212 34468 16264 34474
rect 16212 34410 16264 34416
rect 16028 33924 16080 33930
rect 16028 33866 16080 33872
rect 16040 32502 16068 33866
rect 16316 33658 16344 36042
rect 16592 35290 16620 37062
rect 16684 36650 16712 37198
rect 16672 36644 16724 36650
rect 16672 36586 16724 36592
rect 16776 35698 16804 39200
rect 17224 37664 17276 37670
rect 17224 37606 17276 37612
rect 17236 37466 17264 37606
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17038 37224 17094 37233
rect 17038 37159 17094 37168
rect 17776 37188 17828 37194
rect 16856 36644 16908 36650
rect 16856 36586 16908 36592
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16580 35284 16632 35290
rect 16580 35226 16632 35232
rect 16684 35018 16712 35566
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 16672 35012 16724 35018
rect 16672 34954 16724 34960
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16304 33652 16356 33658
rect 16304 33594 16356 33600
rect 16500 33590 16528 33934
rect 16592 33658 16620 34954
rect 16670 34232 16726 34241
rect 16670 34167 16672 34176
rect 16724 34167 16726 34176
rect 16672 34138 16724 34144
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16488 33584 16540 33590
rect 16488 33526 16540 33532
rect 16868 32842 16896 36586
rect 17052 36553 17080 37159
rect 17776 37130 17828 37136
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 17236 36650 17264 37062
rect 17684 36712 17736 36718
rect 17684 36654 17736 36660
rect 17224 36644 17276 36650
rect 17224 36586 17276 36592
rect 17038 36544 17094 36553
rect 17038 36479 17094 36488
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 17132 36236 17184 36242
rect 17132 36178 17184 36184
rect 16120 32836 16172 32842
rect 16120 32778 16172 32784
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16132 32570 16160 32778
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16028 32496 16080 32502
rect 16028 32438 16080 32444
rect 16396 32020 16448 32026
rect 16396 31962 16448 31968
rect 16408 31822 16436 31962
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 15764 29056 15884 29084
rect 15936 29096 15988 29102
rect 15764 28014 15792 29056
rect 15936 29038 15988 29044
rect 16304 29096 16356 29102
rect 16304 29038 16356 29044
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15948 28490 15976 28562
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 15752 28008 15804 28014
rect 15752 27950 15804 27956
rect 15660 27940 15712 27946
rect 15660 27882 15712 27888
rect 15844 27940 15896 27946
rect 15844 27882 15896 27888
rect 15856 27849 15884 27882
rect 15842 27840 15898 27849
rect 15842 27775 15898 27784
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15568 26580 15620 26586
rect 15568 26522 15620 26528
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15488 22066 15608 22094
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 21690 15332 21898
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 14922 20496 14978 20505
rect 14922 20431 14978 20440
rect 14832 18352 14884 18358
rect 14832 18294 14884 18300
rect 14936 16590 14964 20431
rect 15212 19786 15240 20742
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15120 18902 15148 19178
rect 15580 18902 15608 22066
rect 15108 18896 15160 18902
rect 15108 18838 15160 18844
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13740 13870 13768 15914
rect 14384 15706 14412 16118
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14476 15502 14504 15642
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14618 14412 14894
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14476 13938 14504 15438
rect 15672 14482 15700 25910
rect 15948 24818 15976 27338
rect 16040 25158 16068 28494
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15764 22234 15792 23054
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15948 18290 15976 22170
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 13728 13864 13780 13870
rect 13780 13812 13860 13818
rect 13728 13806 13860 13812
rect 13740 13790 13860 13806
rect 13556 13518 13768 13546
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 13648 5710 13676 13398
rect 13740 10742 13768 13518
rect 13832 13462 13860 13790
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15028 12986 15056 13262
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13740 3126 13768 10542
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 14200 2650 14228 11698
rect 15672 11694 15700 13330
rect 16224 12782 16252 27950
rect 16316 24274 16344 29038
rect 16396 25220 16448 25226
rect 16396 25162 16448 25168
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16408 18714 16436 25162
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16500 24886 16528 25094
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16592 24682 16620 31690
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 16684 30326 16712 30534
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16776 27334 16804 32778
rect 16868 31822 16896 32778
rect 16960 32026 16988 36178
rect 17040 36032 17092 36038
rect 17040 35974 17092 35980
rect 17052 35766 17080 35974
rect 17040 35760 17092 35766
rect 17040 35702 17092 35708
rect 17144 34762 17172 36178
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17052 34734 17172 34762
rect 17052 34105 17080 34734
rect 17236 34610 17264 35430
rect 17500 34672 17552 34678
rect 17500 34614 17552 34620
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17132 34400 17184 34406
rect 17132 34342 17184 34348
rect 17038 34096 17094 34105
rect 17038 34031 17094 34040
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17052 33522 17080 33798
rect 17040 33516 17092 33522
rect 17040 33458 17092 33464
rect 17144 32994 17172 34342
rect 17052 32978 17172 32994
rect 17512 32978 17540 34614
rect 17590 33688 17646 33697
rect 17590 33623 17646 33632
rect 17604 33318 17632 33623
rect 17592 33312 17644 33318
rect 17592 33254 17644 33260
rect 17040 32972 17172 32978
rect 17092 32966 17172 32972
rect 17500 32972 17552 32978
rect 17040 32914 17092 32920
rect 17500 32914 17552 32920
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 17316 31204 17368 31210
rect 17316 31146 17368 31152
rect 17038 31104 17094 31113
rect 17038 31039 17094 31048
rect 16856 30932 16908 30938
rect 16856 30874 16908 30880
rect 16868 30394 16896 30874
rect 17052 30394 17080 31039
rect 17328 30598 17356 31146
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 17040 30388 17092 30394
rect 17040 30330 17092 30336
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16868 29850 16896 30194
rect 16856 29844 16908 29850
rect 16856 29786 16908 29792
rect 16948 28960 17000 28966
rect 16948 28902 17000 28908
rect 16960 28626 16988 28902
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16764 25764 16816 25770
rect 16764 25706 16816 25712
rect 16776 25498 16804 25706
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16580 24676 16632 24682
rect 16580 24618 16632 24624
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16500 20942 16528 24006
rect 16592 22030 16620 24618
rect 16580 22024 16632 22030
rect 16868 22001 16896 27338
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17144 24818 17172 25774
rect 17132 24812 17184 24818
rect 17052 24772 17132 24800
rect 17052 23730 17080 24772
rect 17132 24754 17184 24760
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17420 23118 17448 32438
rect 17592 32020 17644 32026
rect 17592 31962 17644 31968
rect 17500 31204 17552 31210
rect 17500 31146 17552 31152
rect 17512 30666 17540 31146
rect 17500 30660 17552 30666
rect 17500 30602 17552 30608
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 16580 21966 16632 21972
rect 16854 21992 16910 22001
rect 16854 21927 16910 21936
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17236 21622 17264 21830
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16960 20534 16988 21286
rect 17328 20874 17356 22374
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21894 17448 21966
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17316 20868 17368 20874
rect 17316 20810 17368 20816
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16960 19446 16988 20470
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16316 18686 16436 18714
rect 16316 18222 16344 18686
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16316 16182 16344 18158
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 16408 11626 16436 18226
rect 16500 17610 16528 19382
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16776 16782 16988 16810
rect 16776 16522 16804 16782
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16868 14482 16896 16594
rect 16960 16522 16988 16782
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17052 16658 17080 16730
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16182 17080 16390
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 14362 16896 14418
rect 16684 14334 16896 14362
rect 16684 11898 16712 14334
rect 16960 14006 16988 15982
rect 17144 14906 17172 20742
rect 17512 19922 17540 28494
rect 17604 22094 17632 31962
rect 17696 28937 17724 36654
rect 17788 36582 17816 37130
rect 18064 37108 18092 39200
rect 19352 37738 19380 39200
rect 19340 37732 19392 37738
rect 19340 37674 19392 37680
rect 18420 37392 18472 37398
rect 18326 37360 18382 37369
rect 18420 37334 18472 37340
rect 18788 37392 18840 37398
rect 18788 37334 18840 37340
rect 19430 37360 19486 37369
rect 18326 37295 18382 37304
rect 18340 37262 18368 37295
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 18432 37194 18460 37334
rect 18420 37188 18472 37194
rect 18420 37130 18472 37136
rect 17880 37080 18092 37108
rect 17880 36786 17908 37080
rect 17868 36780 17920 36786
rect 17868 36722 17920 36728
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 18420 36712 18472 36718
rect 18420 36654 18472 36660
rect 17776 36576 17828 36582
rect 17776 36518 17828 36524
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 17788 35834 17816 36042
rect 17776 35828 17828 35834
rect 17776 35770 17828 35776
rect 17788 35630 17816 35770
rect 18156 35698 18184 36654
rect 18236 36576 18288 36582
rect 18236 36518 18288 36524
rect 18248 36174 18276 36518
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18144 35692 18196 35698
rect 18144 35634 18196 35640
rect 17776 35624 17828 35630
rect 17776 35566 17828 35572
rect 17958 35320 18014 35329
rect 17958 35255 17960 35264
rect 18012 35255 18014 35264
rect 17960 35226 18012 35232
rect 18156 34474 18184 35634
rect 18144 34468 18196 34474
rect 18144 34410 18196 34416
rect 18156 33454 18184 34410
rect 18144 33448 18196 33454
rect 18144 33390 18196 33396
rect 18432 32910 18460 36654
rect 18512 35760 18564 35766
rect 18512 35702 18564 35708
rect 18524 33266 18552 35702
rect 18602 33280 18658 33289
rect 18524 33238 18602 33266
rect 18602 33215 18658 33224
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17880 31142 17908 32506
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17972 30666 18000 32302
rect 18248 31686 18276 32302
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18248 31346 18276 31622
rect 18510 31376 18566 31385
rect 18236 31340 18288 31346
rect 18510 31311 18566 31320
rect 18236 31282 18288 31288
rect 18144 30796 18196 30802
rect 18248 30784 18276 31282
rect 18524 31278 18552 31311
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18196 30756 18276 30784
rect 18144 30738 18196 30744
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 18248 30258 18276 30756
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17776 28960 17828 28966
rect 17682 28928 17738 28937
rect 17776 28902 17828 28908
rect 17866 28928 17922 28937
rect 17682 28863 17738 28872
rect 17788 28558 17816 28902
rect 17866 28863 17922 28872
rect 17880 28762 17908 28863
rect 17972 28801 18000 29174
rect 18156 29102 18184 29582
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 17958 28792 18014 28801
rect 17868 28756 17920 28762
rect 17958 28727 18014 28736
rect 17868 28698 17920 28704
rect 17776 28552 17828 28558
rect 17682 28520 17738 28529
rect 17776 28494 17828 28500
rect 17682 28455 17684 28464
rect 17736 28455 17738 28464
rect 17684 28426 17736 28432
rect 18156 28014 18184 29038
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 26994 18184 27950
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17880 22982 17908 25230
rect 17972 23662 18000 26522
rect 18248 26194 18276 30058
rect 18432 29073 18460 30738
rect 18616 30190 18644 33215
rect 18800 33153 18828 37334
rect 19430 37295 19486 37304
rect 19340 37256 19392 37262
rect 19260 37204 19340 37210
rect 19260 37198 19392 37204
rect 19260 37182 19380 37198
rect 18972 37120 19024 37126
rect 18972 37062 19024 37068
rect 18984 33454 19012 37062
rect 19260 36174 19288 37182
rect 19444 36718 19472 37295
rect 19996 37126 20024 39200
rect 20352 37732 20404 37738
rect 20352 37674 20404 37680
rect 20260 37460 20312 37466
rect 20260 37402 20312 37408
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19996 36910 20208 36938
rect 19996 36802 20024 36910
rect 20180 36854 20208 36910
rect 19536 36774 20024 36802
rect 20076 36848 20128 36854
rect 20076 36790 20128 36796
rect 20168 36848 20220 36854
rect 20168 36790 20220 36796
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19536 36258 19564 36774
rect 19708 36644 19760 36650
rect 19708 36586 19760 36592
rect 19352 36242 19564 36258
rect 19340 36236 19564 36242
rect 19392 36230 19564 36236
rect 19340 36178 19392 36184
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19156 35012 19208 35018
rect 19156 34954 19208 34960
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18972 33448 19024 33454
rect 18972 33390 19024 33396
rect 18786 33144 18842 33153
rect 18786 33079 18842 33088
rect 18892 33017 18920 33390
rect 18878 33008 18934 33017
rect 18878 32943 18934 32952
rect 18696 32360 18748 32366
rect 18696 32302 18748 32308
rect 18708 30802 18736 32302
rect 18892 30938 18920 32943
rect 18972 32768 19024 32774
rect 18972 32710 19024 32716
rect 18984 31414 19012 32710
rect 19062 31920 19118 31929
rect 19062 31855 19118 31864
rect 19076 31754 19104 31855
rect 19064 31748 19116 31754
rect 19064 31690 19116 31696
rect 18972 31408 19024 31414
rect 18972 31350 19024 31356
rect 19168 30938 19196 34954
rect 19260 34490 19288 36110
rect 19616 36100 19668 36106
rect 19720 36088 19748 36586
rect 19668 36060 19748 36088
rect 19616 36042 19668 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19444 34626 19472 35702
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19616 34740 19668 34746
rect 19616 34682 19668 34688
rect 19628 34626 19656 34682
rect 19892 34672 19944 34678
rect 19812 34632 19892 34660
rect 19812 34626 19840 34632
rect 19444 34598 19564 34626
rect 19628 34598 19840 34626
rect 19892 34614 19944 34620
rect 19260 34474 19472 34490
rect 19248 34468 19472 34474
rect 19300 34462 19472 34468
rect 19248 34410 19300 34416
rect 19260 34379 19288 34410
rect 19444 34406 19472 34462
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19352 33833 19380 34342
rect 19338 33824 19394 33833
rect 19338 33759 19394 33768
rect 19352 32570 19380 33759
rect 19444 32978 19472 34342
rect 19536 33998 19564 34598
rect 19616 34468 19668 34474
rect 19996 34456 20024 35430
rect 19668 34428 20024 34456
rect 19616 34410 19668 34416
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19628 33998 19656 34138
rect 19524 33992 19576 33998
rect 19524 33934 19576 33940
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33658 20024 33798
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19800 33584 19852 33590
rect 19800 33526 19852 33532
rect 19812 33402 19840 33526
rect 19720 33386 19840 33402
rect 19708 33380 19840 33386
rect 19760 33374 19840 33380
rect 19890 33416 19946 33425
rect 19890 33351 19892 33360
rect 19708 33322 19760 33328
rect 19944 33351 19946 33360
rect 19892 33322 19944 33328
rect 19432 32972 19484 32978
rect 19432 32914 19484 32920
rect 19432 32836 19484 32842
rect 19432 32778 19484 32784
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19444 32026 19472 32778
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19444 31482 19472 31962
rect 19628 31754 19656 32506
rect 19982 32328 20038 32337
rect 19982 32263 20038 32272
rect 19996 32230 20024 32263
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 19616 31748 19668 31754
rect 19616 31690 19668 31696
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 19156 30932 19208 30938
rect 19156 30874 19208 30880
rect 19996 30802 20024 31078
rect 18696 30796 18748 30802
rect 18696 30738 18748 30744
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19800 30320 19852 30326
rect 19798 30288 19800 30297
rect 19852 30288 19854 30297
rect 19798 30223 19854 30232
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18878 30152 18934 30161
rect 18878 30087 18934 30096
rect 18892 29220 18920 30087
rect 19062 29880 19118 29889
rect 19062 29815 19064 29824
rect 19116 29815 19118 29824
rect 19798 29880 19854 29889
rect 19798 29815 19800 29824
rect 19064 29786 19116 29792
rect 19852 29815 19854 29824
rect 19800 29786 19852 29792
rect 18972 29776 19024 29782
rect 18972 29718 19024 29724
rect 18984 29345 19012 29718
rect 19338 29608 19394 29617
rect 19338 29543 19394 29552
rect 19352 29510 19380 29543
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19430 29472 19486 29481
rect 19430 29407 19486 29416
rect 18970 29336 19026 29345
rect 18970 29271 19026 29280
rect 19246 29336 19302 29345
rect 19246 29271 19302 29280
rect 18892 29192 19196 29220
rect 18418 29064 18474 29073
rect 18418 28999 18474 29008
rect 18972 28960 19024 28966
rect 18972 28902 19024 28908
rect 18156 26166 18276 26194
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17972 22094 18000 23598
rect 17604 22066 17816 22094
rect 17972 22066 18092 22094
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17604 18834 17632 20334
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17512 18426 17540 18634
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17696 17270 17724 17614
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17788 17134 17816 22066
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 19786 17908 21422
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17316 15972 17368 15978
rect 17316 15914 17368 15920
rect 17328 15638 17356 15914
rect 17604 15910 17632 16730
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17052 14878 17172 14906
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 17052 12434 17080 14878
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14346 17172 14758
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 16776 12406 17080 12434
rect 16776 11898 16804 12406
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16408 11150 16436 11562
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 14936 2446 14964 7142
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 2582 16160 2790
rect 16684 2650 16712 11698
rect 16960 11218 16988 12106
rect 17052 11898 17080 12106
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17144 11354 17172 13942
rect 17512 11762 17540 14214
rect 17788 13870 17816 15098
rect 17880 14482 17908 19314
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17972 17542 18000 17818
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17972 15434 18000 17138
rect 18064 15502 18092 22066
rect 18156 20262 18184 26166
rect 18602 24168 18658 24177
rect 18602 24103 18658 24112
rect 18616 23526 18644 24103
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18248 17202 18276 22646
rect 18616 22438 18644 23462
rect 18800 22710 18828 23462
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18340 18970 18368 20470
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18340 18426 18368 18702
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18892 18358 18920 22034
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 18064 15026 18092 15438
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17604 12306 17632 13806
rect 17880 13326 17908 14282
rect 18248 14006 18276 15302
rect 18892 15162 18920 18294
rect 18984 18193 19012 28902
rect 19168 26926 19196 29192
rect 19260 28966 19288 29271
rect 19338 29200 19394 29209
rect 19338 29135 19394 29144
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19156 26920 19208 26926
rect 19156 26862 19208 26868
rect 19352 26518 19380 29135
rect 19444 28098 19472 29407
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20088 29050 20116 36790
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 20180 33454 20208 36178
rect 20272 35698 20300 37402
rect 20364 36718 20392 37674
rect 21284 37262 21312 39200
rect 22572 37262 22600 39200
rect 22928 37324 22980 37330
rect 22928 37266 22980 37272
rect 20812 37256 20864 37262
rect 20812 37198 20864 37204
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 20352 36712 20404 36718
rect 20352 36654 20404 36660
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20456 36378 20484 36654
rect 20720 36644 20772 36650
rect 20720 36586 20772 36592
rect 20732 36378 20760 36586
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20626 36136 20682 36145
rect 20626 36071 20682 36080
rect 20720 36100 20772 36106
rect 20640 36038 20668 36071
rect 20720 36042 20772 36048
rect 20536 36032 20588 36038
rect 20536 35974 20588 35980
rect 20628 36032 20680 36038
rect 20628 35974 20680 35980
rect 20260 35692 20312 35698
rect 20260 35634 20312 35640
rect 20260 34196 20312 34202
rect 20260 34138 20312 34144
rect 20168 33448 20220 33454
rect 20168 33390 20220 33396
rect 20272 33386 20300 34138
rect 20260 33380 20312 33386
rect 20260 33322 20312 33328
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 20260 32496 20312 32502
rect 20260 32438 20312 32444
rect 20350 32464 20406 32473
rect 20166 31784 20222 31793
rect 20166 31719 20168 31728
rect 20220 31719 20222 31728
rect 20168 31690 20220 31696
rect 20168 30184 20220 30190
rect 20166 30152 20168 30161
rect 20220 30152 20222 30161
rect 20166 30087 20222 30096
rect 20166 29744 20222 29753
rect 20166 29679 20222 29688
rect 20180 29578 20208 29679
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 19984 29028 20036 29034
rect 20088 29022 20208 29050
rect 19984 28970 20036 28976
rect 19996 28490 20024 28970
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 20088 28762 20116 28902
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19524 28144 19576 28150
rect 19444 28092 19524 28098
rect 19444 28086 19576 28092
rect 19444 28070 19564 28086
rect 20076 27396 20128 27402
rect 20076 27338 20128 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25838 19380 26318
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19076 24342 19104 25774
rect 19352 25362 19380 25774
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 19352 24886 19380 25298
rect 19444 24936 19472 26862
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19706 25256 19762 25265
rect 19706 25191 19708 25200
rect 19760 25191 19762 25200
rect 19708 25162 19760 25168
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19444 24908 19564 24936
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18970 18184 19026 18193
rect 18970 18119 19026 18128
rect 18984 16726 19012 18119
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 19076 16658 19104 24278
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19260 20874 19288 24074
rect 19352 23866 19380 24822
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24070 19472 24550
rect 19536 24177 19564 24908
rect 19708 24880 19760 24886
rect 19708 24822 19760 24828
rect 19614 24304 19670 24313
rect 19720 24274 19748 24822
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19614 24239 19616 24248
rect 19668 24239 19670 24248
rect 19708 24268 19760 24274
rect 19616 24210 19668 24216
rect 19708 24210 19760 24216
rect 19522 24168 19578 24177
rect 19522 24103 19578 24112
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19352 23186 19380 23802
rect 19444 23798 19472 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22574 19380 23122
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19338 22400 19394 22409
rect 19338 22335 19394 22344
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19168 18970 19196 19382
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19260 18850 19288 20810
rect 19168 18822 19288 18850
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18510 14376 18566 14385
rect 18510 14311 18566 14320
rect 18524 14278 18552 14311
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18616 13530 18644 13806
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17880 12434 17908 13262
rect 18340 12918 18368 13466
rect 19168 12986 19196 18822
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14074 19288 14826
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 17788 12406 17908 12434
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17052 10742 17080 11018
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 9926 16988 10542
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17052 3058 17080 9522
rect 17328 3126 17356 11086
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16776 2446 16804 2790
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 5184 800 5212 2382
rect 6472 800 6500 2382
rect 7116 800 7144 2382
rect 8404 800 8432 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10336 800 10364 2382
rect 11624 800 11652 2382
rect 12912 800 12940 2382
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 2106 13032 2246
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 13556 800 13584 2382
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 14844 800 14872 2246
rect 16132 800 16160 2246
rect 16776 800 16804 2246
rect 17052 2106 17080 2994
rect 17512 2310 17540 11698
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17604 11558 17632 11630
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11218 17632 11494
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17788 2378 17816 12406
rect 19352 9654 19380 22335
rect 19444 21146 19472 23258
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 19904 23118 19932 23190
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19996 23050 20024 24686
rect 20088 23322 20116 27338
rect 20180 25922 20208 29022
rect 20272 26314 20300 32438
rect 20350 32399 20352 32408
rect 20404 32399 20406 32408
rect 20352 32370 20404 32376
rect 20364 29209 20392 32370
rect 20456 32366 20484 32710
rect 20444 32360 20496 32366
rect 20444 32302 20496 32308
rect 20548 31754 20576 35974
rect 20732 35154 20760 36042
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 20824 35086 20852 37198
rect 21008 36786 21036 37198
rect 21180 37120 21232 37126
rect 21180 37062 21232 37068
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 22100 37120 22152 37126
rect 22100 37062 22152 37068
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21192 36553 21220 37062
rect 22020 36922 22048 37062
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 22112 36802 22140 37062
rect 21928 36774 22140 36802
rect 22744 36780 22796 36786
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 20902 36544 20958 36553
rect 20902 36479 20958 36488
rect 21178 36544 21234 36553
rect 21178 36479 21234 36488
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20628 35012 20680 35018
rect 20628 34954 20680 34960
rect 20456 31726 20576 31754
rect 20350 29200 20406 29209
rect 20350 29135 20406 29144
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20364 28626 20392 28698
rect 20352 28620 20404 28626
rect 20352 28562 20404 28568
rect 20456 28558 20484 31726
rect 20536 31408 20588 31414
rect 20640 31396 20668 34954
rect 20720 34536 20772 34542
rect 20916 34524 20944 36479
rect 21180 36032 21232 36038
rect 21180 35974 21232 35980
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 20772 34496 20944 34524
rect 20720 34478 20772 34484
rect 20718 33960 20774 33969
rect 20718 33895 20774 33904
rect 20732 32842 20760 33895
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20588 31368 20668 31396
rect 20536 31350 20588 31356
rect 20548 29238 20576 31350
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20536 29232 20588 29238
rect 20536 29174 20588 29180
rect 20640 29084 20668 29990
rect 20718 29608 20774 29617
rect 20718 29543 20774 29552
rect 20732 29102 20760 29543
rect 20548 29056 20668 29084
rect 20720 29096 20772 29102
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20456 28150 20484 28494
rect 20444 28144 20496 28150
rect 20444 28086 20496 28092
rect 20260 26308 20312 26314
rect 20312 26268 20484 26296
rect 20260 26250 20312 26256
rect 20180 25894 20300 25922
rect 20168 25832 20220 25838
rect 20168 25774 20220 25780
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19444 20806 19472 21082
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19444 19310 19472 19926
rect 19628 19786 19656 20198
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19304 19484 19310
rect 19484 19264 19564 19292
rect 19432 19246 19484 19252
rect 19536 18834 19564 19264
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 18086 19472 18226
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17678 19472 18022
rect 19996 17746 20024 22986
rect 20074 22808 20130 22817
rect 20074 22743 20076 22752
rect 20128 22743 20130 22752
rect 20076 22714 20128 22720
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20088 19990 20116 20198
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 20088 19174 20116 19654
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 15502 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16250 20024 16594
rect 20088 16454 20116 18906
rect 20180 18698 20208 25774
rect 20272 22817 20300 25894
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20258 22808 20314 22817
rect 20258 22743 20314 22752
rect 20364 22692 20392 24074
rect 20272 22664 20392 22692
rect 20272 22506 20300 22664
rect 20456 22624 20484 26268
rect 20548 25158 20576 29056
rect 20720 29038 20772 29044
rect 20732 28626 20760 29038
rect 20824 28762 20852 33050
rect 21008 31929 21036 35430
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21100 34202 21128 34342
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 20994 31920 21050 31929
rect 20994 31855 21050 31864
rect 21008 31754 21036 31855
rect 21008 31726 21128 31754
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 31278 21036 31622
rect 21100 31346 21128 31726
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 20996 31272 21048 31278
rect 20996 31214 21048 31220
rect 21192 31226 21220 35974
rect 21272 35216 21324 35222
rect 21272 35158 21324 35164
rect 21284 34678 21312 35158
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21376 33114 21404 36654
rect 21928 36106 21956 36774
rect 22744 36722 22796 36728
rect 22756 36553 22784 36722
rect 22742 36544 22798 36553
rect 22742 36479 22798 36488
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21456 34740 21508 34746
rect 21456 34682 21508 34688
rect 21548 34740 21600 34746
rect 21548 34682 21600 34688
rect 21468 33930 21496 34682
rect 21560 34134 21588 34682
rect 21548 34128 21600 34134
rect 21548 34070 21600 34076
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21272 32292 21324 32298
rect 21272 32234 21324 32240
rect 21284 31754 21312 32234
rect 21928 32230 21956 36042
rect 22008 35012 22060 35018
rect 22008 34954 22060 34960
rect 22020 34542 22048 34954
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 22284 34536 22336 34542
rect 22284 34478 22336 34484
rect 22020 33998 22048 34478
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22296 32434 22324 34478
rect 22284 32428 22336 32434
rect 22284 32370 22336 32376
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 22572 31754 22600 34886
rect 22940 33114 22968 37266
rect 23216 37262 23244 39200
rect 24504 39114 24532 39200
rect 24596 39114 24624 39222
rect 24504 39086 24624 39114
rect 24780 37346 24808 39222
rect 25778 39200 25834 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 24780 37318 24900 37346
rect 25792 37330 25820 39200
rect 26330 37360 26386 37369
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 23940 36712 23992 36718
rect 23940 36654 23992 36660
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23572 36576 23624 36582
rect 23572 36518 23624 36524
rect 23308 36106 23336 36518
rect 23584 36242 23612 36518
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 23296 36100 23348 36106
rect 23296 36042 23348 36048
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 23018 35456 23074 35465
rect 23018 35391 23074 35400
rect 23032 33930 23060 35391
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22744 32972 22796 32978
rect 22744 32914 22796 32920
rect 22652 32836 22704 32842
rect 22652 32778 22704 32784
rect 22664 32570 22692 32778
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22756 32434 22784 32914
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 21284 31726 21496 31754
rect 21008 30802 21036 31214
rect 21192 31198 21312 31226
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 21284 30666 21312 31198
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21284 30394 21312 30602
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 20732 28082 20760 28562
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22778 20576 22918
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20640 22624 20668 27270
rect 20916 25498 20944 29718
rect 21192 29186 21220 30262
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 21284 29306 21312 29446
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 21192 29158 21312 29186
rect 20996 29028 21048 29034
rect 20996 28970 21048 28976
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 21008 28762 21036 28970
rect 20996 28756 21048 28762
rect 20996 28698 21048 28704
rect 20996 28484 21048 28490
rect 20996 28426 21048 28432
rect 21008 26926 21036 28426
rect 21100 28014 21128 28970
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21284 26382 21312 29158
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20994 25392 21050 25401
rect 20732 23186 20760 25366
rect 20994 25327 21050 25336
rect 21008 25226 21036 25327
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20824 24274 20852 24618
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21008 23798 21036 24006
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20732 23066 20760 23122
rect 20732 23038 20852 23066
rect 20364 22596 20484 22624
rect 20548 22596 20668 22624
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20180 17338 20208 18294
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19984 16244 20036 16250
rect 20036 16204 20116 16232
rect 19984 16186 20036 16192
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 15706 19840 16050
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19996 15638 20024 15846
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19444 14346 19472 15098
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13530 19472 13806
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19628 13326 19656 13670
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12238 20024 15098
rect 20088 15026 20116 16204
rect 20180 15094 20208 17002
rect 20272 15094 20300 22442
rect 20364 21554 20392 22596
rect 20548 22012 20576 22596
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20456 21984 20576 22012
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 18970 20392 20742
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20364 16114 20392 18634
rect 20456 18086 20484 21984
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20548 20942 20576 21626
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20626 19952 20682 19961
rect 20626 19887 20682 19896
rect 20640 19854 20668 19887
rect 20732 19854 20760 22374
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20640 17354 20668 19790
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19446 20760 19654
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 18358 20760 18770
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20456 17326 20668 17354
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20180 13394 20208 15030
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20088 12442 20116 12854
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19628 11082 19656 11562
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19352 9042 19380 9590
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 3126 17908 3402
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18064 2446 18092 8570
rect 18800 7410 18828 8774
rect 19444 8498 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 8974 19932 9318
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20180 2650 20208 12786
rect 20456 12434 20484 17326
rect 20732 16522 20760 17546
rect 20824 17202 20852 23038
rect 20902 21992 20958 22001
rect 20902 21927 20958 21936
rect 20916 21690 20944 21927
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 21008 20602 21036 23734
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 21008 17202 21036 20538
rect 21100 19378 21128 24006
rect 21192 21350 21220 25910
rect 21284 22506 21312 26318
rect 21468 25226 21496 31726
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22560 31748 22612 31754
rect 22560 31690 22612 31696
rect 21640 31204 21692 31210
rect 21640 31146 21692 31152
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21284 21010 21312 22442
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21270 20632 21326 20641
rect 21270 20567 21326 20576
rect 21284 19378 21312 20567
rect 21376 19514 21404 22578
rect 21468 22166 21496 23462
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21376 17338 21404 17546
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20810 16824 20866 16833
rect 20810 16759 20866 16768
rect 20824 16726 20852 16759
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20548 16046 20576 16458
rect 20626 16144 20682 16153
rect 20626 16079 20682 16088
rect 20720 16108 20772 16114
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20364 12406 20484 12434
rect 20364 7954 20392 12406
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 9178 20484 9454
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20548 2582 20576 15982
rect 20640 15910 20668 16079
rect 20720 16050 20772 16056
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 14074 20668 15030
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20640 11762 20668 14010
rect 20732 14006 20760 16050
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15026 20852 15846
rect 21468 15502 21496 19450
rect 21560 16590 21588 29106
rect 21652 23662 21680 31146
rect 22112 29714 22140 31690
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 21732 28620 21784 28626
rect 21732 28562 21784 28568
rect 21744 28422 21772 28562
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 21732 26036 21784 26042
rect 21732 25978 21784 25984
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21744 22030 21772 25978
rect 22112 25906 22140 29174
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22204 25294 22232 26182
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22296 25362 22324 25774
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 21836 24070 21864 25162
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22112 24410 22140 24550
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21836 20398 21864 23598
rect 21928 21146 21956 24006
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 22020 21486 22048 22646
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 22204 20942 22232 25094
rect 22388 24954 22416 26862
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22480 24834 22508 31282
rect 23492 31278 23520 35974
rect 23848 35488 23900 35494
rect 23848 35430 23900 35436
rect 23860 35290 23888 35430
rect 23848 35284 23900 35290
rect 23848 35226 23900 35232
rect 23952 34542 23980 36654
rect 24780 36582 24808 37198
rect 24872 36786 24900 37318
rect 25504 37324 25556 37330
rect 25504 37266 25556 37272
rect 25780 37324 25832 37330
rect 26330 37295 26386 37304
rect 25780 37266 25832 37272
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24858 36544 24914 36553
rect 24780 36106 24808 36518
rect 24858 36479 24914 36488
rect 24872 36122 24900 36479
rect 24872 36106 25084 36122
rect 24768 36100 24820 36106
rect 24768 36042 24820 36048
rect 24860 36100 25084 36106
rect 24912 36094 25084 36100
rect 24860 36042 24912 36048
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24308 35148 24360 35154
rect 24308 35090 24360 35096
rect 24320 34610 24348 35090
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24688 34542 24716 35634
rect 24780 35630 24808 36042
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24780 35154 24808 35566
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24872 35222 24900 35430
rect 24860 35216 24912 35222
rect 24860 35158 24912 35164
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24964 35018 24992 35974
rect 24952 35012 25004 35018
rect 24952 34954 25004 34960
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23940 34536 23992 34542
rect 23940 34478 23992 34484
rect 24676 34536 24728 34542
rect 24676 34478 24728 34484
rect 23768 32910 23796 34478
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 24688 33658 24716 33866
rect 24768 33856 24820 33862
rect 24768 33798 24820 33804
rect 24860 33856 24912 33862
rect 24860 33798 24912 33804
rect 24780 33658 24808 33798
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24872 33590 24900 33798
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24400 33448 24452 33454
rect 24400 33390 24452 33396
rect 24412 32910 24440 33390
rect 24492 33040 24544 33046
rect 24492 32982 24544 32988
rect 23756 32904 23808 32910
rect 23756 32846 23808 32852
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 23940 32768 23992 32774
rect 23940 32710 23992 32716
rect 23952 32502 23980 32710
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 23940 32496 23992 32502
rect 23940 32438 23992 32444
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23664 32292 23716 32298
rect 23664 32234 23716 32240
rect 23676 32026 23704 32234
rect 23768 32230 23796 32370
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23768 31958 23796 32166
rect 24136 31958 24164 32506
rect 24320 32502 24348 32778
rect 24308 32496 24360 32502
rect 24308 32438 24360 32444
rect 24412 32230 24440 32846
rect 24504 32502 24532 32982
rect 24582 32872 24638 32881
rect 24582 32807 24638 32816
rect 24492 32496 24544 32502
rect 24492 32438 24544 32444
rect 24596 32230 24624 32807
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24584 32224 24636 32230
rect 24584 32166 24636 32172
rect 24412 32008 24440 32166
rect 24584 32020 24636 32026
rect 24412 31980 24584 32008
rect 23756 31952 23808 31958
rect 23756 31894 23808 31900
rect 24124 31952 24176 31958
rect 24124 31894 24176 31900
rect 24308 31952 24360 31958
rect 24308 31894 24360 31900
rect 23480 31272 23532 31278
rect 23480 31214 23532 31220
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22572 28490 22600 29038
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22388 24806 22508 24834
rect 22296 24410 22324 24754
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 22388 20330 22416 24806
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22480 21690 22508 23666
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22572 20466 22600 28426
rect 22664 25158 22692 31078
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22940 29578 22968 30602
rect 23388 30320 23440 30326
rect 23388 30262 23440 30268
rect 22928 29572 22980 29578
rect 22928 29514 22980 29520
rect 22940 29170 22968 29514
rect 23296 29232 23348 29238
rect 23296 29174 23348 29180
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 23020 29096 23072 29102
rect 23020 29038 23072 29044
rect 23032 28558 23060 29038
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 22836 27940 22888 27946
rect 22836 27882 22888 27888
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22848 23322 22876 27882
rect 23032 27130 23060 28494
rect 23308 27402 23336 29174
rect 23400 27606 23428 30262
rect 23492 30258 23520 31214
rect 24320 30666 24348 31894
rect 24308 30660 24360 30666
rect 24308 30602 24360 30608
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 24216 30252 24268 30258
rect 24412 30240 24440 31980
rect 24584 31962 24636 31968
rect 24596 31890 24624 31962
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 24964 31770 24992 31826
rect 24688 31742 24992 31770
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24596 30433 24624 31282
rect 24582 30424 24638 30433
rect 24582 30359 24638 30368
rect 24268 30212 24440 30240
rect 24216 30194 24268 30200
rect 24216 30116 24268 30122
rect 24216 30058 24268 30064
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 24228 30002 24256 30058
rect 24688 30054 24716 31742
rect 25056 30297 25084 36094
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25148 34134 25176 35566
rect 25136 34128 25188 34134
rect 25136 34070 25188 34076
rect 25136 33924 25188 33930
rect 25136 33866 25188 33872
rect 25148 33590 25176 33866
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 25332 33402 25360 36042
rect 25148 33374 25360 33402
rect 25042 30288 25098 30297
rect 25042 30223 25098 30232
rect 24676 30048 24728 30054
rect 23572 29776 23624 29782
rect 23572 29718 23624 29724
rect 23584 29510 23612 29718
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23848 29232 23900 29238
rect 23848 29174 23900 29180
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 23308 26926 23336 27338
rect 23664 27056 23716 27062
rect 23664 26998 23716 27004
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23020 26444 23072 26450
rect 23020 26386 23072 26392
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22848 21962 22876 23258
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22742 21856 22798 21865
rect 22742 21791 22798 21800
rect 22650 20904 22706 20913
rect 22650 20839 22652 20848
rect 22704 20839 22706 20848
rect 22652 20810 22704 20816
rect 22664 20466 22692 20810
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 21730 20088 21786 20097
rect 21730 20023 21732 20032
rect 21784 20023 21786 20032
rect 21824 20052 21876 20058
rect 21732 19994 21784 20000
rect 21824 19994 21876 20000
rect 21836 19854 21864 19994
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 22112 19310 22140 20266
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22756 17898 22784 21791
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22848 20330 22876 20402
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22940 20058 22968 20742
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 23032 19922 23060 26386
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23124 20874 23152 21354
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23216 20058 23244 24822
rect 23480 24744 23532 24750
rect 23400 24704 23480 24732
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23308 21622 23336 24074
rect 23400 23866 23428 24704
rect 23480 24686 23532 24692
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23400 23730 23428 23802
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 23388 21140 23440 21146
rect 23492 21128 23520 22986
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23584 21418 23612 22510
rect 23572 21412 23624 21418
rect 23572 21354 23624 21360
rect 23440 21100 23520 21128
rect 23388 21082 23440 21088
rect 23676 20992 23704 26998
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23322 23796 23462
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23676 20964 23796 20992
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23676 20602 23704 20810
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 22756 17870 22968 17898
rect 22940 17746 22968 17870
rect 23308 17785 23336 20334
rect 23584 19854 23612 20334
rect 23768 20058 23796 20964
rect 23860 20602 23888 29174
rect 23952 28218 23980 29990
rect 24228 29974 24532 30002
rect 24676 29990 24728 29996
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 24504 29866 24532 29974
rect 24872 29866 24900 29990
rect 24504 29838 24900 29866
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29186 24532 29582
rect 24504 29170 24624 29186
rect 24504 29164 24636 29170
rect 24504 29158 24584 29164
rect 24584 29106 24636 29112
rect 24872 29102 24900 29650
rect 25148 29510 25176 33374
rect 25424 33266 25452 36654
rect 25240 33238 25452 33266
rect 25240 31482 25268 33238
rect 25516 32994 25544 37266
rect 26240 37256 26292 37262
rect 25870 37224 25926 37233
rect 26240 37198 26292 37204
rect 25870 37159 25926 37168
rect 25884 36922 25912 37159
rect 25872 36916 25924 36922
rect 25872 36858 25924 36864
rect 26252 36650 26280 37198
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 26240 36644 26292 36650
rect 26240 36586 26292 36592
rect 26160 36106 26188 36586
rect 26344 36310 26372 37295
rect 26436 37194 26464 39200
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 26424 37188 26476 37194
rect 26424 37130 26476 37136
rect 26424 36576 26476 36582
rect 26424 36518 26476 36524
rect 26436 36378 26464 36518
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26332 36304 26384 36310
rect 26332 36246 26384 36252
rect 26148 36100 26200 36106
rect 26148 36042 26200 36048
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 25596 33584 25648 33590
rect 25594 33552 25596 33561
rect 25648 33552 25650 33561
rect 25594 33487 25650 33496
rect 25516 32966 25636 32994
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25516 32337 25544 32778
rect 25502 32328 25558 32337
rect 25502 32263 25558 32272
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 31754 25360 32166
rect 25320 31748 25372 31754
rect 25320 31690 25372 31696
rect 25504 31680 25556 31686
rect 25504 31622 25556 31628
rect 25228 31476 25280 31482
rect 25228 31418 25280 31424
rect 25516 31278 25544 31622
rect 25412 31272 25464 31278
rect 25412 31214 25464 31220
rect 25504 31272 25556 31278
rect 25504 31214 25556 31220
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24872 28626 24900 29038
rect 24952 29028 25004 29034
rect 25240 28994 25268 31078
rect 25424 30802 25452 31214
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25516 30682 25544 31214
rect 24952 28970 25004 28976
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24964 28506 24992 28970
rect 24872 28478 24992 28506
rect 25148 28966 25268 28994
rect 25424 30654 25544 30682
rect 23940 28212 23992 28218
rect 23940 28154 23992 28160
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24044 25770 24072 28154
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24412 26790 24440 27474
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24596 27130 24624 27406
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24596 26450 24624 27066
rect 24872 26586 24900 28478
rect 24952 27872 25004 27878
rect 24952 27814 25004 27820
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 24032 25764 24084 25770
rect 24032 25706 24084 25712
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23952 21078 23980 21830
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18834 23980 19110
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23570 18320 23626 18329
rect 23570 18255 23626 18264
rect 23584 18222 23612 18255
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23294 17776 23350 17785
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22928 17740 22980 17746
rect 23294 17711 23350 17720
rect 22928 17682 22980 17688
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21652 17066 21680 17546
rect 22480 17270 22508 17614
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 15502 21588 16526
rect 22296 16454 22324 17138
rect 22572 16590 22600 17478
rect 22756 16794 22784 17546
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22652 16176 22704 16182
rect 22650 16144 22652 16153
rect 22704 16144 22706 16153
rect 22650 16079 22706 16088
rect 22652 16040 22704 16046
rect 22650 16008 22652 16017
rect 22704 16008 22706 16017
rect 22650 15943 22706 15952
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20732 13530 20760 13806
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20916 13394 20944 13670
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 21008 11898 21036 13466
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20824 11218 20852 11630
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20916 10810 20944 11630
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21008 10674 21036 10950
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20824 9586 20852 9862
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 21192 2514 21220 15302
rect 21468 14414 21496 15438
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21560 13938 21588 15438
rect 22848 14958 22876 17682
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 14006 22600 14214
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21560 11150 21588 13874
rect 22572 12306 22600 13942
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22848 12102 22876 14894
rect 23400 14090 23428 15370
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23400 14062 23520 14090
rect 23492 14006 23520 14062
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23676 13870 23704 14282
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 24044 13326 24072 25094
rect 24412 24886 24440 25842
rect 24964 25226 24992 27814
rect 25056 27402 25084 27814
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 25148 27062 25176 28966
rect 25320 28484 25372 28490
rect 25320 28426 25372 28432
rect 25332 27674 25360 28426
rect 25320 27668 25372 27674
rect 25320 27610 25372 27616
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24136 22438 24164 22714
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12306 22968 13126
rect 23492 12850 23520 13262
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22112 9654 22140 9998
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22388 9382 22416 9862
rect 22756 9450 22784 11630
rect 22848 11354 22876 11630
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 23032 11150 23060 12582
rect 24136 12434 24164 20810
rect 24228 15162 24256 23258
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 24320 21554 24348 21830
rect 24412 21690 24440 24346
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24596 20602 24624 25162
rect 24858 24304 24914 24313
rect 24858 24239 24860 24248
rect 24912 24239 24914 24248
rect 24860 24210 24912 24216
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24688 20874 24716 24074
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 21962 24808 23054
rect 24872 22710 24900 24210
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24872 20874 24900 21490
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 24872 20466 24900 20810
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24872 19854 24900 20402
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24766 18864 24822 18873
rect 24766 18799 24822 18808
rect 24780 18766 24808 18799
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24872 18358 24900 19790
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24964 15706 24992 25162
rect 25148 23662 25176 26998
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25228 25356 25280 25362
rect 25228 25298 25280 25304
rect 25240 24750 25268 25298
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25240 23866 25268 24686
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25240 23118 25268 23802
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25056 21146 25084 22918
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25148 21690 25176 22102
rect 25226 21992 25282 22001
rect 25226 21927 25282 21936
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 25042 21040 25098 21049
rect 25042 20975 25098 20984
rect 25056 17746 25084 20975
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25148 18766 25176 18906
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25056 17338 25084 17682
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 23952 12406 24164 12434
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11558 23152 12038
rect 23952 11898 23980 12406
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23124 10130 23152 11494
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 22744 9444 22796 9450
rect 22744 9386 22796 9392
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 18064 800 18092 2246
rect 19352 800 19380 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2382
rect 21284 800 21312 2382
rect 22572 800 22600 2382
rect 23124 2378 23152 2586
rect 23492 2582 23520 9522
rect 23860 2650 23888 11698
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24688 10130 24716 10542
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24780 9994 24808 10406
rect 24872 10198 24900 13398
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24964 12374 24992 13126
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24964 11082 24992 12310
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24964 10130 24992 11018
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24596 2650 24624 9862
rect 25056 7886 25084 15302
rect 25148 13258 25176 18022
rect 25240 17202 25268 21927
rect 25332 17542 25360 26522
rect 25424 22094 25452 30654
rect 25608 29714 25636 32966
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25792 32065 25820 32302
rect 25778 32056 25834 32065
rect 25778 31991 25834 32000
rect 25596 29708 25648 29714
rect 25596 29650 25648 29656
rect 25608 29034 25636 29650
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26056 28144 26108 28150
rect 26056 28086 26108 28092
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 25596 26444 25648 26450
rect 25596 26386 25648 26392
rect 25608 23594 25636 26386
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25516 22234 25544 22986
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25424 22066 25544 22094
rect 25412 21072 25464 21078
rect 25412 21014 25464 21020
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25424 17202 25452 21014
rect 25516 19378 25544 22066
rect 25608 21554 25636 22714
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25700 19174 25728 27338
rect 25872 26920 25924 26926
rect 25872 26862 25924 26868
rect 25884 26518 25912 26862
rect 25872 26512 25924 26518
rect 25872 26454 25924 26460
rect 25872 25220 25924 25226
rect 25872 25162 25924 25168
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25792 20913 25820 22578
rect 25884 22094 25912 25162
rect 25884 22066 26004 22094
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25884 21690 25912 21830
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25872 20936 25924 20942
rect 25778 20904 25834 20913
rect 25872 20878 25924 20884
rect 25778 20839 25834 20848
rect 25884 20618 25912 20878
rect 25792 20590 25912 20618
rect 25792 19378 25820 20590
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25792 18986 25820 19314
rect 25700 18958 25820 18986
rect 25700 18698 25728 18958
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25240 16969 25268 17138
rect 25424 16998 25452 17138
rect 25412 16992 25464 16998
rect 25226 16960 25282 16969
rect 25412 16934 25464 16940
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25226 16895 25282 16904
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 14074 25268 14282
rect 25516 14278 25544 16594
rect 25608 16522 25636 16934
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 25688 14544 25740 14550
rect 25688 14486 25740 14492
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25700 14006 25728 14486
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25332 11694 25360 13942
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25148 8634 25176 11630
rect 25332 10742 25360 11630
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25424 9654 25452 11018
rect 25884 10266 25912 20334
rect 25976 20058 26004 22066
rect 26068 20516 26096 28086
rect 26160 22778 26188 28562
rect 26252 27946 26280 34954
rect 26528 34474 26556 35430
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 26608 35012 26660 35018
rect 26608 34954 26660 34960
rect 26516 34468 26568 34474
rect 26516 34410 26568 34416
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26436 33318 26464 34342
rect 26528 33454 26556 34410
rect 26620 34066 26648 34954
rect 26700 34944 26752 34950
rect 26700 34886 26752 34892
rect 26712 34202 26740 34886
rect 26700 34196 26752 34202
rect 26700 34138 26752 34144
rect 26608 34060 26660 34066
rect 26608 34002 26660 34008
rect 26516 33448 26568 33454
rect 26516 33390 26568 33396
rect 26424 33312 26476 33318
rect 26424 33254 26476 33260
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26620 32978 26648 33254
rect 26608 32972 26660 32978
rect 26608 32914 26660 32920
rect 26804 31754 26832 35022
rect 26792 31748 26844 31754
rect 26792 31690 26844 31696
rect 26332 30864 26384 30870
rect 26332 30806 26384 30812
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 26344 27606 26372 30806
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 26516 27056 26568 27062
rect 26516 26998 26568 27004
rect 26332 26920 26384 26926
rect 26332 26862 26384 26868
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26160 21146 26188 22714
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26148 20528 26200 20534
rect 26068 20488 26148 20516
rect 26148 20470 26200 20476
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26252 19514 26280 26250
rect 26344 25158 26372 26862
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26332 25152 26384 25158
rect 26332 25094 26384 25100
rect 26332 23656 26384 23662
rect 26332 23598 26384 23604
rect 26344 22001 26372 23598
rect 26436 22982 26464 26250
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26330 21992 26386 22001
rect 26330 21927 26386 21936
rect 26424 21344 26476 21350
rect 26424 21286 26476 21292
rect 26436 21146 26464 21286
rect 26424 21140 26476 21146
rect 26424 21082 26476 21088
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26344 20466 26372 20878
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26344 19854 26372 20402
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 25964 19440 26016 19446
rect 26016 19388 26280 19394
rect 25964 19382 26280 19388
rect 25976 19378 26280 19382
rect 25976 19372 26292 19378
rect 25976 19366 26240 19372
rect 26240 19314 26292 19320
rect 26054 18864 26110 18873
rect 26344 18834 26372 19790
rect 26436 19378 26464 20470
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26054 18799 26110 18808
rect 26332 18828 26384 18834
rect 26068 13326 26096 18799
rect 26332 18770 26384 18776
rect 26528 18426 26556 26998
rect 26620 22574 26648 29514
rect 26804 29306 26832 31690
rect 26884 29844 26936 29850
rect 26884 29786 26936 29792
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26896 29102 26924 29786
rect 26884 29096 26936 29102
rect 26884 29038 26936 29044
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26896 28762 26924 28902
rect 26884 28756 26936 28762
rect 26884 28698 26936 28704
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26712 26790 26740 28562
rect 26976 27872 27028 27878
rect 26976 27814 27028 27820
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26712 24614 26740 26726
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26896 25430 26924 26182
rect 26884 25424 26936 25430
rect 26884 25366 26936 25372
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26988 23866 27016 27814
rect 27080 26858 27108 37198
rect 27724 37194 27752 39200
rect 27896 37664 27948 37670
rect 27896 37606 27948 37612
rect 27712 37188 27764 37194
rect 27712 37130 27764 37136
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 27632 36378 27660 37062
rect 27908 36938 27936 37606
rect 29012 37194 29040 39200
rect 29656 37330 29684 39200
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 30012 37256 30064 37262
rect 30012 37198 30064 37204
rect 29000 37188 29052 37194
rect 29000 37130 29052 37136
rect 27908 36910 28396 36938
rect 27908 36718 27936 36910
rect 27988 36848 28040 36854
rect 27988 36790 28040 36796
rect 28000 36718 28028 36790
rect 27896 36712 27948 36718
rect 27896 36654 27948 36660
rect 27988 36712 28040 36718
rect 27988 36654 28040 36660
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 27896 36576 27948 36582
rect 27896 36518 27948 36524
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 27528 35828 27580 35834
rect 27528 35770 27580 35776
rect 27436 35624 27488 35630
rect 27434 35592 27436 35601
rect 27488 35592 27490 35601
rect 27434 35527 27490 35536
rect 27448 34950 27476 35527
rect 27540 35494 27568 35770
rect 27632 35698 27660 36314
rect 27724 36242 27752 36518
rect 27712 36236 27764 36242
rect 27712 36178 27764 36184
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27724 35630 27752 36178
rect 27804 36100 27856 36106
rect 27804 36042 27856 36048
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27436 34944 27488 34950
rect 27436 34886 27488 34892
rect 27160 33924 27212 33930
rect 27620 33924 27672 33930
rect 27212 33884 27292 33912
rect 27160 33866 27212 33872
rect 27264 30802 27292 33884
rect 27620 33866 27672 33872
rect 27632 33289 27660 33866
rect 27618 33280 27674 33289
rect 27618 33215 27674 33224
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27356 32026 27384 32166
rect 27344 32020 27396 32026
rect 27344 31962 27396 31968
rect 27436 31408 27488 31414
rect 27436 31350 27488 31356
rect 27252 30796 27304 30802
rect 27252 30738 27304 30744
rect 27448 30734 27476 31350
rect 27816 31249 27844 36042
rect 27908 36038 27936 36518
rect 28368 36106 28396 36910
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 28448 36304 28500 36310
rect 28448 36246 28500 36252
rect 28356 36100 28408 36106
rect 28276 36060 28356 36088
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27988 35624 28040 35630
rect 27988 35566 28040 35572
rect 28000 34746 28028 35566
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27802 31240 27858 31249
rect 27802 31175 27858 31184
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 30546 27476 30670
rect 27804 30660 27856 30666
rect 27804 30602 27856 30608
rect 27448 30518 27568 30546
rect 27540 30326 27568 30518
rect 27528 30320 27580 30326
rect 27528 30262 27580 30268
rect 27540 30190 27568 30262
rect 27528 30184 27580 30190
rect 27528 30126 27580 30132
rect 27436 29504 27488 29510
rect 27436 29446 27488 29452
rect 27068 26852 27120 26858
rect 27068 26794 27120 26800
rect 27448 24750 27476 29446
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27632 28014 27660 28494
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27632 27538 27660 27950
rect 27712 27668 27764 27674
rect 27712 27610 27764 27616
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 27632 27130 27660 27474
rect 27724 27402 27752 27610
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27172 24614 27200 24686
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26608 22568 26660 22574
rect 26608 22510 26660 22516
rect 26804 22234 26832 22918
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26608 22092 26660 22098
rect 26608 22034 26660 22040
rect 26620 20942 26648 22034
rect 26608 20936 26660 20942
rect 26608 20878 26660 20884
rect 26698 20904 26754 20913
rect 26698 20839 26754 20848
rect 26606 20632 26662 20641
rect 26606 20567 26662 20576
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26436 18306 26464 18362
rect 26620 18306 26648 20567
rect 26712 19786 26740 20839
rect 26700 19780 26752 19786
rect 26700 19722 26752 19728
rect 26712 19553 26740 19722
rect 26698 19544 26754 19553
rect 26698 19479 26754 19488
rect 26436 18278 26648 18306
rect 26620 17678 26648 18278
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26148 16720 26200 16726
rect 26148 16662 26200 16668
rect 26160 13870 26188 16662
rect 26804 16658 26832 22170
rect 26884 18692 26936 18698
rect 26884 18634 26936 18640
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26516 16516 26568 16522
rect 26516 16458 26568 16464
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26344 14006 26372 15846
rect 26528 15638 26556 16458
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26514 15328 26570 15337
rect 26514 15263 26570 15272
rect 26528 15162 26556 15263
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26160 13462 26188 13806
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26436 12986 26464 13262
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26804 12434 26832 16594
rect 26896 14958 26924 18634
rect 26988 18290 27016 23802
rect 27172 23730 27200 24550
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27172 22642 27200 23666
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27448 22094 27476 24686
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 27632 23497 27660 23530
rect 27618 23488 27674 23497
rect 27618 23423 27674 23432
rect 27632 23254 27660 23423
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 27528 23044 27580 23050
rect 27528 22986 27580 22992
rect 27264 22066 27476 22094
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27080 20942 27108 21490
rect 27068 20936 27120 20942
rect 27066 20904 27068 20913
rect 27120 20904 27122 20913
rect 27066 20839 27122 20848
rect 27158 20088 27214 20097
rect 27158 20023 27214 20032
rect 27172 19922 27200 20023
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27172 18834 27200 19314
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27080 18358 27108 18702
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27080 17882 27108 18158
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26988 16794 27016 17546
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 27080 17105 27108 17274
rect 27066 17096 27122 17105
rect 27066 17031 27122 17040
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 27080 16538 27108 17031
rect 27172 16658 27200 17682
rect 27264 17490 27292 22066
rect 27436 21956 27488 21962
rect 27436 21898 27488 21904
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27356 19242 27384 21014
rect 27344 19236 27396 19242
rect 27344 19178 27396 19184
rect 27448 18970 27476 21898
rect 27540 20058 27568 22986
rect 27618 21584 27674 21593
rect 27618 21519 27674 21528
rect 27632 21418 27660 21519
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27632 20398 27660 21354
rect 27724 20777 27752 27338
rect 27710 20768 27766 20777
rect 27710 20703 27766 20712
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27528 19236 27580 19242
rect 27528 19178 27580 19184
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 27356 18850 27384 18906
rect 27540 18850 27568 19178
rect 27356 18822 27568 18850
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27356 18358 27384 18566
rect 27344 18352 27396 18358
rect 27344 18294 27396 18300
rect 27264 17462 27384 17490
rect 27250 17368 27306 17377
rect 27250 17303 27252 17312
rect 27304 17303 27306 17312
rect 27252 17274 27304 17280
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27080 16510 27200 16538
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26976 14884 27028 14890
rect 26976 14826 27028 14832
rect 26988 14482 27016 14826
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 13462 27108 14282
rect 27068 13456 27120 13462
rect 27068 13398 27120 13404
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 26712 12406 26832 12434
rect 26712 11762 26740 12406
rect 26896 12170 26924 13126
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26252 10674 26280 11698
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 27172 9586 27200 16510
rect 27264 15638 27292 17002
rect 27252 15632 27304 15638
rect 27252 15574 27304 15580
rect 27356 15450 27384 17462
rect 27448 17202 27476 18702
rect 27526 18320 27582 18329
rect 27526 18255 27582 18264
rect 27540 18222 27568 18255
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27356 15422 27476 15450
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27356 15094 27384 15302
rect 27344 15088 27396 15094
rect 27344 15030 27396 15036
rect 27252 14952 27304 14958
rect 27252 14894 27304 14900
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 23216 800 23244 2382
rect 24504 800 24532 2382
rect 25148 2310 25176 8434
rect 27264 8362 27292 14894
rect 27448 14346 27476 15422
rect 27632 15366 27660 16390
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27632 14958 27660 15302
rect 27620 14952 27672 14958
rect 27620 14894 27672 14900
rect 27816 14618 27844 30602
rect 28092 30054 28120 35974
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 28080 29504 28132 29510
rect 28080 29446 28132 29452
rect 28092 29306 28120 29446
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28092 28490 28120 29242
rect 28080 28484 28132 28490
rect 28080 28426 28132 28432
rect 27896 27056 27948 27062
rect 27896 26998 27948 27004
rect 27908 19446 27936 26998
rect 28276 26217 28304 36060
rect 28356 36042 28408 36048
rect 28460 35193 28488 36246
rect 29012 36009 29040 36722
rect 29564 36310 29592 36722
rect 29918 36408 29974 36417
rect 29918 36343 29974 36352
rect 29552 36304 29604 36310
rect 29552 36246 29604 36252
rect 29932 36106 29960 36343
rect 30024 36281 30052 37198
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30300 36786 30328 37062
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30010 36272 30066 36281
rect 30010 36207 30066 36216
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 28998 36000 29054 36009
rect 28998 35935 29054 35944
rect 30300 35698 30328 36722
rect 30746 36408 30802 36417
rect 30746 36343 30802 36352
rect 30472 36100 30524 36106
rect 30392 36060 30472 36088
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 28446 35184 28502 35193
rect 28446 35119 28502 35128
rect 28356 33856 28408 33862
rect 28356 33798 28408 33804
rect 28368 27674 28396 33798
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28262 26208 28318 26217
rect 28262 26143 28318 26152
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 28000 21486 28028 21966
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 28092 19854 28120 21558
rect 28184 19922 28212 23734
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 27986 19544 28042 19553
rect 27986 19479 28042 19488
rect 27896 19440 27948 19446
rect 27896 19382 27948 19388
rect 28000 19378 28028 19479
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27356 13530 27384 13806
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27448 12850 27476 14282
rect 27908 13258 27936 18634
rect 28092 17678 28120 19246
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 28000 16017 28028 17070
rect 28092 16522 28120 17614
rect 28080 16516 28132 16522
rect 28080 16458 28132 16464
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16250 28212 16458
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28276 16114 28304 23598
rect 28460 22094 28488 35119
rect 29380 32570 29408 35430
rect 29736 35012 29788 35018
rect 29736 34954 29788 34960
rect 29748 34066 29776 34954
rect 29736 34060 29788 34066
rect 29736 34002 29788 34008
rect 29368 32564 29420 32570
rect 29368 32506 29420 32512
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28644 30433 28672 31282
rect 29828 31272 29880 31278
rect 29880 31232 29960 31260
rect 29828 31214 29880 31220
rect 29932 30734 29960 31232
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 28630 30424 28686 30433
rect 28630 30359 28686 30368
rect 29552 30388 29604 30394
rect 29552 30330 29604 30336
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28552 27146 28580 30194
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 28920 28014 28948 29990
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28552 27118 28672 27146
rect 28920 27130 28948 27406
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 28540 24676 28592 24682
rect 28540 24618 28592 24624
rect 28552 23526 28580 24618
rect 28540 23520 28592 23526
rect 28540 23462 28592 23468
rect 28368 22066 28488 22094
rect 28368 19394 28396 22066
rect 28446 21040 28502 21049
rect 28446 20975 28448 20984
rect 28500 20975 28502 20984
rect 28448 20946 28500 20952
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28460 19854 28488 20742
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28368 19366 28488 19394
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28368 18290 28396 19246
rect 28460 18698 28488 19366
rect 28552 18766 28580 23462
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 27986 16008 28042 16017
rect 27986 15943 28042 15952
rect 28368 15162 28396 18226
rect 28538 17776 28594 17785
rect 28538 17711 28594 17720
rect 28552 17678 28580 17711
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28644 17610 28672 27118
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 28908 26784 28960 26790
rect 28908 26726 28960 26732
rect 28920 25265 28948 26726
rect 29012 26586 29040 26862
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 29104 26450 29132 27270
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 29092 26444 29144 26450
rect 29092 26386 29144 26392
rect 29196 26330 29224 26522
rect 29104 26302 29224 26330
rect 29104 25838 29132 26302
rect 29288 26194 29316 30262
rect 29564 29578 29592 30330
rect 29552 29572 29604 29578
rect 29552 29514 29604 29520
rect 29644 29504 29696 29510
rect 29644 29446 29696 29452
rect 29656 28994 29684 29446
rect 29656 28966 29776 28994
rect 29748 28150 29776 28966
rect 29736 28144 29788 28150
rect 29736 28086 29788 28092
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29368 27872 29420 27878
rect 29368 27814 29420 27820
rect 29380 26926 29408 27814
rect 29368 26920 29420 26926
rect 29368 26862 29420 26868
rect 29196 26166 29316 26194
rect 29092 25832 29144 25838
rect 29092 25774 29144 25780
rect 28906 25256 28962 25265
rect 28906 25191 28962 25200
rect 28816 24812 28868 24818
rect 28816 24754 28868 24760
rect 28724 24676 28776 24682
rect 28724 24618 28776 24624
rect 28736 21894 28764 24618
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28448 17332 28500 17338
rect 28448 17274 28500 17280
rect 28460 17134 28488 17274
rect 28448 17128 28500 17134
rect 28540 17128 28592 17134
rect 28448 17070 28500 17076
rect 28538 17096 28540 17105
rect 28592 17096 28594 17105
rect 28538 17031 28594 17040
rect 28736 16114 28764 21830
rect 28828 18698 28856 24754
rect 29000 24608 29052 24614
rect 28920 24556 29000 24562
rect 28920 24550 29052 24556
rect 28920 24534 29040 24550
rect 28920 23662 28948 24534
rect 28908 23656 28960 23662
rect 28908 23598 28960 23604
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 28920 20602 28948 21558
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28920 19854 28948 19994
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28920 18766 28948 19790
rect 29012 19446 29040 20810
rect 29104 20466 29132 25774
rect 29196 20534 29224 26166
rect 29460 24744 29512 24750
rect 29460 24686 29512 24692
rect 29472 24206 29500 24686
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29472 23730 29500 24142
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29276 23588 29328 23594
rect 29276 23530 29328 23536
rect 29184 20528 29236 20534
rect 29184 20470 29236 20476
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 29104 19334 29132 19654
rect 29012 19306 29132 19334
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28816 18692 28868 18698
rect 28816 18634 28868 18640
rect 29012 18290 29040 19306
rect 29092 19168 29144 19174
rect 29092 19110 29144 19116
rect 29104 18426 29132 19110
rect 29092 18420 29144 18426
rect 29092 18362 29144 18368
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29196 17864 29224 18294
rect 29104 17836 29224 17864
rect 29104 17746 29132 17836
rect 29182 17776 29238 17785
rect 29092 17740 29144 17746
rect 29182 17711 29238 17720
rect 29092 17682 29144 17688
rect 29196 17678 29224 17711
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29196 16794 29224 17206
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29288 16522 29316 23530
rect 29472 23186 29500 23666
rect 29368 23180 29420 23186
rect 29368 23122 29420 23128
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29380 21418 29408 23122
rect 29472 22642 29500 23122
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29368 21412 29420 21418
rect 29368 21354 29420 21360
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28552 13938 28580 15574
rect 28724 15428 28776 15434
rect 28724 15370 28776 15376
rect 28632 14408 28684 14414
rect 28632 14350 28684 14356
rect 28540 13932 28592 13938
rect 28540 13874 28592 13880
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27252 8356 27304 8362
rect 27252 8298 27304 8304
rect 27816 2650 27844 10542
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 28092 8974 28120 9318
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28644 3602 28672 14350
rect 28632 3596 28684 3602
rect 28632 3538 28684 3544
rect 28736 2650 28764 15370
rect 29196 15094 29224 15846
rect 29288 15502 29316 16458
rect 29380 16130 29408 21354
rect 29552 20868 29604 20874
rect 29552 20810 29604 20816
rect 29564 20602 29592 20810
rect 29552 20596 29604 20602
rect 29552 20538 29604 20544
rect 29460 19780 29512 19786
rect 29460 19722 29512 19728
rect 29472 17678 29500 19722
rect 29656 19378 29684 27950
rect 29748 25226 29776 28086
rect 29840 26926 29868 30534
rect 29932 30190 29960 30670
rect 30196 30592 30248 30598
rect 30196 30534 30248 30540
rect 30208 30326 30236 30534
rect 30196 30320 30248 30326
rect 30196 30262 30248 30268
rect 29920 30184 29972 30190
rect 29920 30126 29972 30132
rect 29932 29714 29960 30126
rect 29920 29708 29972 29714
rect 29920 29650 29972 29656
rect 30012 27532 30064 27538
rect 30012 27474 30064 27480
rect 30024 27402 30052 27474
rect 30012 27396 30064 27402
rect 30012 27338 30064 27344
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 30024 26058 30052 27338
rect 30392 26518 30420 36060
rect 30472 36042 30524 36048
rect 30470 35728 30526 35737
rect 30470 35663 30472 35672
rect 30524 35663 30526 35672
rect 30472 35634 30524 35640
rect 30564 35012 30616 35018
rect 30564 34954 30616 34960
rect 30576 34746 30604 34954
rect 30564 34740 30616 34746
rect 30564 34682 30616 34688
rect 30576 32978 30604 34682
rect 30760 34542 30788 36343
rect 30944 35698 30972 39200
rect 32232 37346 32260 39200
rect 32232 37318 32352 37346
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 31036 36922 31064 37062
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 32232 36718 32260 37198
rect 32324 36922 32352 37318
rect 32876 36922 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 34060 37324 34112 37330
rect 34060 37266 34112 37272
rect 33140 37188 33192 37194
rect 33140 37130 33192 37136
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 32864 36916 32916 36922
rect 32864 36858 32916 36864
rect 32312 36780 32364 36786
rect 32312 36722 32364 36728
rect 33048 36780 33100 36786
rect 33048 36722 33100 36728
rect 32220 36712 32272 36718
rect 32220 36654 32272 36660
rect 31668 36576 31720 36582
rect 31668 36518 31720 36524
rect 31392 36032 31444 36038
rect 31392 35974 31444 35980
rect 31404 35850 31432 35974
rect 31220 35822 31432 35850
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30932 35692 30984 35698
rect 30932 35634 30984 35640
rect 30852 34610 30880 35634
rect 31024 34944 31076 34950
rect 31024 34886 31076 34892
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30748 34536 30800 34542
rect 30748 34478 30800 34484
rect 31036 33930 31064 34886
rect 31024 33924 31076 33930
rect 31024 33866 31076 33872
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 30656 32836 30708 32842
rect 30656 32778 30708 32784
rect 30564 31408 30616 31414
rect 30564 31350 30616 31356
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30484 30802 30512 31078
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30576 30433 30604 31350
rect 30562 30424 30618 30433
rect 30562 30359 30618 30368
rect 30668 27130 30696 32778
rect 31220 31142 31248 35822
rect 31392 35760 31444 35766
rect 31392 35702 31444 35708
rect 31300 34536 31352 34542
rect 31300 34478 31352 34484
rect 31312 31686 31340 34478
rect 31300 31680 31352 31686
rect 31300 31622 31352 31628
rect 31208 31136 31260 31142
rect 31208 31078 31260 31084
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 31312 29073 31340 30194
rect 31404 30054 31432 35702
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31496 35154 31524 35430
rect 31484 35148 31536 35154
rect 31484 35090 31536 35096
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 31484 34672 31536 34678
rect 31484 34614 31536 34620
rect 31496 30326 31524 34614
rect 31588 33658 31616 34954
rect 31576 33652 31628 33658
rect 31576 33594 31628 33600
rect 31680 32842 31708 36518
rect 32232 36242 32260 36654
rect 32324 36417 32352 36722
rect 32310 36408 32366 36417
rect 33060 36378 33088 36722
rect 33152 36553 33180 37130
rect 33876 36848 33928 36854
rect 33876 36790 33928 36796
rect 33784 36576 33836 36582
rect 33138 36544 33194 36553
rect 33784 36518 33836 36524
rect 33138 36479 33194 36488
rect 33796 36378 33824 36518
rect 32310 36343 32366 36352
rect 33048 36372 33100 36378
rect 33048 36314 33100 36320
rect 33784 36372 33836 36378
rect 33784 36314 33836 36320
rect 33888 36310 33916 36790
rect 33876 36304 33928 36310
rect 33876 36246 33928 36252
rect 32220 36236 32272 36242
rect 32220 36178 32272 36184
rect 31760 36100 31812 36106
rect 31760 36042 31812 36048
rect 31668 32836 31720 32842
rect 31668 32778 31720 32784
rect 31772 32434 31800 36042
rect 32232 35154 32260 36178
rect 33968 36032 34020 36038
rect 33968 35974 34020 35980
rect 33980 35834 34008 35974
rect 33968 35828 34020 35834
rect 33968 35770 34020 35776
rect 32864 35556 32916 35562
rect 32864 35498 32916 35504
rect 31852 35148 31904 35154
rect 31852 35090 31904 35096
rect 32220 35148 32272 35154
rect 32220 35090 32272 35096
rect 31864 33930 31892 35090
rect 32876 35018 32904 35498
rect 34072 35306 34100 37266
rect 34440 37244 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35162 37360 35218 37369
rect 35162 37295 35164 37304
rect 35216 37295 35218 37304
rect 35164 37266 35216 37272
rect 34520 37256 34572 37262
rect 34440 37216 34520 37244
rect 34520 37198 34572 37204
rect 34152 37120 34204 37126
rect 34152 37062 34204 37068
rect 34164 35894 34192 37062
rect 34428 36712 34480 36718
rect 34428 36654 34480 36660
rect 34704 36712 34756 36718
rect 34704 36654 34756 36660
rect 34440 36242 34468 36654
rect 34428 36236 34480 36242
rect 34428 36178 34480 36184
rect 34520 36100 34572 36106
rect 34520 36042 34572 36048
rect 34612 36100 34664 36106
rect 34612 36042 34664 36048
rect 34164 35866 34284 35894
rect 34072 35278 34192 35306
rect 32956 35148 33008 35154
rect 32956 35090 33008 35096
rect 32864 35012 32916 35018
rect 32864 34954 32916 34960
rect 31852 33924 31904 33930
rect 31852 33866 31904 33872
rect 31864 33833 31892 33866
rect 32404 33856 32456 33862
rect 31850 33824 31906 33833
rect 32404 33798 32456 33804
rect 31850 33759 31906 33768
rect 32416 33658 32444 33798
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32876 33590 32904 34954
rect 32968 33930 32996 35090
rect 33416 34672 33468 34678
rect 33416 34614 33468 34620
rect 33428 34474 33456 34614
rect 34164 34610 34192 35278
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 33416 34468 33468 34474
rect 33416 34410 33468 34416
rect 34164 33998 34192 34546
rect 34152 33992 34204 33998
rect 34152 33934 34204 33940
rect 32956 33924 33008 33930
rect 32956 33866 33008 33872
rect 32864 33584 32916 33590
rect 32864 33526 32916 33532
rect 32968 33522 32996 33866
rect 33416 33856 33468 33862
rect 33416 33798 33468 33804
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32312 33380 32364 33386
rect 32312 33322 32364 33328
rect 32324 32774 32352 33322
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 32312 32768 32364 32774
rect 32312 32710 32364 32716
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 32128 31272 32180 31278
rect 32128 31214 32180 31220
rect 31576 31136 31628 31142
rect 31576 31078 31628 31084
rect 31484 30320 31536 30326
rect 31484 30262 31536 30268
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31588 29170 31616 31078
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 32048 30433 32076 30602
rect 32034 30424 32090 30433
rect 32034 30359 32090 30368
rect 32140 30054 32168 31214
rect 31668 30048 31720 30054
rect 31666 30016 31668 30025
rect 32128 30048 32180 30054
rect 31720 30016 31722 30025
rect 32128 29990 32180 29996
rect 31666 29951 31722 29960
rect 31668 29572 31720 29578
rect 31668 29514 31720 29520
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31298 29064 31354 29073
rect 31298 28999 31354 29008
rect 31116 28552 31168 28558
rect 31116 28494 31168 28500
rect 31128 28014 31156 28494
rect 31680 28422 31708 29514
rect 32140 28914 32168 29990
rect 32220 29572 32272 29578
rect 32220 29514 32272 29520
rect 32232 29073 32260 29514
rect 32324 29102 32352 32710
rect 32404 31272 32456 31278
rect 32404 31214 32456 31220
rect 32772 31272 32824 31278
rect 32772 31214 32824 31220
rect 32416 30734 32444 31214
rect 32404 30728 32456 30734
rect 32404 30670 32456 30676
rect 32416 29714 32444 30670
rect 32404 29708 32456 29714
rect 32404 29650 32456 29656
rect 32416 29170 32444 29650
rect 32404 29164 32456 29170
rect 32404 29106 32456 29112
rect 32312 29096 32364 29102
rect 32218 29064 32274 29073
rect 32312 29038 32364 29044
rect 32218 28999 32274 29008
rect 32588 28960 32640 28966
rect 32140 28886 32260 28914
rect 32588 28902 32640 28908
rect 32036 28484 32088 28490
rect 32036 28426 32088 28432
rect 31668 28416 31720 28422
rect 31668 28358 31720 28364
rect 31300 28076 31352 28082
rect 31300 28018 31352 28024
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 30656 27124 30708 27130
rect 30656 27066 30708 27072
rect 30380 26512 30432 26518
rect 30380 26454 30432 26460
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30104 26308 30156 26314
rect 30104 26250 30156 26256
rect 29932 26030 30052 26058
rect 29736 25220 29788 25226
rect 29736 25162 29788 25168
rect 29748 23118 29776 25162
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29828 22500 29880 22506
rect 29828 22442 29880 22448
rect 29840 21486 29868 22442
rect 29932 22030 29960 26030
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 29736 21412 29788 21418
rect 29736 21354 29788 21360
rect 29748 20942 29776 21354
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29748 19922 29776 20334
rect 29932 19922 29960 21830
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29550 19136 29606 19145
rect 29550 19071 29606 19080
rect 29460 17672 29512 17678
rect 29458 17640 29460 17649
rect 29512 17640 29514 17649
rect 29458 17575 29514 17584
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29472 16250 29500 17206
rect 29460 16244 29512 16250
rect 29460 16186 29512 16192
rect 29380 16102 29500 16130
rect 29564 16114 29592 19071
rect 29748 18222 29776 19858
rect 29920 19236 29972 19242
rect 29920 19178 29972 19184
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29644 17808 29696 17814
rect 29644 17750 29696 17756
rect 29656 17270 29684 17750
rect 29644 17264 29696 17270
rect 29644 17206 29696 17212
rect 29276 15496 29328 15502
rect 29276 15438 29328 15444
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28908 14000 28960 14006
rect 28908 13942 28960 13948
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28828 11218 28856 12718
rect 28816 11212 28868 11218
rect 28816 11154 28868 11160
rect 28920 10674 28948 13942
rect 29012 13938 29040 14214
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29380 12986 29408 15438
rect 29472 14346 29500 16102
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29748 14958 29776 18158
rect 29932 16454 29960 19178
rect 30024 17882 30052 25910
rect 30116 23662 30144 26250
rect 30576 25906 30604 26318
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 30012 17876 30064 17882
rect 30012 17818 30064 17824
rect 30116 16946 30144 23598
rect 30208 22574 30236 24686
rect 30380 23792 30432 23798
rect 30380 23734 30432 23740
rect 30196 22568 30248 22574
rect 30196 22510 30248 22516
rect 30392 20602 30420 23734
rect 30472 22704 30524 22710
rect 30472 22646 30524 22652
rect 30380 20596 30432 20602
rect 30380 20538 30432 20544
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 18850 30420 19314
rect 30484 18970 30512 22646
rect 30564 22568 30616 22574
rect 30564 22510 30616 22516
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30392 18822 30512 18850
rect 30484 18766 30512 18822
rect 30380 18760 30432 18766
rect 30380 18702 30432 18708
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30392 18601 30420 18702
rect 30378 18592 30434 18601
rect 30378 18527 30434 18536
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30208 17882 30236 18362
rect 30472 18352 30524 18358
rect 30472 18294 30524 18300
rect 30378 17912 30434 17921
rect 30196 17876 30248 17882
rect 30378 17847 30434 17856
rect 30196 17818 30248 17824
rect 30392 17814 30420 17847
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30300 16946 30328 17138
rect 30116 16918 30328 16946
rect 30116 16658 30144 16918
rect 30392 16726 30420 17614
rect 30380 16720 30432 16726
rect 30380 16662 30432 16668
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 30484 16590 30512 18294
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 30208 16114 30236 16458
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 30576 14414 30604 22510
rect 30668 21418 30696 27066
rect 31024 27056 31076 27062
rect 31024 26998 31076 27004
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30944 26314 30972 26386
rect 30932 26308 30984 26314
rect 30932 26250 30984 26256
rect 30748 25832 30800 25838
rect 30748 25774 30800 25780
rect 30760 24993 30788 25774
rect 30746 24984 30802 24993
rect 30746 24919 30802 24928
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30656 21412 30708 21418
rect 30656 21354 30708 21360
rect 30852 21146 30880 24754
rect 31036 22094 31064 26998
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 31128 23322 31156 24006
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31128 22778 31156 23258
rect 31220 23089 31248 26726
rect 31206 23080 31262 23089
rect 31206 23015 31262 23024
rect 31312 22930 31340 28018
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31392 27668 31444 27674
rect 31392 27610 31444 27616
rect 31404 23526 31432 27610
rect 31680 27538 31708 27950
rect 31668 27532 31720 27538
rect 31668 27474 31720 27480
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31220 22902 31340 22930
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 30944 22066 31064 22094
rect 30840 21140 30892 21146
rect 30840 21082 30892 21088
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30760 20890 30788 20946
rect 30668 20862 30788 20890
rect 30668 19530 30696 20862
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 30852 20534 30880 20742
rect 30840 20528 30892 20534
rect 30746 20496 30802 20505
rect 30840 20470 30892 20476
rect 30746 20431 30802 20440
rect 30760 20398 30788 20431
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30668 19502 30788 19530
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30668 18426 30696 19382
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30760 17066 30788 19502
rect 30852 18630 30880 19654
rect 30944 18737 30972 22066
rect 31220 19009 31248 22902
rect 31300 22160 31352 22166
rect 31300 22102 31352 22108
rect 31312 19174 31340 22102
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 31206 19000 31262 19009
rect 31206 18935 31262 18944
rect 30930 18728 30986 18737
rect 30930 18663 30986 18672
rect 31116 18692 31168 18698
rect 31116 18634 31168 18640
rect 30840 18624 30892 18630
rect 30840 18566 30892 18572
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 30746 16008 30802 16017
rect 30852 15994 30880 18566
rect 31128 18222 31156 18634
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31022 17640 31078 17649
rect 31022 17575 31078 17584
rect 30932 17060 30984 17066
rect 30932 17002 30984 17008
rect 30944 16833 30972 17002
rect 30930 16824 30986 16833
rect 30930 16759 30986 16768
rect 31036 16590 31064 17575
rect 31312 16640 31340 19110
rect 31404 18290 31432 21422
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31220 16612 31340 16640
rect 31024 16584 31076 16590
rect 31116 16584 31168 16590
rect 31024 16526 31076 16532
rect 31114 16552 31116 16561
rect 31168 16552 31170 16561
rect 31036 16153 31064 16526
rect 31114 16487 31170 16496
rect 31022 16144 31078 16153
rect 31022 16079 31078 16088
rect 30802 15966 30880 15994
rect 30746 15943 30802 15952
rect 30760 15502 30788 15943
rect 30930 15736 30986 15745
rect 30930 15671 30986 15680
rect 30944 15638 30972 15671
rect 30932 15632 30984 15638
rect 30932 15574 30984 15580
rect 30748 15496 30800 15502
rect 30748 15438 30800 15444
rect 30760 14482 30788 15438
rect 31220 15026 31248 16612
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 31312 16114 31340 16458
rect 31496 16250 31524 27338
rect 31680 26994 31708 27474
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31668 26988 31720 26994
rect 31668 26930 31720 26936
rect 31680 25906 31708 26930
rect 31772 26926 31800 27406
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31668 25900 31720 25906
rect 31668 25842 31720 25848
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31588 22094 31616 24142
rect 31588 22066 31708 22094
rect 31680 21010 31708 22066
rect 31668 21004 31720 21010
rect 31668 20946 31720 20952
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 31576 19712 31628 19718
rect 31576 19654 31628 19660
rect 31588 19446 31616 19654
rect 31680 19446 31708 19790
rect 31576 19440 31628 19446
rect 31576 19382 31628 19388
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 31668 19168 31720 19174
rect 31668 19110 31720 19116
rect 31574 18864 31630 18873
rect 31574 18799 31630 18808
rect 31588 18766 31616 18799
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31588 18630 31616 18702
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 31680 18442 31708 19110
rect 31588 18414 31708 18442
rect 31484 16244 31536 16250
rect 31484 16186 31536 16192
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31588 15570 31616 18414
rect 31772 18272 31800 26862
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31864 22817 31892 22986
rect 31850 22808 31906 22817
rect 31850 22743 31906 22752
rect 31852 22704 31904 22710
rect 31852 22646 31904 22652
rect 31864 21418 31892 22646
rect 32048 22094 32076 28426
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 32140 24410 32168 26250
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32232 22234 32260 28886
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32324 25294 32352 25638
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32324 24818 32352 25230
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32324 24274 32352 24754
rect 32404 24404 32456 24410
rect 32404 24346 32456 24352
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 32324 23730 32352 24210
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32324 23186 32352 23666
rect 32312 23180 32364 23186
rect 32312 23122 32364 23128
rect 32324 22574 32352 23122
rect 32312 22568 32364 22574
rect 32312 22510 32364 22516
rect 32416 22522 32444 24346
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32324 22098 32352 22510
rect 32416 22494 32536 22522
rect 32404 22228 32456 22234
rect 32404 22170 32456 22176
rect 31956 22066 32076 22094
rect 32312 22092 32364 22098
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31852 20392 31904 20398
rect 31852 20334 31904 20340
rect 31864 19990 31892 20334
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 31956 18358 31984 22066
rect 32312 22034 32364 22040
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32140 20534 32168 20878
rect 32128 20528 32180 20534
rect 32128 20470 32180 20476
rect 32140 20058 32168 20470
rect 32416 20466 32444 22170
rect 32508 20942 32536 22494
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32600 20641 32628 28902
rect 32678 23080 32734 23089
rect 32678 23015 32734 23024
rect 32692 22982 32720 23015
rect 32680 22976 32732 22982
rect 32680 22918 32732 22924
rect 32680 22568 32732 22574
rect 32680 22510 32732 22516
rect 32586 20632 32642 20641
rect 32586 20567 32642 20576
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 32048 19530 32076 19790
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32048 19502 32168 19530
rect 32036 19372 32088 19378
rect 32036 19314 32088 19320
rect 31944 18352 31996 18358
rect 31944 18294 31996 18300
rect 31852 18284 31904 18290
rect 31772 18244 31852 18272
rect 31852 18226 31904 18232
rect 31852 18080 31904 18086
rect 31852 18022 31904 18028
rect 31864 17134 31892 18022
rect 31944 17740 31996 17746
rect 31944 17682 31996 17688
rect 31852 17128 31904 17134
rect 31852 17070 31904 17076
rect 31758 16960 31814 16969
rect 31758 16895 31814 16904
rect 31772 16658 31800 16895
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31760 16448 31812 16454
rect 31760 16390 31812 16396
rect 31668 16040 31720 16046
rect 31668 15982 31720 15988
rect 31576 15564 31628 15570
rect 31576 15506 31628 15512
rect 31392 15360 31444 15366
rect 31392 15302 31444 15308
rect 31404 15026 31432 15302
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 29460 14340 29512 14346
rect 29460 14282 29512 14288
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 29012 7886 29040 10406
rect 29000 7880 29052 7886
rect 29000 7822 29052 7828
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 29288 2582 29316 12786
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 29840 5710 29868 12174
rect 30392 9654 30420 14214
rect 30852 14006 30880 14758
rect 30840 14000 30892 14006
rect 30840 13942 30892 13948
rect 31680 13870 31708 15982
rect 31772 15366 31800 16390
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31864 15178 31892 17070
rect 31956 17066 31984 17682
rect 31944 17060 31996 17066
rect 31944 17002 31996 17008
rect 31956 15434 31984 17002
rect 32048 16046 32076 19314
rect 32140 17746 32168 19502
rect 32232 18426 32260 19722
rect 32324 19553 32352 20198
rect 32310 19544 32366 19553
rect 32310 19479 32366 19488
rect 32508 19310 32536 20198
rect 32496 19304 32548 19310
rect 32496 19246 32548 19252
rect 32312 19236 32364 19242
rect 32312 19178 32364 19184
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 32128 17740 32180 17746
rect 32128 17682 32180 17688
rect 32220 16176 32272 16182
rect 32220 16118 32272 16124
rect 32036 16040 32088 16046
rect 32036 15982 32088 15988
rect 32036 15904 32088 15910
rect 32036 15846 32088 15852
rect 31944 15428 31996 15434
rect 31944 15370 31996 15376
rect 31772 15150 31892 15178
rect 31772 14618 31800 15150
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31864 14482 31892 14758
rect 32048 14618 32076 15846
rect 32232 15638 32260 16118
rect 32220 15632 32272 15638
rect 32220 15574 32272 15580
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 32128 14884 32180 14890
rect 32128 14826 32180 14832
rect 32036 14612 32088 14618
rect 32036 14554 32088 14560
rect 31852 14476 31904 14482
rect 31852 14418 31904 14424
rect 31668 13864 31720 13870
rect 31668 13806 31720 13812
rect 31852 13864 31904 13870
rect 31852 13806 31904 13812
rect 31680 11218 31708 13806
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31864 11150 31892 13806
rect 32048 11150 32076 14554
rect 32140 14482 32168 14826
rect 32232 14618 32260 14894
rect 32324 14890 32352 19178
rect 32402 19000 32458 19009
rect 32402 18935 32458 18944
rect 32416 18902 32444 18935
rect 32404 18896 32456 18902
rect 32404 18838 32456 18844
rect 32586 18728 32642 18737
rect 32586 18663 32588 18672
rect 32640 18663 32642 18672
rect 32588 18634 32640 18640
rect 32692 16658 32720 22510
rect 32784 19242 32812 31214
rect 33048 30048 33100 30054
rect 33048 29990 33100 29996
rect 33060 29782 33088 29990
rect 33048 29776 33100 29782
rect 33048 29718 33100 29724
rect 33152 29510 33180 32778
rect 33428 32570 33456 33798
rect 34164 33046 34192 33934
rect 34152 33040 34204 33046
rect 34152 32982 34204 32988
rect 33968 32972 34020 32978
rect 33968 32914 34020 32920
rect 33416 32564 33468 32570
rect 33416 32506 33468 32512
rect 33784 31340 33836 31346
rect 33784 31282 33836 31288
rect 33416 30660 33468 30666
rect 33416 30602 33468 30608
rect 33140 29504 33192 29510
rect 33140 29446 33192 29452
rect 33152 29050 33180 29446
rect 33232 29232 33284 29238
rect 33230 29200 33232 29209
rect 33284 29200 33286 29209
rect 33230 29135 33286 29144
rect 33060 29022 33180 29050
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32876 27674 32904 28358
rect 32864 27668 32916 27674
rect 32864 27610 32916 27616
rect 32772 19236 32824 19242
rect 32772 19178 32824 19184
rect 32772 18896 32824 18902
rect 32772 18838 32824 18844
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32784 16590 32812 18838
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 32772 16584 32824 16590
rect 32772 16526 32824 16532
rect 32416 16182 32444 16526
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32404 16176 32456 16182
rect 32404 16118 32456 16124
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32128 14476 32180 14482
rect 32128 14418 32180 14424
rect 32312 14408 32364 14414
rect 32312 14350 32364 14356
rect 32324 12986 32352 14350
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32324 12238 32352 12922
rect 32312 12232 32364 12238
rect 32312 12174 32364 12180
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 32416 10810 32444 15982
rect 32508 15094 32536 16390
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32600 15706 32628 15846
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32876 15570 32904 27610
rect 32956 23520 33008 23526
rect 32956 23462 33008 23468
rect 32968 21962 32996 23462
rect 32956 21956 33008 21962
rect 32956 21898 33008 21904
rect 32968 21049 32996 21898
rect 32954 21040 33010 21049
rect 32954 20975 33010 20984
rect 33060 18902 33088 29022
rect 33428 28150 33456 30602
rect 33600 29300 33652 29306
rect 33600 29242 33652 29248
rect 33416 28144 33468 28150
rect 33416 28086 33468 28092
rect 33416 27872 33468 27878
rect 33416 27814 33468 27820
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 33140 21072 33192 21078
rect 33140 21014 33192 21020
rect 33048 18896 33100 18902
rect 33048 18838 33100 18844
rect 32956 18760 33008 18766
rect 33008 18720 33088 18748
rect 32956 18702 33008 18708
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 32968 18193 32996 18226
rect 32954 18184 33010 18193
rect 32954 18119 33010 18128
rect 33060 17785 33088 18720
rect 33046 17776 33102 17785
rect 33046 17711 33102 17720
rect 33060 16658 33088 17711
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 32864 15564 32916 15570
rect 32864 15506 32916 15512
rect 32956 15360 33008 15366
rect 32956 15302 33008 15308
rect 33046 15328 33102 15337
rect 32496 15088 32548 15094
rect 32496 15030 32548 15036
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32494 13424 32550 13433
rect 32494 13359 32550 13368
rect 32508 12850 32536 13359
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30012 7744 30064 7750
rect 30012 7686 30064 7692
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 29276 2576 29328 2582
rect 29276 2518 29328 2524
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25792 800 25820 2382
rect 27080 800 27108 2382
rect 27724 800 27752 2382
rect 29012 800 29040 2382
rect 29840 2378 29868 5646
rect 30024 2514 30052 7686
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30392 2446 30420 8774
rect 32508 4622 32536 11018
rect 32784 7546 32812 14010
rect 32862 13560 32918 13569
rect 32862 13495 32864 13504
rect 32916 13495 32918 13504
rect 32864 13466 32916 13472
rect 32968 13394 32996 15302
rect 33046 15263 33102 15272
rect 33060 15162 33088 15263
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33152 13462 33180 21014
rect 33244 18970 33272 27270
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 33232 18760 33284 18766
rect 33232 18702 33284 18708
rect 33244 18601 33272 18702
rect 33230 18592 33286 18601
rect 33230 18527 33286 18536
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 33244 17610 33272 18022
rect 33232 17604 33284 17610
rect 33232 17546 33284 17552
rect 33230 16824 33286 16833
rect 33230 16759 33286 16768
rect 33244 15638 33272 16759
rect 33322 16688 33378 16697
rect 33322 16623 33378 16632
rect 33336 16046 33364 16623
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33428 15858 33456 27814
rect 33612 26926 33640 29242
rect 33600 26920 33652 26926
rect 33600 26862 33652 26868
rect 33508 20936 33560 20942
rect 33508 20878 33560 20884
rect 33520 17082 33548 20878
rect 33612 17218 33640 26862
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33704 24993 33732 25842
rect 33690 24984 33746 24993
rect 33690 24919 33746 24928
rect 33796 22522 33824 31282
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 33888 25702 33916 25978
rect 33876 25696 33928 25702
rect 33876 25638 33928 25644
rect 33876 24744 33928 24750
rect 33876 24686 33928 24692
rect 33704 22494 33824 22522
rect 33704 20262 33732 22494
rect 33888 22094 33916 24686
rect 33796 22066 33916 22094
rect 33796 21894 33824 22066
rect 33784 21888 33836 21894
rect 33784 21830 33836 21836
rect 33796 20942 33824 21830
rect 33980 21690 34008 32914
rect 34256 32502 34284 35866
rect 34336 35828 34388 35834
rect 34336 35770 34388 35776
rect 34348 35222 34376 35770
rect 34532 35290 34560 36042
rect 34520 35284 34572 35290
rect 34520 35226 34572 35232
rect 34336 35216 34388 35222
rect 34336 35158 34388 35164
rect 34336 34944 34388 34950
rect 34336 34886 34388 34892
rect 34244 32496 34296 32502
rect 34244 32438 34296 32444
rect 34348 31278 34376 34886
rect 34624 34626 34652 36042
rect 34716 35766 34744 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35452 35894 35480 39200
rect 36096 37126 36124 39200
rect 37186 37496 37242 37505
rect 37186 37431 37242 37440
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 35716 36848 35768 36854
rect 35716 36790 35768 36796
rect 35360 35866 35480 35894
rect 34704 35760 34756 35766
rect 34704 35702 34756 35708
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 34532 34598 34652 34626
rect 34532 33454 34560 34598
rect 34612 34536 34664 34542
rect 34612 34478 34664 34484
rect 34624 34066 34652 34478
rect 34612 34060 34664 34066
rect 34612 34002 34664 34008
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 34336 31272 34388 31278
rect 34336 31214 34388 31220
rect 34244 31136 34296 31142
rect 34244 31078 34296 31084
rect 34256 30802 34284 31078
rect 34244 30796 34296 30802
rect 34244 30738 34296 30744
rect 34532 30138 34560 33254
rect 34624 33114 34652 34002
rect 34716 33590 34744 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34536 34848 34542
rect 34796 34478 34848 34484
rect 34808 34202 34836 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 34796 33924 34848 33930
rect 34796 33866 34848 33872
rect 34704 33584 34756 33590
rect 34704 33526 34756 33532
rect 34612 33108 34664 33114
rect 34612 33050 34664 33056
rect 34808 32978 34836 33866
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 34808 32434 34836 32914
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34610 30968 34666 30977
rect 34934 30971 35242 30980
rect 34610 30903 34612 30912
rect 34664 30903 34666 30912
rect 34612 30874 34664 30880
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 34716 30258 34744 30670
rect 35072 30320 35124 30326
rect 35072 30262 35124 30268
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 34440 30110 34560 30138
rect 34612 30184 34664 30190
rect 34612 30126 34664 30132
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34440 29458 34468 30110
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 34072 24750 34100 28426
rect 34060 24744 34112 24750
rect 34060 24686 34112 24692
rect 33968 21684 34020 21690
rect 33968 21626 34020 21632
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 33980 21146 34008 21286
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 33876 21072 33928 21078
rect 33876 21014 33928 21020
rect 33888 20942 33916 21014
rect 33784 20936 33836 20942
rect 33784 20878 33836 20884
rect 33876 20936 33928 20942
rect 33876 20878 33928 20884
rect 33784 20596 33836 20602
rect 33784 20538 33836 20544
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33796 19718 33824 20538
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33874 19952 33930 19961
rect 33874 19887 33876 19896
rect 33928 19887 33930 19896
rect 33876 19858 33928 19864
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33690 19272 33746 19281
rect 33690 19207 33746 19216
rect 33704 18970 33732 19207
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33796 17610 33824 19654
rect 33876 18624 33928 18630
rect 33876 18566 33928 18572
rect 33888 18290 33916 18566
rect 33876 18284 33928 18290
rect 33876 18226 33928 18232
rect 33888 18154 33916 18226
rect 33876 18148 33928 18154
rect 33876 18090 33928 18096
rect 33980 17746 34008 20334
rect 33968 17740 34020 17746
rect 33968 17682 34020 17688
rect 33784 17604 33836 17610
rect 33784 17546 33836 17552
rect 33980 17338 34008 17682
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 33612 17190 33916 17218
rect 33520 17054 33640 17082
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33520 16017 33548 16526
rect 33506 16008 33562 16017
rect 33506 15943 33562 15952
rect 33336 15830 33456 15858
rect 33232 15632 33284 15638
rect 33232 15574 33284 15580
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 33244 13938 33272 14962
rect 33336 14958 33364 15830
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33336 14346 33364 14894
rect 33416 14816 33468 14822
rect 33416 14758 33468 14764
rect 33428 14346 33456 14758
rect 33520 14550 33548 14894
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 33416 14340 33468 14346
rect 33416 14282 33468 14288
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33508 13796 33560 13802
rect 33508 13738 33560 13744
rect 33140 13456 33192 13462
rect 33140 13398 33192 13404
rect 32956 13388 33008 13394
rect 32956 13330 33008 13336
rect 33138 13288 33194 13297
rect 32864 13252 32916 13258
rect 33138 13223 33194 13232
rect 32864 13194 32916 13200
rect 32876 12442 32904 13194
rect 33152 12850 33180 13223
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33520 12714 33548 13738
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 32772 7540 32824 7546
rect 32772 7482 32824 7488
rect 33152 7410 33180 12582
rect 33416 12436 33468 12442
rect 33416 12378 33468 12384
rect 33428 12345 33456 12378
rect 33414 12336 33470 12345
rect 33414 12271 33470 12280
rect 33612 12238 33640 17054
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33704 16250 33732 16390
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33784 16176 33836 16182
rect 33784 16118 33836 16124
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33704 13802 33732 15982
rect 33796 15706 33824 16118
rect 33784 15700 33836 15706
rect 33784 15642 33836 15648
rect 33692 13796 33744 13802
rect 33692 13738 33744 13744
rect 33690 13696 33746 13705
rect 33690 13631 33746 13640
rect 33704 13326 33732 13631
rect 33692 13320 33744 13326
rect 33692 13262 33744 13268
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 33690 12744 33746 12753
rect 33690 12679 33692 12688
rect 33744 12679 33746 12688
rect 33692 12650 33744 12656
rect 33600 12232 33652 12238
rect 33600 12174 33652 12180
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 32496 4616 32548 4622
rect 32496 4558 32548 4564
rect 33796 3738 33824 12854
rect 33888 11218 33916 17190
rect 33968 17060 34020 17066
rect 33968 17002 34020 17008
rect 33980 14482 34008 17002
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 33968 14000 34020 14006
rect 33968 13942 34020 13948
rect 33980 13530 34008 13942
rect 33968 13524 34020 13530
rect 33968 13466 34020 13472
rect 34072 11762 34100 24686
rect 34164 24410 34192 29446
rect 34440 29430 34560 29458
rect 34428 27056 34480 27062
rect 34428 26998 34480 27004
rect 34440 26353 34468 26998
rect 34426 26344 34482 26353
rect 34426 26279 34482 26288
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 34164 20942 34192 24346
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 34256 22642 34284 24210
rect 34428 24132 34480 24138
rect 34428 24074 34480 24080
rect 34336 23656 34388 23662
rect 34336 23598 34388 23604
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34256 21622 34284 22578
rect 34348 22438 34376 23598
rect 34336 22432 34388 22438
rect 34336 22374 34388 22380
rect 34244 21616 34296 21622
rect 34244 21558 34296 21564
rect 34348 21554 34376 22374
rect 34336 21548 34388 21554
rect 34336 21490 34388 21496
rect 34336 21412 34388 21418
rect 34336 21354 34388 21360
rect 34244 21072 34296 21078
rect 34244 21014 34296 21020
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 34152 20596 34204 20602
rect 34152 20538 34204 20544
rect 34164 20398 34192 20538
rect 34152 20392 34204 20398
rect 34152 20334 34204 20340
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 34164 19446 34192 19994
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 34164 17270 34192 19110
rect 34256 18154 34284 21014
rect 34348 18426 34376 21354
rect 34440 21078 34468 24074
rect 34532 23526 34560 29430
rect 34624 25770 34652 30126
rect 34716 29714 34744 30194
rect 35084 30190 35112 30262
rect 35072 30184 35124 30190
rect 35072 30126 35124 30132
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29850 35388 35866
rect 35728 35834 35756 36790
rect 36188 36689 36216 37198
rect 36728 36916 36780 36922
rect 36728 36858 36780 36864
rect 36174 36680 36230 36689
rect 35808 36644 35860 36650
rect 36174 36615 36230 36624
rect 35808 36586 35860 36592
rect 35820 36242 35848 36586
rect 36176 36576 36228 36582
rect 36176 36518 36228 36524
rect 35808 36236 35860 36242
rect 35808 36178 35860 36184
rect 35716 35828 35768 35834
rect 35716 35770 35768 35776
rect 35820 35698 35848 36178
rect 36188 36122 36216 36518
rect 35912 36094 36216 36122
rect 35912 36038 35940 36094
rect 35900 36032 35952 36038
rect 35900 35974 35952 35980
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35808 35692 35860 35698
rect 35808 35634 35860 35640
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 35452 34066 35480 35566
rect 36004 35562 36032 35974
rect 36740 35834 36768 36858
rect 36820 36576 36872 36582
rect 36820 36518 36872 36524
rect 36832 36106 36860 36518
rect 37200 36174 37228 37431
rect 37384 36922 37412 39200
rect 37462 38856 37518 38865
rect 37462 38791 37518 38800
rect 37476 37330 37504 38791
rect 37464 37324 37516 37330
rect 37464 37266 37516 37272
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 37554 36816 37610 36825
rect 37554 36751 37610 36760
rect 37568 36310 37596 36751
rect 37924 36372 37976 36378
rect 37924 36314 37976 36320
rect 37556 36304 37608 36310
rect 37556 36246 37608 36252
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 36820 36100 36872 36106
rect 36820 36042 36872 36048
rect 36728 35828 36780 35834
rect 36728 35770 36780 35776
rect 36820 35692 36872 35698
rect 36820 35634 36872 35640
rect 35992 35556 36044 35562
rect 35992 35498 36044 35504
rect 35624 34672 35676 34678
rect 35624 34614 35676 34620
rect 35636 34406 35664 34614
rect 35900 34536 35952 34542
rect 35900 34478 35952 34484
rect 35624 34400 35676 34406
rect 35624 34342 35676 34348
rect 35440 34060 35492 34066
rect 35440 34002 35492 34008
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 34704 29708 34756 29714
rect 34704 29650 34756 29656
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34808 28014 34836 28494
rect 34796 28008 34848 28014
rect 34796 27950 34848 27956
rect 34808 27538 34836 27950
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 34704 26784 34756 26790
rect 34704 26726 34756 26732
rect 34716 25974 34744 26726
rect 34808 26450 34836 27474
rect 35452 26790 35480 34002
rect 35532 33516 35584 33522
rect 35532 33458 35584 33464
rect 35544 33425 35572 33458
rect 35530 33416 35586 33425
rect 35530 33351 35586 33360
rect 35636 31754 35664 34342
rect 35912 32366 35940 34478
rect 35900 32360 35952 32366
rect 35900 32302 35952 32308
rect 35544 31726 35664 31754
rect 35440 26784 35492 26790
rect 35440 26726 35492 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 34612 25764 34664 25770
rect 34612 25706 34664 25712
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34624 22114 34652 25706
rect 34532 22086 34652 22114
rect 34428 21072 34480 21078
rect 34428 21014 34480 21020
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34336 18420 34388 18426
rect 34336 18362 34388 18368
rect 34244 18148 34296 18154
rect 34244 18090 34296 18096
rect 34440 18034 34468 19654
rect 34532 19530 34560 22086
rect 34612 21548 34664 21554
rect 34612 21490 34664 21496
rect 34624 19718 34652 21490
rect 34612 19712 34664 19718
rect 34612 19654 34664 19660
rect 34532 19502 34652 19530
rect 34624 19334 34652 19502
rect 34256 18006 34468 18034
rect 34532 19306 34652 19334
rect 34152 17264 34204 17270
rect 34152 17206 34204 17212
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34164 16046 34192 17070
rect 34152 16040 34204 16046
rect 34152 15982 34204 15988
rect 34256 15026 34284 18006
rect 34532 17746 34560 19306
rect 34612 19236 34664 19242
rect 34612 19178 34664 19184
rect 34624 18698 34652 19178
rect 34716 18902 34744 25910
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34808 23798 34836 24142
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 34796 23792 34848 23798
rect 34796 23734 34848 23740
rect 34808 23186 34836 23734
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23180 34848 23186
rect 34796 23122 34848 23128
rect 34808 22642 34836 23122
rect 35072 23044 35124 23050
rect 35072 22986 35124 22992
rect 35084 22930 35112 22986
rect 35084 22902 35388 22930
rect 34796 22636 34848 22642
rect 34796 22578 34848 22584
rect 34808 22098 34836 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 34808 21554 34836 22034
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 20868 34848 20874
rect 34796 20810 34848 20816
rect 34808 20040 34836 20810
rect 35164 20800 35216 20806
rect 35216 20760 35296 20788
rect 35164 20742 35216 20748
rect 35268 20244 35296 20760
rect 35360 20602 35388 22902
rect 35452 22574 35480 24006
rect 35440 22568 35492 22574
rect 35440 22510 35492 22516
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 35348 20596 35400 20602
rect 35348 20538 35400 20544
rect 35268 20216 35388 20244
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20074 35388 20216
rect 35268 20046 35388 20074
rect 34808 20012 35204 20040
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 34808 19553 34836 19790
rect 35176 19786 35204 20012
rect 35268 19922 35296 20046
rect 35348 19984 35400 19990
rect 35348 19926 35400 19932
rect 35452 19938 35480 21558
rect 35544 20398 35572 31726
rect 35900 27328 35952 27334
rect 35900 27270 35952 27276
rect 35714 22808 35770 22817
rect 35714 22743 35770 22752
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 35636 22098 35664 22374
rect 35624 22092 35676 22098
rect 35624 22034 35676 22040
rect 35624 20528 35676 20534
rect 35624 20470 35676 20476
rect 35532 20392 35584 20398
rect 35532 20334 35584 20340
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 35164 19780 35216 19786
rect 35164 19722 35216 19728
rect 34794 19544 34850 19553
rect 34794 19479 34850 19488
rect 34796 19440 34848 19446
rect 35256 19440 35308 19446
rect 34796 19382 34848 19388
rect 34978 19408 35034 19417
rect 34704 18896 34756 18902
rect 34704 18838 34756 18844
rect 34612 18692 34664 18698
rect 34612 18634 34664 18640
rect 34808 18426 34836 19382
rect 35256 19382 35308 19388
rect 34978 19343 35034 19352
rect 34992 19310 35020 19343
rect 34980 19304 35032 19310
rect 34980 19246 35032 19252
rect 35268 19242 35296 19382
rect 35256 19236 35308 19242
rect 35256 19178 35308 19184
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34704 17740 34756 17746
rect 34704 17682 34756 17688
rect 34336 17604 34388 17610
rect 34336 17546 34388 17552
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 34244 14476 34296 14482
rect 34244 14418 34296 14424
rect 34152 14272 34204 14278
rect 34152 14214 34204 14220
rect 34164 13870 34192 14214
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34164 12850 34192 13806
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 34256 12442 34284 14418
rect 34348 14074 34376 17546
rect 34520 15972 34572 15978
rect 34520 15914 34572 15920
rect 34532 15314 34560 15914
rect 34612 15428 34664 15434
rect 34612 15370 34664 15376
rect 34440 15286 34560 15314
rect 34440 15094 34468 15286
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34520 15088 34572 15094
rect 34520 15030 34572 15036
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34532 12918 34560 15030
rect 34520 12912 34572 12918
rect 34520 12854 34572 12860
rect 34244 12436 34296 12442
rect 34244 12378 34296 12384
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 34336 11552 34388 11558
rect 34336 11494 34388 11500
rect 33876 11212 33928 11218
rect 33876 11154 33928 11160
rect 34348 11150 34376 11494
rect 34440 11150 34468 12174
rect 34624 11898 34652 15370
rect 34716 13512 34744 17682
rect 35360 17678 35388 19926
rect 35452 19910 35572 19938
rect 35438 19544 35494 19553
rect 35438 19479 35494 19488
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 34808 15706 34836 17206
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35164 16720 35216 16726
rect 35164 16662 35216 16668
rect 34980 16448 35032 16454
rect 34978 16416 34980 16425
rect 35032 16416 35034 16425
rect 34978 16351 35034 16360
rect 35176 15978 35204 16662
rect 35254 16552 35310 16561
rect 35254 16487 35310 16496
rect 35268 16250 35296 16487
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35164 15972 35216 15978
rect 35164 15914 35216 15920
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 34886 15600 34942 15609
rect 34886 15535 34942 15544
rect 34900 15502 34928 15535
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34886 15192 34942 15201
rect 34886 15127 34942 15136
rect 34900 15026 34928 15127
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34716 13484 35020 13512
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 34888 13184 34940 13190
rect 34888 13126 34940 13132
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34716 11354 34744 12854
rect 34808 12646 34836 13126
rect 34900 12986 34928 13126
rect 34888 12980 34940 12986
rect 34888 12922 34940 12928
rect 34992 12850 35020 13484
rect 35360 12986 35388 17206
rect 35452 16046 35480 19479
rect 35544 16794 35572 19910
rect 35636 18426 35664 20470
rect 35728 19334 35756 22743
rect 35912 21146 35940 27270
rect 36004 26874 36032 35498
rect 36832 35290 36860 35634
rect 36820 35284 36872 35290
rect 36820 35226 36872 35232
rect 37936 35086 37964 36314
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 38198 36136 38254 36145
rect 38028 35290 38056 36110
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38292 35624 38344 35630
rect 38292 35566 38344 35572
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38016 35284 38068 35290
rect 38016 35226 38068 35232
rect 36452 35080 36504 35086
rect 36452 35022 36504 35028
rect 37556 35080 37608 35086
rect 37556 35022 37608 35028
rect 37924 35080 37976 35086
rect 37924 35022 37976 35028
rect 36176 34944 36228 34950
rect 36176 34886 36228 34892
rect 36084 34400 36136 34406
rect 36084 34342 36136 34348
rect 36096 30410 36124 34342
rect 36188 31822 36216 34886
rect 36360 33856 36412 33862
rect 36360 33798 36412 33804
rect 36372 33522 36400 33798
rect 36464 33658 36492 35022
rect 36820 35012 36872 35018
rect 36820 34954 36872 34960
rect 36832 34746 36860 34954
rect 36820 34740 36872 34746
rect 36820 34682 36872 34688
rect 36912 33856 36964 33862
rect 36912 33798 36964 33804
rect 36452 33652 36504 33658
rect 36452 33594 36504 33600
rect 36360 33516 36412 33522
rect 36360 33458 36412 33464
rect 36728 32564 36780 32570
rect 36728 32506 36780 32512
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36176 31816 36228 31822
rect 36280 31793 36308 32370
rect 36452 32360 36504 32366
rect 36452 32302 36504 32308
rect 36176 31758 36228 31764
rect 36266 31784 36322 31793
rect 36266 31719 36322 31728
rect 36096 30382 36216 30410
rect 36084 30252 36136 30258
rect 36084 30194 36136 30200
rect 36096 29073 36124 30194
rect 36082 29064 36138 29073
rect 36082 28999 36138 29008
rect 36188 28082 36216 30382
rect 36360 30184 36412 30190
rect 36360 30126 36412 30132
rect 36176 28076 36228 28082
rect 36176 28018 36228 28024
rect 36004 26846 36308 26874
rect 36176 24268 36228 24274
rect 36176 24210 36228 24216
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35820 19922 35848 20742
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35900 19780 35952 19786
rect 35900 19722 35952 19728
rect 35912 19446 35940 19722
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35728 19306 35848 19334
rect 35716 18896 35768 18902
rect 35716 18838 35768 18844
rect 35624 18420 35676 18426
rect 35624 18362 35676 18368
rect 35728 18290 35756 18838
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35728 17134 35756 17682
rect 35716 17128 35768 17134
rect 35716 17070 35768 17076
rect 35532 16788 35584 16794
rect 35532 16730 35584 16736
rect 35544 16114 35572 16730
rect 35532 16108 35584 16114
rect 35532 16050 35584 16056
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35438 15736 35494 15745
rect 35728 15722 35756 17070
rect 35438 15671 35494 15680
rect 35636 15694 35756 15722
rect 35452 15366 35480 15671
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35636 14958 35664 15694
rect 35716 15632 35768 15638
rect 35716 15574 35768 15580
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35728 14414 35756 15574
rect 35624 14408 35676 14414
rect 35624 14350 35676 14356
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 35532 14000 35584 14006
rect 35532 13942 35584 13948
rect 35440 13864 35492 13870
rect 35440 13806 35492 13812
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 34980 12844 35032 12850
rect 34980 12786 35032 12792
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35452 11898 35480 13806
rect 35544 13530 35572 13942
rect 35532 13524 35584 13530
rect 35532 13466 35584 13472
rect 35532 13388 35584 13394
rect 35532 13330 35584 13336
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34336 11144 34388 11150
rect 34336 11086 34388 11092
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34426 10976 34482 10985
rect 34426 10911 34482 10920
rect 34440 10674 34468 10911
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35544 10198 35572 13330
rect 35636 11626 35664 14350
rect 35728 12442 35756 14350
rect 35820 13326 35848 19306
rect 36004 18873 36032 20878
rect 36096 20602 36124 22714
rect 36188 21350 36216 24210
rect 36176 21344 36228 21350
rect 36176 21286 36228 21292
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 36280 20210 36308 26846
rect 36372 22094 36400 30126
rect 36464 28218 36492 32302
rect 36740 31346 36768 32506
rect 36820 32428 36872 32434
rect 36820 32370 36872 32376
rect 36832 31482 36860 32370
rect 36924 31890 36952 33798
rect 37568 33114 37596 35022
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38016 33312 38068 33318
rect 38016 33254 38068 33260
rect 37556 33108 37608 33114
rect 37556 33050 37608 33056
rect 38028 32910 38056 33254
rect 37832 32904 37884 32910
rect 37832 32846 37884 32852
rect 38016 32904 38068 32910
rect 38016 32846 38068 32852
rect 37844 32230 37872 32846
rect 38120 32745 38148 33458
rect 38200 32768 38252 32774
rect 38106 32736 38162 32745
rect 38200 32710 38252 32716
rect 38106 32671 38162 32680
rect 37832 32224 37884 32230
rect 37832 32166 37884 32172
rect 37004 32020 37056 32026
rect 37004 31962 37056 31968
rect 36912 31884 36964 31890
rect 36912 31826 36964 31832
rect 36912 31680 36964 31686
rect 36912 31622 36964 31628
rect 36820 31476 36872 31482
rect 36820 31418 36872 31424
rect 36728 31340 36780 31346
rect 36728 31282 36780 31288
rect 36636 30592 36688 30598
rect 36636 30534 36688 30540
rect 36648 28966 36676 30534
rect 36740 29646 36768 31282
rect 36728 29640 36780 29646
rect 36728 29582 36780 29588
rect 36636 28960 36688 28966
rect 36636 28902 36688 28908
rect 36452 28212 36504 28218
rect 36452 28154 36504 28160
rect 36636 27328 36688 27334
rect 36636 27270 36688 27276
rect 36648 27130 36676 27270
rect 36636 27124 36688 27130
rect 36636 27066 36688 27072
rect 36544 26308 36596 26314
rect 36544 26250 36596 26256
rect 36452 24608 36504 24614
rect 36452 24550 36504 24556
rect 36464 23730 36492 24550
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36464 23497 36492 23666
rect 36450 23488 36506 23497
rect 36450 23423 36506 23432
rect 36450 22808 36506 22817
rect 36450 22743 36452 22752
rect 36504 22743 36506 22752
rect 36452 22714 36504 22720
rect 36372 22066 36492 22094
rect 36464 20942 36492 22066
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36464 20466 36492 20878
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36280 20182 36400 20210
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 35990 18864 36046 18873
rect 35900 18828 35952 18834
rect 35990 18799 35992 18808
rect 35900 18770 35952 18776
rect 36044 18799 36046 18808
rect 35992 18770 36044 18776
rect 35912 17134 35940 18770
rect 36004 18739 36032 18770
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 35900 17128 35952 17134
rect 35900 17070 35952 17076
rect 35912 16726 35940 17070
rect 35900 16720 35952 16726
rect 35900 16662 35952 16668
rect 35900 16516 35952 16522
rect 35900 16458 35952 16464
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35912 12986 35940 16458
rect 36004 14550 36032 17478
rect 35992 14544 36044 14550
rect 35992 14486 36044 14492
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 35716 12436 35768 12442
rect 35716 12378 35768 12384
rect 35624 11620 35676 11626
rect 35624 11562 35676 11568
rect 36004 10810 36032 13330
rect 36096 12238 36124 19382
rect 36188 19378 36216 19790
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36268 18692 36320 18698
rect 36268 18634 36320 18640
rect 36176 18624 36228 18630
rect 36176 18566 36228 18572
rect 36188 18034 36216 18566
rect 36280 18426 36308 18634
rect 36268 18420 36320 18426
rect 36268 18362 36320 18368
rect 36372 18222 36400 20182
rect 36360 18216 36412 18222
rect 36360 18158 36412 18164
rect 36188 18006 36400 18034
rect 36176 17672 36228 17678
rect 36174 17640 36176 17649
rect 36228 17640 36230 17649
rect 36174 17575 36230 17584
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36280 16998 36308 17478
rect 36268 16992 36320 16998
rect 36268 16934 36320 16940
rect 36268 16652 36320 16658
rect 36268 16594 36320 16600
rect 36176 15972 36228 15978
rect 36176 15914 36228 15920
rect 36188 15162 36216 15914
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 36174 13560 36230 13569
rect 36174 13495 36230 13504
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 35992 10804 36044 10810
rect 35992 10746 36044 10752
rect 36096 10674 36124 11222
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 35532 10192 35584 10198
rect 35532 10134 35584 10140
rect 36188 10062 36216 13495
rect 36280 12986 36308 16594
rect 36372 16096 36400 18006
rect 36464 17542 36492 20402
rect 36452 17536 36504 17542
rect 36452 17478 36504 17484
rect 36450 16280 36506 16289
rect 36450 16215 36452 16224
rect 36504 16215 36506 16224
rect 36452 16186 36504 16192
rect 36452 16108 36504 16114
rect 36372 16068 36452 16096
rect 36452 16050 36504 16056
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36372 14618 36400 15506
rect 36464 15094 36492 16050
rect 36556 15162 36584 26250
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 36636 22976 36688 22982
rect 36636 22918 36688 22924
rect 36648 22234 36676 22918
rect 36636 22228 36688 22234
rect 36636 22170 36688 22176
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 36648 18358 36676 21286
rect 36728 20460 36780 20466
rect 36728 20402 36780 20408
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36648 16153 36676 17478
rect 36634 16144 36690 16153
rect 36634 16079 36690 16088
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36452 15088 36504 15094
rect 36452 15030 36504 15036
rect 36648 15026 36676 16079
rect 36740 15978 36768 20402
rect 36728 15972 36780 15978
rect 36728 15914 36780 15920
rect 36636 15020 36688 15026
rect 36636 14962 36688 14968
rect 36360 14612 36412 14618
rect 36360 14554 36412 14560
rect 36372 13530 36400 14554
rect 36452 14000 36504 14006
rect 36452 13942 36504 13948
rect 36360 13524 36412 13530
rect 36360 13466 36412 13472
rect 36360 13388 36412 13394
rect 36360 13330 36412 13336
rect 36268 12980 36320 12986
rect 36268 12922 36320 12928
rect 36372 12481 36400 13330
rect 36358 12472 36414 12481
rect 36358 12407 36414 12416
rect 36266 12336 36322 12345
rect 36266 12271 36322 12280
rect 36280 11830 36308 12271
rect 36268 11824 36320 11830
rect 36268 11766 36320 11772
rect 36360 11824 36412 11830
rect 36360 11766 36412 11772
rect 36266 11656 36322 11665
rect 36266 11591 36322 11600
rect 36280 11354 36308 11591
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 36372 10742 36400 11766
rect 36360 10736 36412 10742
rect 36360 10678 36412 10684
rect 36176 10056 36228 10062
rect 36176 9998 36228 10004
rect 35992 9920 36044 9926
rect 35992 9862 36044 9868
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 33784 3732 33836 3738
rect 33784 3674 33836 3680
rect 34440 2922 34468 7142
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35348 4480 35400 4486
rect 35348 4422 35400 4428
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34520 3460 34572 3466
rect 34520 3402 34572 3408
rect 34428 2916 34480 2922
rect 34428 2858 34480 2864
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 32324 2446 32352 2790
rect 34532 2650 34560 3402
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 35360 2378 35388 4422
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 35348 2372 35400 2378
rect 35348 2314 35400 2320
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 30300 800 30328 2246
rect 30944 800 30972 2246
rect 32232 800 32260 2246
rect 33520 800 33548 2246
rect 34164 800 34192 2314
rect 35452 800 35480 2926
rect 35898 2680 35954 2689
rect 35898 2615 35954 2624
rect 35912 2446 35940 2615
rect 36004 2514 36032 9862
rect 36464 9654 36492 13942
rect 36636 13932 36688 13938
rect 36636 13874 36688 13880
rect 36544 12640 36596 12646
rect 36544 12582 36596 12588
rect 36556 12238 36584 12582
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36556 11830 36584 12174
rect 36544 11824 36596 11830
rect 36544 11766 36596 11772
rect 36556 11150 36584 11766
rect 36544 11144 36596 11150
rect 36544 11086 36596 11092
rect 36648 10062 36676 13874
rect 36832 12782 36860 25638
rect 36924 25294 36952 31622
rect 37016 30258 37044 31962
rect 37464 31272 37516 31278
rect 37464 31214 37516 31220
rect 37476 30802 37504 31214
rect 37844 30938 37872 32166
rect 38212 32065 38240 32710
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38304 31822 38332 35566
rect 38672 34542 38700 39200
rect 39316 35290 39344 39200
rect 39672 37256 39724 37262
rect 39672 37198 39724 37204
rect 39684 35894 39712 37198
rect 39684 35866 39896 35894
rect 39304 35284 39356 35290
rect 39304 35226 39356 35232
rect 39028 34604 39080 34610
rect 39028 34546 39080 34552
rect 38660 34536 38712 34542
rect 38660 34478 38712 34484
rect 38844 33380 38896 33386
rect 38844 33322 38896 33328
rect 38568 32836 38620 32842
rect 38568 32778 38620 32784
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 37832 30932 37884 30938
rect 37832 30874 37884 30880
rect 38384 30864 38436 30870
rect 38384 30806 38436 30812
rect 37464 30796 37516 30802
rect 37464 30738 37516 30744
rect 37556 30728 37608 30734
rect 37556 30670 37608 30676
rect 38198 30696 38254 30705
rect 37004 30252 37056 30258
rect 37004 30194 37056 30200
rect 37568 28762 37596 30670
rect 38198 30631 38254 30640
rect 38212 30394 38240 30631
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37648 29504 37700 29510
rect 37648 29446 37700 29452
rect 37556 28756 37608 28762
rect 37556 28698 37608 28704
rect 37660 28558 37688 29446
rect 37648 28552 37700 28558
rect 37648 28494 37700 28500
rect 37556 27396 37608 27402
rect 37556 27338 37608 27344
rect 37004 26240 37056 26246
rect 37004 26182 37056 26188
rect 37016 25498 37044 26182
rect 37096 25968 37148 25974
rect 37096 25910 37148 25916
rect 37004 25492 37056 25498
rect 37004 25434 37056 25440
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 36912 23860 36964 23866
rect 36912 23802 36964 23808
rect 36924 18970 36952 23802
rect 37004 23044 37056 23050
rect 37004 22986 37056 22992
rect 37016 22234 37044 22986
rect 37004 22228 37056 22234
rect 37004 22170 37056 22176
rect 37004 21956 37056 21962
rect 37004 21898 37056 21904
rect 37016 21418 37044 21898
rect 37004 21412 37056 21418
rect 37004 21354 37056 21360
rect 36912 18964 36964 18970
rect 36912 18906 36964 18912
rect 36910 17096 36966 17105
rect 36910 17031 36966 17040
rect 36820 12776 36872 12782
rect 36820 12718 36872 12724
rect 36728 12640 36780 12646
rect 36728 12582 36780 12588
rect 36740 11558 36768 12582
rect 36924 11558 36952 17031
rect 37004 14816 37056 14822
rect 37004 14758 37056 14764
rect 37016 12186 37044 14758
rect 37108 12442 37136 25910
rect 37464 24200 37516 24206
rect 37464 24142 37516 24148
rect 37476 23905 37504 24142
rect 37462 23896 37518 23905
rect 37568 23866 37596 27338
rect 37648 27328 37700 27334
rect 37648 27270 37700 27276
rect 37660 25809 37688 27270
rect 37646 25800 37702 25809
rect 37646 25735 37702 25744
rect 37462 23831 37518 23840
rect 37556 23860 37608 23866
rect 37556 23802 37608 23808
rect 37648 23792 37700 23798
rect 37648 23734 37700 23740
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37280 22976 37332 22982
rect 37280 22918 37332 22924
rect 37188 22704 37240 22710
rect 37188 22646 37240 22652
rect 37200 17746 37228 22646
rect 37292 21622 37320 22918
rect 37476 22030 37504 23054
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37292 21146 37320 21422
rect 37476 21146 37504 21966
rect 37280 21140 37332 21146
rect 37280 21082 37332 21088
rect 37464 21140 37516 21146
rect 37464 21082 37516 21088
rect 37278 21040 37334 21049
rect 37278 20975 37334 20984
rect 37464 21004 37516 21010
rect 37188 17740 37240 17746
rect 37188 17682 37240 17688
rect 37292 17678 37320 20975
rect 37464 20946 37516 20952
rect 37372 20868 37424 20874
rect 37372 20810 37424 20816
rect 37384 17882 37412 20810
rect 37476 19990 37504 20946
rect 37464 19984 37516 19990
rect 37464 19926 37516 19932
rect 37464 19304 37516 19310
rect 37464 19246 37516 19252
rect 37476 19145 37504 19246
rect 37462 19136 37518 19145
rect 37462 19071 37518 19080
rect 37462 19000 37518 19009
rect 37462 18935 37518 18944
rect 37476 18306 37504 18935
rect 37568 18426 37596 22578
rect 37660 18970 37688 23734
rect 37844 22001 37872 29582
rect 37924 29572 37976 29578
rect 37924 29514 37976 29520
rect 37830 21992 37886 22001
rect 37830 21927 37886 21936
rect 37832 21888 37884 21894
rect 37832 21830 37884 21836
rect 37740 21412 37792 21418
rect 37740 21354 37792 21360
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37556 18420 37608 18426
rect 37556 18362 37608 18368
rect 37476 18278 37596 18306
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37476 18086 37504 18158
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37476 17678 37504 18022
rect 37280 17672 37332 17678
rect 37280 17614 37332 17620
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 17264 37424 17270
rect 37372 17206 37424 17212
rect 37188 14952 37240 14958
rect 37188 14894 37240 14900
rect 37200 13326 37228 14894
rect 37188 13320 37240 13326
rect 37188 13262 37240 13268
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37292 12866 37320 12922
rect 37200 12838 37320 12866
rect 37096 12436 37148 12442
rect 37096 12378 37148 12384
rect 37016 12170 37136 12186
rect 37016 12164 37148 12170
rect 37016 12158 37096 12164
rect 37096 12106 37148 12112
rect 37200 11898 37228 12838
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 37188 11892 37240 11898
rect 37188 11834 37240 11840
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 36726 10568 36782 10577
rect 36726 10503 36782 10512
rect 36740 10266 36768 10503
rect 36728 10260 36780 10266
rect 36728 10202 36780 10208
rect 36636 10056 36688 10062
rect 36636 9998 36688 10004
rect 37292 9654 37320 12718
rect 37384 10810 37412 17206
rect 37476 16658 37504 17614
rect 37568 17134 37596 18278
rect 37648 18284 37700 18290
rect 37648 18226 37700 18232
rect 37660 17814 37688 18226
rect 37752 17882 37780 21354
rect 37740 17876 37792 17882
rect 37740 17818 37792 17824
rect 37648 17808 37700 17814
rect 37648 17750 37700 17756
rect 37844 17610 37872 21830
rect 37832 17604 37884 17610
rect 37832 17546 37884 17552
rect 37556 17128 37608 17134
rect 37556 17070 37608 17076
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37476 12646 37504 15438
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37462 12472 37518 12481
rect 37462 12407 37518 12416
rect 37372 10804 37424 10810
rect 37372 10746 37424 10752
rect 37476 10674 37504 12407
rect 37568 12306 37596 17070
rect 37936 16522 37964 29514
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38212 29345 38240 29446
rect 38198 29336 38254 29345
rect 38198 29271 38254 29280
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38028 20466 38056 28358
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38200 26784 38252 26790
rect 38200 26726 38252 26732
rect 38212 26314 38240 26726
rect 38200 26308 38252 26314
rect 38200 26250 38252 26256
rect 38290 25936 38346 25945
rect 38290 25871 38292 25880
rect 38344 25871 38346 25880
rect 38292 25842 38344 25848
rect 38198 25256 38254 25265
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38292 24812 38344 24818
rect 38292 24754 38344 24760
rect 38108 24200 38160 24206
rect 38108 24142 38160 24148
rect 38120 21010 38148 24142
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38304 22094 38332 24754
rect 38212 22066 38332 22094
rect 38108 21004 38160 21010
rect 38108 20946 38160 20952
rect 38212 20754 38240 22066
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38292 21344 38344 21350
rect 38292 21286 38344 21292
rect 38120 20726 38240 20754
rect 38016 20460 38068 20466
rect 38016 20402 38068 20408
rect 38016 18760 38068 18766
rect 38016 18702 38068 18708
rect 38028 18222 38056 18702
rect 38016 18216 38068 18222
rect 38016 18158 38068 18164
rect 37924 16516 37976 16522
rect 37924 16458 37976 16464
rect 37740 16176 37792 16182
rect 37740 16118 37792 16124
rect 37648 16040 37700 16046
rect 37648 15982 37700 15988
rect 37556 12300 37608 12306
rect 37556 12242 37608 12248
rect 37554 11928 37610 11937
rect 37554 11863 37556 11872
rect 37608 11863 37610 11872
rect 37556 11834 37608 11840
rect 37556 11756 37608 11762
rect 37556 11698 37608 11704
rect 37568 11626 37596 11698
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37464 10668 37516 10674
rect 37464 10610 37516 10616
rect 37568 10062 37596 11562
rect 37660 11218 37688 15982
rect 37648 11212 37700 11218
rect 37648 11154 37700 11160
rect 37752 11082 37780 16118
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 37924 15428 37976 15434
rect 37924 15370 37976 15376
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37740 11076 37792 11082
rect 37740 11018 37792 11024
rect 37740 10532 37792 10538
rect 37740 10474 37792 10480
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 36452 9648 36504 9654
rect 36452 9590 36504 9596
rect 37280 9648 37332 9654
rect 37280 9590 37332 9596
rect 36464 4146 36492 9590
rect 37752 9586 37780 10474
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 37844 9450 37872 13262
rect 37936 12986 37964 15370
rect 38028 15337 38056 15438
rect 38014 15328 38070 15337
rect 38014 15263 38070 15272
rect 38120 15162 38148 20726
rect 38200 20596 38252 20602
rect 38200 20538 38252 20544
rect 38212 20505 38240 20538
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 38198 20360 38254 20369
rect 38198 20295 38254 20304
rect 38212 15910 38240 20295
rect 38304 17241 38332 21286
rect 38290 17232 38346 17241
rect 38290 17167 38346 17176
rect 38292 17128 38344 17134
rect 38292 17070 38344 17076
rect 38304 16046 38332 17070
rect 38292 16040 38344 16046
rect 38292 15982 38344 15988
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38108 15156 38160 15162
rect 38108 15098 38160 15104
rect 38212 15065 38240 15302
rect 38198 15056 38254 15065
rect 38108 15020 38160 15026
rect 38198 14991 38254 15000
rect 38108 14962 38160 14968
rect 38120 14414 38148 14962
rect 38108 14408 38160 14414
rect 38108 14350 38160 14356
rect 38120 13938 38148 14350
rect 38108 13932 38160 13938
rect 38108 13874 38160 13880
rect 38016 13184 38068 13190
rect 38016 13126 38068 13132
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 37924 12980 37976 12986
rect 37924 12922 37976 12928
rect 37936 12782 37964 12922
rect 37924 12776 37976 12782
rect 37924 12718 37976 12724
rect 37832 9444 37884 9450
rect 37832 9386 37884 9392
rect 38028 8974 38056 13126
rect 38108 12708 38160 12714
rect 38108 12650 38160 12656
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38120 8634 38148 12650
rect 38212 12345 38240 13126
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38304 11778 38332 15982
rect 38396 12434 38424 30806
rect 38476 26444 38528 26450
rect 38476 26386 38528 26392
rect 38488 17270 38516 26386
rect 38476 17264 38528 17270
rect 38476 17206 38528 17212
rect 38580 14074 38608 32778
rect 38660 28484 38712 28490
rect 38660 28426 38712 28432
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38672 14006 38700 28426
rect 38752 21004 38804 21010
rect 38752 20946 38804 20952
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 38396 12406 38516 12434
rect 38384 12368 38436 12374
rect 38384 12310 38436 12316
rect 38212 11762 38332 11778
rect 38200 11756 38332 11762
rect 38252 11750 38332 11756
rect 38200 11698 38252 11704
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38212 10305 38240 10406
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 38304 8498 38332 10911
rect 38396 10606 38424 12310
rect 38488 10742 38516 12406
rect 38764 12102 38792 20946
rect 38856 17354 38884 33322
rect 38936 26512 38988 26518
rect 38936 26454 38988 26460
rect 38948 18902 38976 26454
rect 38936 18896 38988 18902
rect 38936 18838 38988 18844
rect 38856 17326 38976 17354
rect 38844 17264 38896 17270
rect 38844 17206 38896 17212
rect 38856 12374 38884 17206
rect 38948 15201 38976 17326
rect 39040 15706 39068 34546
rect 39396 31816 39448 31822
rect 39396 31758 39448 31764
rect 39212 30660 39264 30666
rect 39212 30602 39264 30608
rect 39120 29164 39172 29170
rect 39120 29106 39172 29112
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 38934 15192 38990 15201
rect 38934 15127 38990 15136
rect 39132 12442 39160 29106
rect 39224 13530 39252 30602
rect 39304 25696 39356 25702
rect 39304 25638 39356 25644
rect 39316 14482 39344 25638
rect 39408 19922 39436 31758
rect 39868 31754 39896 35866
rect 39684 31726 39896 31754
rect 39488 24132 39540 24138
rect 39488 24074 39540 24080
rect 39396 19916 39448 19922
rect 39396 19858 39448 19864
rect 39500 16454 39528 24074
rect 39684 21350 39712 31726
rect 39764 23724 39816 23730
rect 39764 23666 39816 23672
rect 39672 21344 39724 21350
rect 39672 21286 39724 21292
rect 39672 21208 39724 21214
rect 39672 21150 39724 21156
rect 39580 21140 39632 21146
rect 39580 21082 39632 21088
rect 39592 18766 39620 21082
rect 39580 18760 39632 18766
rect 39580 18702 39632 18708
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 39304 14476 39356 14482
rect 39304 14418 39356 14424
rect 39212 13524 39264 13530
rect 39212 13466 39264 13472
rect 39120 12436 39172 12442
rect 39120 12378 39172 12384
rect 38844 12368 38896 12374
rect 38844 12310 38896 12316
rect 38752 12096 38804 12102
rect 38752 12038 38804 12044
rect 38476 10736 38528 10742
rect 38476 10678 38528 10684
rect 38384 10600 38436 10606
rect 38384 10542 38436 10548
rect 38764 8566 38792 12038
rect 39684 9586 39712 21150
rect 39776 15026 39804 23666
rect 39856 22160 39908 22166
rect 39856 22102 39908 22108
rect 39764 15020 39816 15026
rect 39764 14962 39816 14968
rect 39868 14618 39896 22102
rect 39856 14612 39908 14618
rect 39856 14554 39908 14560
rect 39672 9580 39724 9586
rect 39672 9522 39724 9528
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 36636 8356 36688 8362
rect 36636 8298 36688 8304
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 35992 2508 36044 2514
rect 35992 2450 36044 2456
rect 36648 2446 36676 8298
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38212 7585 38240 7686
rect 38198 7576 38254 7585
rect 38198 7511 38254 7520
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4185 38332 4558
rect 38290 4176 38346 4185
rect 38016 4140 38068 4146
rect 38290 4111 38346 4120
rect 38016 4082 38068 4088
rect 36912 3936 36964 3942
rect 36912 3878 36964 3884
rect 36924 3058 36952 3878
rect 37464 3528 37516 3534
rect 37462 3496 37464 3505
rect 37516 3496 37518 3505
rect 37462 3431 37518 3440
rect 38028 3194 38056 4082
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 37188 2576 37240 2582
rect 37188 2518 37240 2524
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 36636 2440 36688 2446
rect 36636 2382 36688 2388
rect 36820 2304 36872 2310
rect 36820 2246 36872 2252
rect 37004 2304 37056 2310
rect 37004 2246 37056 2252
rect 36832 2145 36860 2246
rect 36818 2136 36874 2145
rect 36818 2071 36874 2080
rect 36740 870 36860 898
rect 36740 800 36768 870
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 36832 762 36860 870
rect 37016 762 37044 2246
rect 36832 734 37044 762
rect 37200 105 37228 2518
rect 37384 800 37412 2790
rect 37370 200 37426 800
rect 38212 785 38240 3878
rect 38660 3460 38712 3466
rect 38660 3402 38712 3408
rect 38672 800 38700 3402
rect 38198 776 38254 785
rect 38198 711 38254 720
rect 38658 200 38714 800
rect 37186 96 37242 105
rect 37186 31 37242 40
<< via2 >>
rect 1582 38800 1638 38856
rect 1674 36896 1730 36952
rect 1766 36116 1768 36136
rect 1768 36116 1820 36136
rect 1820 36116 1822 36136
rect 1766 36080 1822 36116
rect 1674 35708 1676 35728
rect 1676 35708 1728 35728
rect 1728 35708 1730 35728
rect 1674 35672 1730 35708
rect 1766 34040 1822 34096
rect 1766 32716 1768 32736
rect 1768 32716 1820 32736
rect 1820 32716 1822 32736
rect 1766 32680 1822 32716
rect 1766 32000 1822 32056
rect 1766 30640 1822 30696
rect 1766 29280 1822 29336
rect 1766 28600 1822 28656
rect 1766 27240 1822 27296
rect 1766 25880 1822 25936
rect 1766 24556 1768 24576
rect 1768 24556 1820 24576
rect 1820 24556 1822 24576
rect 1766 24520 1822 24556
rect 1766 23840 1822 23896
rect 1674 22480 1730 22536
rect 1766 21120 1822 21176
rect 1766 20440 1822 20496
rect 3422 39480 3478 39536
rect 2870 37440 2926 37496
rect 2410 35536 2466 35592
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1582 19080 1638 19136
rect 1582 17076 1584 17096
rect 1584 17076 1636 17096
rect 1636 17076 1638 17096
rect 1582 17040 1638 17076
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 6458 36216 6514 36272
rect 7010 36780 7066 36816
rect 7010 36760 7012 36780
rect 7012 36760 7064 36780
rect 7064 36760 7066 36780
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 10506 37304 10562 37360
rect 8574 36644 8630 36680
rect 8574 36624 8576 36644
rect 8576 36624 8628 36644
rect 8628 36624 8630 36644
rect 9034 36488 9090 36544
rect 8298 32408 8354 32464
rect 8206 31320 8262 31376
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 9310 34448 9366 34504
rect 10138 36524 10140 36544
rect 10140 36524 10192 36544
rect 10192 36524 10194 36544
rect 10138 36488 10194 36524
rect 10138 35400 10194 35456
rect 11702 37204 11704 37224
rect 11704 37204 11756 37224
rect 11756 37204 11758 37224
rect 11702 37168 11758 37204
rect 10322 35944 10378 36000
rect 10598 35808 10654 35864
rect 11058 36080 11114 36136
rect 10874 35264 10930 35320
rect 11242 35944 11298 36000
rect 10966 35128 11022 35184
rect 10690 34620 10692 34640
rect 10692 34620 10744 34640
rect 10744 34620 10746 34640
rect 10690 34584 10746 34620
rect 10138 32952 10194 33008
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1766 17720 1822 17776
rect 1766 15680 1822 15736
rect 1766 14320 1822 14376
rect 1766 13640 1822 13696
rect 1766 12280 1822 12336
rect 1766 10920 1822 10976
rect 1766 10240 1822 10296
rect 1766 8916 1768 8936
rect 1768 8916 1820 8936
rect 1820 8916 1822 8936
rect 1766 8880 1822 8916
rect 1766 7520 1822 7576
rect 1582 6840 1638 6896
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1582 5480 1638 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1766 4120 1822 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1766 3440 1822 3496
rect 3146 2080 3202 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10782 33360 10838 33416
rect 10506 28756 10562 28792
rect 10506 28736 10508 28756
rect 10508 28736 10560 28756
rect 10560 28736 10562 28756
rect 11058 33224 11114 33280
rect 11058 31204 11114 31240
rect 11058 31184 11060 31204
rect 11060 31184 11112 31204
rect 11112 31184 11114 31204
rect 11794 36896 11850 36952
rect 11886 36488 11942 36544
rect 12070 36488 12126 36544
rect 12162 35808 12218 35864
rect 11886 34620 11888 34640
rect 11888 34620 11940 34640
rect 11940 34620 11942 34640
rect 11886 34584 11942 34620
rect 11978 33768 12034 33824
rect 11702 33088 11758 33144
rect 10874 29824 10930 29880
rect 10966 29008 11022 29064
rect 11518 21528 11574 21584
rect 13174 35264 13230 35320
rect 12898 34076 12900 34096
rect 12900 34076 12952 34096
rect 12952 34076 12954 34096
rect 12898 34040 12954 34076
rect 13634 35284 13690 35320
rect 13634 35264 13636 35284
rect 13636 35264 13688 35284
rect 13688 35264 13690 35284
rect 13174 33632 13230 33688
rect 14370 33904 14426 33960
rect 15106 34448 15162 34504
rect 15106 33496 15162 33552
rect 12806 31320 12862 31376
rect 13542 32272 13598 32328
rect 13542 31084 13544 31104
rect 13544 31084 13596 31104
rect 13596 31084 13598 31104
rect 13542 31048 13598 31084
rect 13174 30252 13230 30288
rect 13174 30232 13176 30252
rect 13176 30232 13228 30252
rect 13228 30232 13230 30252
rect 12806 29280 12862 29336
rect 13634 29552 13690 29608
rect 14462 32836 14518 32872
rect 14462 32816 14464 32836
rect 14464 32816 14516 32836
rect 14516 32816 14518 32836
rect 13082 27784 13138 27840
rect 13634 25336 13690 25392
rect 14370 30368 14426 30424
rect 15290 36896 15346 36952
rect 16302 36488 16358 36544
rect 15566 34584 15622 34640
rect 15566 34196 15622 34232
rect 15566 34176 15568 34196
rect 15568 34176 15620 34196
rect 15620 34176 15622 34196
rect 15566 33632 15622 33688
rect 15750 31728 15806 31784
rect 15106 29008 15162 29064
rect 14922 28500 14924 28520
rect 14924 28500 14976 28520
rect 14976 28500 14978 28520
rect 14922 28464 14978 28500
rect 17038 37168 17094 37224
rect 16670 34196 16726 34232
rect 16670 34176 16672 34196
rect 16672 34176 16724 34196
rect 16724 34176 16726 34196
rect 17038 36488 17094 36544
rect 15842 27784 15898 27840
rect 14922 20440 14978 20496
rect 17038 34040 17094 34096
rect 17590 33632 17646 33688
rect 17038 31048 17094 31104
rect 16854 21936 16910 21992
rect 18326 37304 18382 37360
rect 17958 35284 18014 35320
rect 17958 35264 17960 35284
rect 17960 35264 18012 35284
rect 18012 35264 18014 35284
rect 18602 33224 18658 33280
rect 18510 31320 18566 31376
rect 17682 28872 17738 28928
rect 17866 28872 17922 28928
rect 17958 28736 18014 28792
rect 17682 28484 17738 28520
rect 17682 28464 17684 28484
rect 17684 28464 17736 28484
rect 17736 28464 17738 28484
rect 19430 37304 19486 37360
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 18786 33088 18842 33144
rect 18878 32952 18934 33008
rect 19062 31864 19118 31920
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19338 33768 19394 33824
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19890 33380 19946 33416
rect 19890 33360 19892 33380
rect 19892 33360 19944 33380
rect 19944 33360 19946 33380
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19982 32272 20038 32328
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19798 30268 19800 30288
rect 19800 30268 19852 30288
rect 19852 30268 19854 30288
rect 19798 30232 19854 30268
rect 18878 30096 18934 30152
rect 19062 29844 19118 29880
rect 19062 29824 19064 29844
rect 19064 29824 19116 29844
rect 19116 29824 19118 29844
rect 19798 29844 19854 29880
rect 19798 29824 19800 29844
rect 19800 29824 19852 29844
rect 19852 29824 19854 29844
rect 19338 29552 19394 29608
rect 19430 29416 19486 29472
rect 18970 29280 19026 29336
rect 19246 29280 19302 29336
rect 18418 29008 18474 29064
rect 18602 24112 18658 24168
rect 19338 29144 19394 29200
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 20626 36080 20682 36136
rect 20166 31748 20222 31784
rect 20166 31728 20168 31748
rect 20168 31728 20220 31748
rect 20220 31728 20222 31748
rect 20166 30132 20168 30152
rect 20168 30132 20220 30152
rect 20220 30132 20222 30152
rect 20166 30096 20222 30132
rect 20166 29688 20222 29744
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19706 25220 19762 25256
rect 19706 25200 19708 25220
rect 19708 25200 19760 25220
rect 19760 25200 19762 25220
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 18970 18128 19026 18184
rect 19614 24268 19670 24304
rect 19614 24248 19616 24268
rect 19616 24248 19668 24268
rect 19668 24248 19670 24268
rect 19522 24112 19578 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19338 22344 19394 22400
rect 18510 14320 18566 14376
rect 20350 32428 20406 32464
rect 20350 32408 20352 32428
rect 20352 32408 20404 32428
rect 20404 32408 20406 32428
rect 20902 36488 20958 36544
rect 21178 36488 21234 36544
rect 20350 29144 20406 29200
rect 20718 33904 20774 33960
rect 20718 29552 20774 29608
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20074 22772 20130 22808
rect 20074 22752 20076 22772
rect 20076 22752 20128 22772
rect 20128 22752 20130 22772
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20258 22752 20314 22808
rect 20994 31864 21050 31920
rect 22742 36488 22798 36544
rect 23018 35400 23074 35456
rect 20994 25336 21050 25392
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20626 19896 20682 19952
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20902 21936 20958 21992
rect 21270 20576 21326 20632
rect 20810 16768 20866 16824
rect 20626 16088 20682 16144
rect 26330 37304 26386 37360
rect 24858 36488 24914 36544
rect 24582 32816 24638 32872
rect 24582 30368 24638 30424
rect 25042 30232 25098 30288
rect 22742 21800 22798 21856
rect 22650 20868 22706 20904
rect 22650 20848 22652 20868
rect 22652 20848 22704 20868
rect 22704 20848 22706 20868
rect 21730 20052 21786 20088
rect 21730 20032 21732 20052
rect 21732 20032 21784 20052
rect 21784 20032 21786 20052
rect 25870 37168 25926 37224
rect 25594 33532 25596 33552
rect 25596 33532 25648 33552
rect 25648 33532 25650 33552
rect 25594 33496 25650 33532
rect 25502 32272 25558 32328
rect 23570 18264 23626 18320
rect 23294 17720 23350 17776
rect 22650 16124 22652 16144
rect 22652 16124 22704 16144
rect 22704 16124 22706 16144
rect 22650 16088 22706 16124
rect 22650 15988 22652 16008
rect 22652 15988 22704 16008
rect 22704 15988 22706 16008
rect 22650 15952 22706 15988
rect 24858 24268 24914 24304
rect 24858 24248 24860 24268
rect 24860 24248 24912 24268
rect 24912 24248 24914 24268
rect 24766 18808 24822 18864
rect 25226 21936 25282 21992
rect 25042 20984 25098 21040
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 25778 32000 25834 32056
rect 25778 20848 25834 20904
rect 25226 16904 25282 16960
rect 26330 21936 26386 21992
rect 26054 18808 26110 18864
rect 27434 35572 27436 35592
rect 27436 35572 27488 35592
rect 27488 35572 27490 35592
rect 27434 35536 27490 35572
rect 27618 33224 27674 33280
rect 27802 31184 27858 31240
rect 26698 20848 26754 20904
rect 26606 20576 26662 20632
rect 26698 19488 26754 19544
rect 26514 15272 26570 15328
rect 27618 23432 27674 23488
rect 27066 20884 27068 20904
rect 27068 20884 27120 20904
rect 27120 20884 27122 20904
rect 27066 20848 27122 20884
rect 27158 20032 27214 20088
rect 27066 17040 27122 17096
rect 27618 21528 27674 21584
rect 27710 20712 27766 20768
rect 27250 17332 27306 17368
rect 27250 17312 27252 17332
rect 27252 17312 27304 17332
rect 27304 17312 27306 17332
rect 27526 18264 27582 18320
rect 29918 36352 29974 36408
rect 30010 36216 30066 36272
rect 28998 35944 29054 36000
rect 30746 36352 30802 36408
rect 28446 35128 28502 35184
rect 28262 26152 28318 26208
rect 27986 19488 28042 19544
rect 28630 30368 28686 30424
rect 28446 21004 28502 21040
rect 28446 20984 28448 21004
rect 28448 20984 28500 21004
rect 28500 20984 28502 21004
rect 27986 15952 28042 16008
rect 28538 17720 28594 17776
rect 28906 25200 28962 25256
rect 28538 17076 28540 17096
rect 28540 17076 28592 17096
rect 28592 17076 28594 17096
rect 28538 17040 28594 17076
rect 29182 17720 29238 17776
rect 30470 35692 30526 35728
rect 30470 35672 30472 35692
rect 30472 35672 30524 35692
rect 30524 35672 30526 35692
rect 30562 30368 30618 30424
rect 32310 36352 32366 36408
rect 33138 36488 33194 36544
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35162 37324 35218 37360
rect 35162 37304 35164 37324
rect 35164 37304 35216 37324
rect 35216 37304 35218 37324
rect 31850 33768 31906 33824
rect 32034 30368 32090 30424
rect 31666 29996 31668 30016
rect 31668 29996 31720 30016
rect 31720 29996 31722 30016
rect 31666 29960 31722 29996
rect 31298 29008 31354 29064
rect 32218 29008 32274 29064
rect 29550 19080 29606 19136
rect 29458 17620 29460 17640
rect 29460 17620 29512 17640
rect 29512 17620 29514 17640
rect 29458 17584 29514 17620
rect 30378 18536 30434 18592
rect 30378 17856 30434 17912
rect 30746 24928 30802 24984
rect 31206 23024 31262 23080
rect 30746 20440 30802 20496
rect 31206 18944 31262 19000
rect 30930 18672 30986 18728
rect 30746 15952 30802 16008
rect 31022 17584 31078 17640
rect 30930 16768 30986 16824
rect 31114 16532 31116 16552
rect 31116 16532 31168 16552
rect 31168 16532 31170 16552
rect 31114 16496 31170 16532
rect 31022 16088 31078 16144
rect 30930 15680 30986 15736
rect 31574 18808 31630 18864
rect 31850 22752 31906 22808
rect 32678 23024 32734 23080
rect 32586 20576 32642 20632
rect 31758 16904 31814 16960
rect 32310 19488 32366 19544
rect 32402 18944 32458 19000
rect 32586 18692 32642 18728
rect 32586 18672 32588 18692
rect 32588 18672 32640 18692
rect 32640 18672 32642 18692
rect 33230 29180 33232 29200
rect 33232 29180 33284 29200
rect 33284 29180 33286 29200
rect 33230 29144 33286 29180
rect 32954 20984 33010 21040
rect 32954 18128 33010 18184
rect 33046 17720 33102 17776
rect 32494 13368 32550 13424
rect 32862 13524 32918 13560
rect 32862 13504 32864 13524
rect 32864 13504 32916 13524
rect 32916 13504 32918 13524
rect 33046 15272 33102 15328
rect 33230 18536 33286 18592
rect 33230 16768 33286 16824
rect 33322 16632 33378 16688
rect 33690 24928 33746 24984
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 37186 37440 37242 37496
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34610 30932 34666 30968
rect 34610 30912 34612 30932
rect 34612 30912 34664 30932
rect 34664 30912 34666 30932
rect 33874 19916 33930 19952
rect 33874 19896 33876 19916
rect 33876 19896 33928 19916
rect 33928 19896 33930 19916
rect 33690 19216 33746 19272
rect 33506 15952 33562 16008
rect 33138 13232 33194 13288
rect 33414 12280 33470 12336
rect 33690 13640 33746 13696
rect 33690 12708 33746 12744
rect 33690 12688 33692 12708
rect 33692 12688 33744 12708
rect 33744 12688 33746 12708
rect 34426 26288 34482 26344
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 36174 36624 36230 36680
rect 37462 38800 37518 38856
rect 37554 36760 37610 36816
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35530 33360 35586 33416
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35714 22752 35770 22808
rect 34794 19488 34850 19544
rect 34978 19352 35034 19408
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35438 19488 35494 19544
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34978 16396 34980 16416
rect 34980 16396 35032 16416
rect 35032 16396 35034 16416
rect 34978 16360 35034 16396
rect 35254 16496 35310 16552
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34886 15544 34942 15600
rect 34886 15136 34942 15192
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 36266 31728 36322 31784
rect 36082 29008 36138 29064
rect 35438 15680 35494 15736
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34426 10920 34482 10976
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38198 34040 38254 34096
rect 38106 32680 38162 32736
rect 36450 23432 36506 23488
rect 36450 22772 36506 22808
rect 36450 22752 36452 22772
rect 36452 22752 36504 22772
rect 36504 22752 36506 22772
rect 35990 18828 36046 18864
rect 35990 18808 35992 18828
rect 35992 18808 36044 18828
rect 36044 18808 36046 18828
rect 36174 17620 36176 17640
rect 36176 17620 36228 17640
rect 36228 17620 36230 17640
rect 36174 17584 36230 17620
rect 36174 13504 36230 13560
rect 36450 16244 36506 16280
rect 36450 16224 36452 16244
rect 36452 16224 36504 16244
rect 36504 16224 36506 16244
rect 36634 16088 36690 16144
rect 36358 12416 36414 12472
rect 36266 12280 36322 12336
rect 36266 11600 36322 11656
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 2624 35954 2680
rect 38198 32000 38254 32056
rect 38198 30640 38254 30696
rect 36910 17040 36966 17096
rect 37462 23840 37518 23896
rect 37646 25744 37702 25800
rect 37278 20984 37334 21040
rect 37462 19080 37518 19136
rect 37462 18944 37518 19000
rect 37830 21936 37886 21992
rect 36726 10512 36782 10568
rect 37462 12416 37518 12472
rect 38198 29280 38254 29336
rect 38198 28600 38254 28656
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25900 38346 25936
rect 38290 25880 38292 25900
rect 38292 25880 38344 25900
rect 38344 25880 38346 25900
rect 38198 25200 38254 25256
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38290 21800 38346 21856
rect 37554 11892 37610 11928
rect 37554 11872 37556 11892
rect 37556 11872 37608 11892
rect 37608 11872 37610 11892
rect 38014 15272 38070 15328
rect 38198 20440 38254 20496
rect 38198 20304 38254 20360
rect 38290 17176 38346 17232
rect 38198 15000 38254 15056
rect 38198 12280 38254 12336
rect 38290 10920 38346 10976
rect 38198 10240 38254 10296
rect 38198 8880 38254 8936
rect 38934 15136 38990 15192
rect 38198 7520 38254 7576
rect 38290 6840 38346 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 38290 4120 38346 4176
rect 37462 3476 37464 3496
rect 37464 3476 37516 3496
rect 37516 3476 37518 3496
rect 37462 3440 37518 3476
rect 36818 2080 36874 2136
rect 1398 720 1454 776
rect 38198 720 38254 776
rect 37186 40 37242 96
<< metal3 >>
rect 200 39538 800 39568
rect 3417 39538 3483 39541
rect 200 39536 3483 39538
rect 200 39480 3422 39536
rect 3478 39480 3483 39536
rect 200 39478 3483 39480
rect 200 39448 800 39478
rect 3417 39475 3483 39478
rect 200 38858 800 38888
rect 1577 38858 1643 38861
rect 200 38856 1643 38858
rect 200 38800 1582 38856
rect 1638 38800 1643 38856
rect 200 38798 1643 38800
rect 200 38768 800 38798
rect 1577 38795 1643 38798
rect 37457 38858 37523 38861
rect 39200 38858 39800 38888
rect 37457 38856 39800 38858
rect 37457 38800 37462 38856
rect 37518 38800 39800 38856
rect 37457 38798 39800 38800
rect 37457 38795 37523 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2865 37498 2931 37501
rect 200 37496 2931 37498
rect 200 37440 2870 37496
rect 2926 37440 2931 37496
rect 200 37438 2931 37440
rect 200 37408 800 37438
rect 2865 37435 2931 37438
rect 37181 37498 37247 37501
rect 39200 37498 39800 37528
rect 37181 37496 39800 37498
rect 37181 37440 37186 37496
rect 37242 37440 39800 37496
rect 37181 37438 39800 37440
rect 37181 37435 37247 37438
rect 39200 37408 39800 37438
rect 10501 37362 10567 37365
rect 18321 37362 18387 37365
rect 10501 37360 18387 37362
rect 10501 37304 10506 37360
rect 10562 37304 18326 37360
rect 18382 37304 18387 37360
rect 10501 37302 18387 37304
rect 10501 37299 10567 37302
rect 18321 37299 18387 37302
rect 19425 37362 19491 37365
rect 26325 37362 26391 37365
rect 19425 37360 26391 37362
rect 19425 37304 19430 37360
rect 19486 37304 26330 37360
rect 26386 37304 26391 37360
rect 19425 37302 26391 37304
rect 19425 37299 19491 37302
rect 26325 37299 26391 37302
rect 35157 37362 35223 37365
rect 35566 37362 35572 37364
rect 35157 37360 35572 37362
rect 35157 37304 35162 37360
rect 35218 37304 35572 37360
rect 35157 37302 35572 37304
rect 35157 37299 35223 37302
rect 35566 37300 35572 37302
rect 35636 37300 35642 37364
rect 11697 37226 11763 37229
rect 17033 37226 17099 37229
rect 25865 37226 25931 37229
rect 11697 37224 17099 37226
rect 11697 37168 11702 37224
rect 11758 37168 17038 37224
rect 17094 37168 17099 37224
rect 11697 37166 17099 37168
rect 11697 37163 11763 37166
rect 17033 37163 17099 37166
rect 17174 37224 25931 37226
rect 17174 37168 25870 37224
rect 25926 37168 25931 37224
rect 17174 37166 25931 37168
rect 17174 37090 17234 37166
rect 25865 37163 25931 37166
rect 2730 37030 17234 37090
rect 1669 36954 1735 36957
rect 2730 36954 2790 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 1669 36952 2790 36954
rect 1669 36896 1674 36952
rect 1730 36896 2790 36952
rect 1669 36894 2790 36896
rect 11789 36954 11855 36957
rect 15285 36954 15351 36957
rect 11789 36952 15351 36954
rect 11789 36896 11794 36952
rect 11850 36896 15290 36952
rect 15346 36896 15351 36952
rect 11789 36894 15351 36896
rect 1669 36891 1735 36894
rect 11789 36891 11855 36894
rect 15285 36891 15351 36894
rect 7005 36818 7071 36821
rect 37549 36818 37615 36821
rect 7005 36816 37615 36818
rect 7005 36760 7010 36816
rect 7066 36760 37554 36816
rect 37610 36760 37615 36816
rect 7005 36758 37615 36760
rect 7005 36755 7071 36758
rect 37549 36755 37615 36758
rect 8569 36682 8635 36685
rect 36169 36682 36235 36685
rect 8569 36680 36235 36682
rect 8569 36624 8574 36680
rect 8630 36624 36174 36680
rect 36230 36624 36235 36680
rect 8569 36622 36235 36624
rect 8569 36619 8635 36622
rect 36169 36619 36235 36622
rect 9029 36546 9095 36549
rect 9438 36546 9444 36548
rect 9029 36544 9444 36546
rect 9029 36488 9034 36544
rect 9090 36488 9444 36544
rect 9029 36486 9444 36488
rect 9029 36483 9095 36486
rect 9438 36484 9444 36486
rect 9508 36484 9514 36548
rect 10133 36546 10199 36549
rect 11881 36546 11947 36549
rect 10133 36544 11947 36546
rect 10133 36488 10138 36544
rect 10194 36488 11886 36544
rect 11942 36488 11947 36544
rect 10133 36486 11947 36488
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 9446 36410 9506 36484
rect 10133 36483 10199 36486
rect 11881 36483 11947 36486
rect 12065 36546 12131 36549
rect 16297 36546 16363 36549
rect 12065 36544 16363 36546
rect 12065 36488 12070 36544
rect 12126 36488 16302 36544
rect 16358 36488 16363 36544
rect 12065 36486 16363 36488
rect 12065 36483 12131 36486
rect 16297 36483 16363 36486
rect 17033 36546 17099 36549
rect 20897 36546 20963 36549
rect 21173 36546 21239 36549
rect 17033 36544 21239 36546
rect 17033 36488 17038 36544
rect 17094 36488 20902 36544
rect 20958 36488 21178 36544
rect 21234 36488 21239 36544
rect 17033 36486 21239 36488
rect 17033 36483 17099 36486
rect 20897 36483 20963 36486
rect 21173 36483 21239 36486
rect 22737 36546 22803 36549
rect 24853 36546 24919 36549
rect 22737 36544 24919 36546
rect 22737 36488 22742 36544
rect 22798 36488 24858 36544
rect 24914 36488 24919 36544
rect 22737 36486 24919 36488
rect 22737 36483 22803 36486
rect 24853 36483 24919 36486
rect 33133 36548 33199 36549
rect 33133 36544 33180 36548
rect 33244 36546 33250 36548
rect 33133 36488 33138 36544
rect 33133 36484 33180 36488
rect 33244 36486 33290 36546
rect 33244 36484 33250 36486
rect 33133 36483 33199 36484
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 29913 36410 29979 36413
rect 30741 36410 30807 36413
rect 9446 36408 30807 36410
rect 9446 36352 29918 36408
rect 29974 36352 30746 36408
rect 30802 36352 30807 36408
rect 9446 36350 30807 36352
rect 29913 36347 29979 36350
rect 30741 36347 30807 36350
rect 32305 36410 32371 36413
rect 32438 36410 32444 36412
rect 32305 36408 32444 36410
rect 32305 36352 32310 36408
rect 32366 36352 32444 36408
rect 32305 36350 32444 36352
rect 32305 36347 32371 36350
rect 32438 36348 32444 36350
rect 32508 36348 32514 36412
rect 6453 36274 6519 36277
rect 30005 36274 30071 36277
rect 6453 36272 30071 36274
rect 6453 36216 6458 36272
rect 6514 36216 30010 36272
rect 30066 36216 30071 36272
rect 6453 36214 30071 36216
rect 6453 36211 6519 36214
rect 30005 36211 30071 36214
rect 200 36138 800 36168
rect 1761 36138 1827 36141
rect 200 36136 1827 36138
rect 200 36080 1766 36136
rect 1822 36080 1827 36136
rect 200 36078 1827 36080
rect 200 36048 800 36078
rect 1761 36075 1827 36078
rect 11053 36138 11119 36141
rect 20621 36138 20687 36141
rect 11053 36136 20687 36138
rect 11053 36080 11058 36136
rect 11114 36080 20626 36136
rect 20682 36080 20687 36136
rect 11053 36078 20687 36080
rect 11053 36075 11119 36078
rect 20621 36075 20687 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 10317 36002 10383 36005
rect 11237 36002 11303 36005
rect 10317 36000 11303 36002
rect 10317 35944 10322 36000
rect 10378 35944 11242 36000
rect 11298 35944 11303 36000
rect 10317 35942 11303 35944
rect 10317 35939 10383 35942
rect 11237 35939 11303 35942
rect 28993 36002 29059 36005
rect 29126 36002 29132 36004
rect 28993 36000 29132 36002
rect 28993 35944 28998 36000
rect 29054 35944 29132 36000
rect 28993 35942 29132 35944
rect 28993 35939 29059 35942
rect 29126 35940 29132 35942
rect 29196 35940 29202 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 10593 35866 10659 35869
rect 12157 35866 12223 35869
rect 10593 35864 12223 35866
rect 10593 35808 10598 35864
rect 10654 35808 12162 35864
rect 12218 35808 12223 35864
rect 10593 35806 12223 35808
rect 10593 35803 10659 35806
rect 12157 35803 12223 35806
rect 1669 35730 1735 35733
rect 30465 35730 30531 35733
rect 1669 35728 30531 35730
rect 1669 35672 1674 35728
rect 1730 35672 30470 35728
rect 30526 35672 30531 35728
rect 1669 35670 30531 35672
rect 1669 35667 1735 35670
rect 30465 35667 30531 35670
rect 2405 35594 2471 35597
rect 27429 35594 27495 35597
rect 2405 35592 27495 35594
rect 2405 35536 2410 35592
rect 2466 35536 27434 35592
rect 27490 35536 27495 35592
rect 2405 35534 27495 35536
rect 2405 35531 2471 35534
rect 27429 35531 27495 35534
rect 200 35368 800 35488
rect 10133 35458 10199 35461
rect 23013 35458 23079 35461
rect 10133 35456 23079 35458
rect 10133 35400 10138 35456
rect 10194 35400 23018 35456
rect 23074 35400 23079 35456
rect 10133 35398 23079 35400
rect 10133 35395 10199 35398
rect 23013 35395 23079 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 10869 35322 10935 35325
rect 13169 35322 13235 35325
rect 10869 35320 13235 35322
rect 10869 35264 10874 35320
rect 10930 35264 13174 35320
rect 13230 35264 13235 35320
rect 10869 35262 13235 35264
rect 10869 35259 10935 35262
rect 13169 35259 13235 35262
rect 13629 35322 13695 35325
rect 17953 35322 18019 35325
rect 13629 35320 18019 35322
rect 13629 35264 13634 35320
rect 13690 35264 17958 35320
rect 18014 35264 18019 35320
rect 13629 35262 18019 35264
rect 13629 35259 13695 35262
rect 17953 35259 18019 35262
rect 10961 35186 11027 35189
rect 28441 35186 28507 35189
rect 10961 35184 28507 35186
rect 10961 35128 10966 35184
rect 11022 35128 28446 35184
rect 28502 35128 28507 35184
rect 10961 35126 28507 35128
rect 10961 35123 11027 35126
rect 28441 35123 28507 35126
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 10685 34642 10751 34645
rect 11881 34642 11947 34645
rect 10685 34640 11947 34642
rect 10685 34584 10690 34640
rect 10746 34584 11886 34640
rect 11942 34584 11947 34640
rect 10685 34582 11947 34584
rect 10685 34579 10751 34582
rect 11881 34579 11947 34582
rect 15561 34642 15627 34645
rect 15694 34642 15700 34644
rect 15561 34640 15700 34642
rect 15561 34584 15566 34640
rect 15622 34584 15700 34640
rect 15561 34582 15700 34584
rect 15561 34579 15627 34582
rect 15694 34580 15700 34582
rect 15764 34580 15770 34644
rect 9305 34506 9371 34509
rect 15101 34506 15167 34509
rect 9305 34504 15167 34506
rect 9305 34448 9310 34504
rect 9366 34448 15106 34504
rect 15162 34448 15167 34504
rect 9305 34446 15167 34448
rect 9305 34443 9371 34446
rect 15101 34443 15167 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 15561 34234 15627 34237
rect 16665 34234 16731 34237
rect 15561 34232 16731 34234
rect 15561 34176 15566 34232
rect 15622 34176 16670 34232
rect 16726 34176 16731 34232
rect 15561 34174 16731 34176
rect 15561 34171 15627 34174
rect 16665 34171 16731 34174
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 12893 34098 12959 34101
rect 17033 34098 17099 34101
rect 12893 34096 17099 34098
rect 12893 34040 12898 34096
rect 12954 34040 17038 34096
rect 17094 34040 17099 34096
rect 12893 34038 17099 34040
rect 12893 34035 12959 34038
rect 17033 34035 17099 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 14365 33962 14431 33965
rect 20713 33962 20779 33965
rect 14365 33960 20779 33962
rect 14365 33904 14370 33960
rect 14426 33904 20718 33960
rect 20774 33904 20779 33960
rect 14365 33902 20779 33904
rect 14365 33899 14431 33902
rect 20713 33899 20779 33902
rect 11973 33826 12039 33829
rect 19333 33826 19399 33829
rect 11973 33824 19399 33826
rect 11973 33768 11978 33824
rect 12034 33768 19338 33824
rect 19394 33768 19399 33824
rect 11973 33766 19399 33768
rect 11973 33763 12039 33766
rect 19333 33763 19399 33766
rect 31845 33826 31911 33829
rect 33910 33826 33916 33828
rect 31845 33824 33916 33826
rect 31845 33768 31850 33824
rect 31906 33768 33916 33824
rect 31845 33766 33916 33768
rect 31845 33763 31911 33766
rect 33910 33764 33916 33766
rect 33980 33764 33986 33828
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 13169 33690 13235 33693
rect 15561 33690 15627 33693
rect 17585 33690 17651 33693
rect 13169 33688 17651 33690
rect 13169 33632 13174 33688
rect 13230 33632 15566 33688
rect 15622 33632 17590 33688
rect 17646 33632 17651 33688
rect 13169 33630 17651 33632
rect 13169 33627 13235 33630
rect 15561 33627 15627 33630
rect 17585 33627 17651 33630
rect 15101 33554 15167 33557
rect 25589 33554 25655 33557
rect 15101 33552 25655 33554
rect 15101 33496 15106 33552
rect 15162 33496 25594 33552
rect 25650 33496 25655 33552
rect 15101 33494 25655 33496
rect 15101 33491 15167 33494
rect 25589 33491 25655 33494
rect 10777 33418 10843 33421
rect 19885 33418 19951 33421
rect 10777 33416 19951 33418
rect 10777 33360 10782 33416
rect 10838 33360 19890 33416
rect 19946 33360 19951 33416
rect 10777 33358 19951 33360
rect 10777 33355 10843 33358
rect 19885 33355 19951 33358
rect 34646 33356 34652 33420
rect 34716 33418 34722 33420
rect 35525 33418 35591 33421
rect 34716 33416 35591 33418
rect 34716 33360 35530 33416
rect 35586 33360 35591 33416
rect 34716 33358 35591 33360
rect 34716 33356 34722 33358
rect 35525 33355 35591 33358
rect 11053 33282 11119 33285
rect 18597 33282 18663 33285
rect 11053 33280 18663 33282
rect 11053 33224 11058 33280
rect 11114 33224 18602 33280
rect 18658 33224 18663 33280
rect 11053 33222 18663 33224
rect 11053 33219 11119 33222
rect 18597 33219 18663 33222
rect 27613 33284 27679 33285
rect 27613 33280 27660 33284
rect 27724 33282 27730 33284
rect 27613 33224 27618 33280
rect 27613 33220 27660 33224
rect 27724 33222 27770 33282
rect 27724 33220 27730 33222
rect 27613 33219 27679 33220
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 11697 33146 11763 33149
rect 18781 33146 18847 33149
rect 11697 33144 18847 33146
rect 11697 33088 11702 33144
rect 11758 33088 18786 33144
rect 18842 33088 18847 33144
rect 11697 33086 18847 33088
rect 11697 33083 11763 33086
rect 18781 33083 18847 33086
rect 10133 33010 10199 33013
rect 18873 33010 18939 33013
rect 10133 33008 18939 33010
rect 10133 32952 10138 33008
rect 10194 32952 18878 33008
rect 18934 32952 18939 33008
rect 10133 32950 18939 32952
rect 10133 32947 10199 32950
rect 18873 32947 18939 32950
rect 14457 32874 14523 32877
rect 24577 32874 24643 32877
rect 14457 32872 24643 32874
rect 14457 32816 14462 32872
rect 14518 32816 24582 32872
rect 24638 32816 24643 32872
rect 14457 32814 24643 32816
rect 14457 32811 14523 32814
rect 24577 32811 24643 32814
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 38101 32738 38167 32741
rect 39200 32738 39800 32768
rect 38101 32736 39800 32738
rect 38101 32680 38106 32736
rect 38162 32680 39800 32736
rect 38101 32678 39800 32680
rect 38101 32675 38167 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 8293 32466 8359 32469
rect 20345 32466 20411 32469
rect 8293 32464 20411 32466
rect 8293 32408 8298 32464
rect 8354 32408 20350 32464
rect 20406 32408 20411 32464
rect 8293 32406 20411 32408
rect 8293 32403 8359 32406
rect 20345 32403 20411 32406
rect 13537 32330 13603 32333
rect 19977 32330 20043 32333
rect 25497 32332 25563 32333
rect 25446 32330 25452 32332
rect 13537 32328 20043 32330
rect 13537 32272 13542 32328
rect 13598 32272 19982 32328
rect 20038 32272 20043 32328
rect 13537 32270 20043 32272
rect 25406 32270 25452 32330
rect 25516 32328 25563 32332
rect 25558 32272 25563 32328
rect 13537 32267 13603 32270
rect 19977 32267 20043 32270
rect 25446 32268 25452 32270
rect 25516 32268 25563 32272
rect 25497 32267 25563 32268
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 25630 31996 25636 32060
rect 25700 32058 25706 32060
rect 25773 32058 25839 32061
rect 25700 32056 25839 32058
rect 25700 32000 25778 32056
rect 25834 32000 25839 32056
rect 25700 31998 25839 32000
rect 25700 31996 25706 31998
rect 25773 31995 25839 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 19057 31922 19123 31925
rect 20989 31922 21055 31925
rect 19057 31920 21055 31922
rect 19057 31864 19062 31920
rect 19118 31864 20994 31920
rect 21050 31864 21055 31920
rect 19057 31862 21055 31864
rect 19057 31859 19123 31862
rect 20989 31859 21055 31862
rect 15745 31786 15811 31789
rect 20161 31786 20227 31789
rect 15745 31784 20227 31786
rect 15745 31728 15750 31784
rect 15806 31728 20166 31784
rect 20222 31728 20227 31784
rect 15745 31726 20227 31728
rect 15745 31723 15811 31726
rect 20161 31723 20227 31726
rect 36261 31788 36327 31789
rect 36261 31784 36308 31788
rect 36372 31786 36378 31788
rect 36261 31728 36266 31784
rect 36261 31724 36308 31728
rect 36372 31726 36418 31786
rect 36372 31724 36378 31726
rect 36261 31723 36327 31724
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 8201 31378 8267 31381
rect 12801 31378 12867 31381
rect 18505 31378 18571 31381
rect 8201 31376 18571 31378
rect 8201 31320 8206 31376
rect 8262 31320 12806 31376
rect 12862 31320 18510 31376
rect 18566 31320 18571 31376
rect 8201 31318 18571 31320
rect 8201 31315 8267 31318
rect 12801 31315 12867 31318
rect 18505 31315 18571 31318
rect 11053 31242 11119 31245
rect 27797 31242 27863 31245
rect 11053 31240 27863 31242
rect 11053 31184 11058 31240
rect 11114 31184 27802 31240
rect 27858 31184 27863 31240
rect 11053 31182 27863 31184
rect 11053 31179 11119 31182
rect 27797 31179 27863 31182
rect 13537 31106 13603 31109
rect 17033 31106 17099 31109
rect 13537 31104 17099 31106
rect 13537 31048 13542 31104
rect 13598 31048 17038 31104
rect 17094 31048 17099 31104
rect 13537 31046 17099 31048
rect 13537 31043 13603 31046
rect 17033 31043 17099 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 34605 30972 34671 30973
rect 34605 30970 34652 30972
rect 34560 30968 34652 30970
rect 34560 30912 34610 30968
rect 34560 30910 34652 30912
rect 34605 30908 34652 30910
rect 34716 30908 34722 30972
rect 34605 30907 34671 30908
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 38193 30698 38259 30701
rect 39200 30698 39800 30728
rect 38193 30696 39800 30698
rect 38193 30640 38198 30696
rect 38254 30640 39800 30696
rect 38193 30638 39800 30640
rect 38193 30635 38259 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 14365 30426 14431 30429
rect 19374 30426 19380 30428
rect 14365 30424 19380 30426
rect 14365 30368 14370 30424
rect 14426 30368 19380 30424
rect 14365 30366 19380 30368
rect 14365 30363 14431 30366
rect 19374 30364 19380 30366
rect 19444 30364 19450 30428
rect 24577 30426 24643 30429
rect 24710 30426 24716 30428
rect 24577 30424 24716 30426
rect 24577 30368 24582 30424
rect 24638 30368 24716 30424
rect 24577 30366 24716 30368
rect 24577 30363 24643 30366
rect 24710 30364 24716 30366
rect 24780 30364 24786 30428
rect 28625 30426 28691 30429
rect 28758 30426 28764 30428
rect 28625 30424 28764 30426
rect 28625 30368 28630 30424
rect 28686 30368 28764 30424
rect 28625 30366 28764 30368
rect 28625 30363 28691 30366
rect 28758 30364 28764 30366
rect 28828 30364 28834 30428
rect 30230 30364 30236 30428
rect 30300 30426 30306 30428
rect 30557 30426 30623 30429
rect 30300 30424 30623 30426
rect 30300 30368 30562 30424
rect 30618 30368 30623 30424
rect 30300 30366 30623 30368
rect 30300 30364 30306 30366
rect 30557 30363 30623 30366
rect 31886 30364 31892 30428
rect 31956 30426 31962 30428
rect 32029 30426 32095 30429
rect 31956 30424 32095 30426
rect 31956 30368 32034 30424
rect 32090 30368 32095 30424
rect 31956 30366 32095 30368
rect 31956 30364 31962 30366
rect 32029 30363 32095 30366
rect 13169 30290 13235 30293
rect 19793 30290 19859 30293
rect 13169 30288 19859 30290
rect 13169 30232 13174 30288
rect 13230 30232 19798 30288
rect 19854 30232 19859 30288
rect 13169 30230 19859 30232
rect 13169 30227 13235 30230
rect 19793 30227 19859 30230
rect 21398 30228 21404 30292
rect 21468 30290 21474 30292
rect 25037 30290 25103 30293
rect 21468 30288 25103 30290
rect 21468 30232 25042 30288
rect 25098 30232 25103 30288
rect 21468 30230 25103 30232
rect 21468 30228 21474 30230
rect 25037 30227 25103 30230
rect 18873 30154 18939 30157
rect 20161 30154 20227 30157
rect 18873 30152 20227 30154
rect 18873 30096 18878 30152
rect 18934 30096 20166 30152
rect 20222 30096 20227 30152
rect 18873 30094 20227 30096
rect 18873 30091 18939 30094
rect 20161 30091 20227 30094
rect 31518 29956 31524 30020
rect 31588 30018 31594 30020
rect 31661 30018 31727 30021
rect 31588 30016 31727 30018
rect 31588 29960 31666 30016
rect 31722 29960 31727 30016
rect 31588 29958 31727 29960
rect 31588 29956 31594 29958
rect 31661 29955 31727 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 9438 29820 9444 29884
rect 9508 29882 9514 29884
rect 10869 29882 10935 29885
rect 9508 29880 10935 29882
rect 9508 29824 10874 29880
rect 10930 29824 10935 29880
rect 9508 29822 10935 29824
rect 9508 29820 9514 29822
rect 10869 29819 10935 29822
rect 19057 29882 19123 29885
rect 19793 29882 19859 29885
rect 19057 29880 19859 29882
rect 19057 29824 19062 29880
rect 19118 29824 19798 29880
rect 19854 29824 19859 29880
rect 19057 29822 19859 29824
rect 19057 29819 19123 29822
rect 19793 29819 19859 29822
rect 20161 29746 20227 29749
rect 17910 29744 20227 29746
rect 17910 29688 20166 29744
rect 20222 29688 20227 29744
rect 17910 29686 20227 29688
rect 13629 29610 13695 29613
rect 17910 29610 17970 29686
rect 20161 29683 20227 29686
rect 13629 29608 17970 29610
rect 13629 29552 13634 29608
rect 13690 29552 17970 29608
rect 13629 29550 17970 29552
rect 19333 29610 19399 29613
rect 20713 29610 20779 29613
rect 19333 29608 20779 29610
rect 19333 29552 19338 29608
rect 19394 29552 20718 29608
rect 20774 29552 20779 29608
rect 19333 29550 20779 29552
rect 13629 29547 13695 29550
rect 19333 29547 19399 29550
rect 20713 29547 20779 29550
rect 19425 29476 19491 29477
rect 19374 29474 19380 29476
rect 19334 29414 19380 29474
rect 19444 29472 19491 29476
rect 19486 29416 19491 29472
rect 19374 29412 19380 29414
rect 19444 29412 19491 29416
rect 19425 29411 19491 29412
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 12801 29338 12867 29341
rect 18965 29338 19031 29341
rect 19241 29338 19307 29341
rect 12801 29336 19307 29338
rect 12801 29280 12806 29336
rect 12862 29280 18970 29336
rect 19026 29280 19246 29336
rect 19302 29280 19307 29336
rect 12801 29278 19307 29280
rect 12801 29275 12867 29278
rect 18965 29275 19031 29278
rect 19241 29275 19307 29278
rect 38193 29338 38259 29341
rect 39200 29338 39800 29368
rect 38193 29336 39800 29338
rect 38193 29280 38198 29336
rect 38254 29280 39800 29336
rect 38193 29278 39800 29280
rect 38193 29275 38259 29278
rect 39200 29248 39800 29278
rect 19333 29202 19399 29205
rect 20345 29202 20411 29205
rect 19333 29200 20411 29202
rect 19333 29144 19338 29200
rect 19394 29144 20350 29200
rect 20406 29144 20411 29200
rect 19333 29142 20411 29144
rect 19333 29139 19399 29142
rect 20345 29139 20411 29142
rect 25998 29140 26004 29204
rect 26068 29202 26074 29204
rect 33225 29202 33291 29205
rect 26068 29200 33291 29202
rect 26068 29144 33230 29200
rect 33286 29144 33291 29200
rect 26068 29142 33291 29144
rect 26068 29140 26074 29142
rect 33225 29139 33291 29142
rect 10961 29066 11027 29069
rect 15101 29066 15167 29069
rect 18413 29066 18479 29069
rect 10961 29064 18479 29066
rect 10961 29008 10966 29064
rect 11022 29008 15106 29064
rect 15162 29008 18418 29064
rect 18474 29008 18479 29064
rect 10961 29006 18479 29008
rect 10961 29003 11027 29006
rect 15101 29003 15167 29006
rect 18413 29003 18479 29006
rect 31293 29068 31359 29069
rect 32213 29068 32279 29069
rect 31293 29064 31340 29068
rect 31404 29066 31410 29068
rect 31293 29008 31298 29064
rect 31293 29004 31340 29008
rect 31404 29006 31450 29066
rect 32213 29064 32260 29068
rect 32324 29066 32330 29068
rect 32213 29008 32218 29064
rect 31404 29004 31410 29006
rect 32213 29004 32260 29008
rect 32324 29006 32370 29066
rect 32324 29004 32330 29006
rect 32990 29004 32996 29068
rect 33060 29066 33066 29068
rect 36077 29066 36143 29069
rect 33060 29064 36143 29066
rect 33060 29008 36082 29064
rect 36138 29008 36143 29064
rect 33060 29006 36143 29008
rect 33060 29004 33066 29006
rect 31293 29003 31359 29004
rect 32213 29003 32279 29004
rect 36077 29003 36143 29006
rect 17677 28930 17743 28933
rect 17861 28930 17927 28933
rect 17677 28928 17927 28930
rect 17677 28872 17682 28928
rect 17738 28872 17866 28928
rect 17922 28872 17927 28928
rect 17677 28870 17927 28872
rect 17677 28867 17743 28870
rect 17861 28867 17927 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 10501 28794 10567 28797
rect 17953 28794 18019 28797
rect 10501 28792 18019 28794
rect 10501 28736 10506 28792
rect 10562 28736 17958 28792
rect 18014 28736 18019 28792
rect 10501 28734 18019 28736
rect 10501 28731 10567 28734
rect 17953 28731 18019 28734
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 14917 28522 14983 28525
rect 17677 28522 17743 28525
rect 14917 28520 17743 28522
rect 14917 28464 14922 28520
rect 14978 28464 17682 28520
rect 17738 28464 17743 28520
rect 14917 28462 17743 28464
rect 14917 28459 14983 28462
rect 17677 28459 17743 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 13077 27842 13143 27845
rect 15837 27842 15903 27845
rect 13077 27840 15903 27842
rect 13077 27784 13082 27840
rect 13138 27784 15842 27840
rect 15898 27784 15903 27840
rect 13077 27782 15903 27784
rect 13077 27779 13143 27782
rect 15837 27779 15903 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 34421 26348 34487 26349
rect 34421 26344 34468 26348
rect 34532 26346 34538 26348
rect 34421 26288 34426 26344
rect 34421 26284 34468 26288
rect 34532 26286 34578 26346
rect 34532 26284 34538 26286
rect 34421 26283 34487 26284
rect 23422 26148 23428 26212
rect 23492 26210 23498 26212
rect 28257 26210 28323 26213
rect 23492 26208 28323 26210
rect 23492 26152 28262 26208
rect 28318 26152 28323 26208
rect 23492 26150 28323 26152
rect 23492 26148 23498 26150
rect 28257 26147 28323 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1761 25938 1827 25941
rect 200 25936 1827 25938
rect 200 25880 1766 25936
rect 1822 25880 1827 25936
rect 200 25878 1827 25880
rect 200 25848 800 25878
rect 1761 25875 1827 25878
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 24894 25740 24900 25804
rect 24964 25802 24970 25804
rect 37641 25802 37707 25805
rect 24964 25800 37707 25802
rect 24964 25744 37646 25800
rect 37702 25744 37707 25800
rect 24964 25742 37707 25744
rect 24964 25740 24970 25742
rect 37641 25739 37707 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 13629 25394 13695 25397
rect 20989 25394 21055 25397
rect 13629 25392 21055 25394
rect 13629 25336 13634 25392
rect 13690 25336 20994 25392
rect 21050 25336 21055 25392
rect 13629 25334 21055 25336
rect 13629 25331 13695 25334
rect 20989 25331 21055 25334
rect 19374 25196 19380 25260
rect 19444 25258 19450 25260
rect 19701 25258 19767 25261
rect 28901 25258 28967 25261
rect 19444 25256 28967 25258
rect 19444 25200 19706 25256
rect 19762 25200 28906 25256
rect 28962 25200 28967 25256
rect 19444 25198 28967 25200
rect 19444 25196 19450 25198
rect 19701 25195 19767 25198
rect 28901 25195 28967 25198
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 30414 24924 30420 24988
rect 30484 24986 30490 24988
rect 30741 24986 30807 24989
rect 30484 24984 30807 24986
rect 30484 24928 30746 24984
rect 30802 24928 30807 24984
rect 30484 24926 30807 24928
rect 30484 24924 30490 24926
rect 30741 24923 30807 24926
rect 33685 24988 33751 24989
rect 33685 24984 33732 24988
rect 33796 24986 33802 24988
rect 33685 24928 33690 24984
rect 33685 24924 33732 24928
rect 33796 24926 33842 24986
rect 33796 24924 33802 24926
rect 33685 24923 33751 24924
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19609 24306 19675 24309
rect 24853 24306 24919 24309
rect 19609 24304 24919 24306
rect 19609 24248 19614 24304
rect 19670 24248 24858 24304
rect 24914 24248 24919 24304
rect 19609 24246 24919 24248
rect 19609 24243 19675 24246
rect 24853 24243 24919 24246
rect 18597 24170 18663 24173
rect 19517 24170 19583 24173
rect 18597 24168 19583 24170
rect 18597 24112 18602 24168
rect 18658 24112 19522 24168
rect 19578 24112 19583 24168
rect 18597 24110 19583 24112
rect 18597 24107 18663 24110
rect 19517 24107 19583 24110
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 37457 23898 37523 23901
rect 39200 23898 39800 23928
rect 37457 23896 39800 23898
rect 37457 23840 37462 23896
rect 37518 23840 39800 23896
rect 37457 23838 39800 23840
rect 37457 23835 37523 23838
rect 39200 23808 39800 23838
rect 27613 23490 27679 23493
rect 27838 23490 27844 23492
rect 27613 23488 27844 23490
rect 27613 23432 27618 23488
rect 27674 23432 27844 23488
rect 27613 23430 27844 23432
rect 27613 23427 27679 23430
rect 27838 23428 27844 23430
rect 27908 23428 27914 23492
rect 35750 23428 35756 23492
rect 35820 23490 35826 23492
rect 36445 23490 36511 23493
rect 35820 23488 36511 23490
rect 35820 23432 36450 23488
rect 36506 23432 36511 23488
rect 35820 23430 36511 23432
rect 35820 23428 35826 23430
rect 36445 23427 36511 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 30046 23020 30052 23084
rect 30116 23082 30122 23084
rect 31201 23082 31267 23085
rect 32673 23082 32739 23085
rect 30116 23080 32739 23082
rect 30116 23024 31206 23080
rect 31262 23024 32678 23080
rect 32734 23024 32739 23080
rect 30116 23022 32739 23024
rect 30116 23020 30122 23022
rect 31201 23019 31267 23022
rect 32673 23019 32739 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 20069 22810 20135 22813
rect 20253 22810 20319 22813
rect 20069 22808 20319 22810
rect 20069 22752 20074 22808
rect 20130 22752 20258 22808
rect 20314 22752 20319 22808
rect 20069 22750 20319 22752
rect 20069 22747 20135 22750
rect 20253 22747 20319 22750
rect 31845 22810 31911 22813
rect 35709 22810 35775 22813
rect 36445 22810 36511 22813
rect 31845 22808 36511 22810
rect 31845 22752 31850 22808
rect 31906 22752 35714 22808
rect 35770 22752 36450 22808
rect 36506 22752 36511 22808
rect 31845 22750 36511 22752
rect 31845 22747 31911 22750
rect 35709 22747 35775 22750
rect 36445 22747 36511 22750
rect 15694 22612 15700 22676
rect 15764 22674 15770 22676
rect 23606 22674 23612 22676
rect 15764 22614 23612 22674
rect 15764 22612 15770 22614
rect 23606 22612 23612 22614
rect 23676 22612 23682 22676
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 19333 22404 19399 22405
rect 19333 22400 19380 22404
rect 19444 22402 19450 22404
rect 19333 22344 19338 22400
rect 19333 22340 19380 22344
rect 19444 22342 19490 22402
rect 19444 22340 19450 22342
rect 19333 22339 19399 22340
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 16849 21994 16915 21997
rect 20897 21994 20963 21997
rect 23422 21994 23428 21996
rect 16849 21992 20730 21994
rect 16849 21936 16854 21992
rect 16910 21936 20730 21992
rect 16849 21934 20730 21936
rect 16849 21931 16915 21934
rect 20670 21858 20730 21934
rect 20897 21992 23428 21994
rect 20897 21936 20902 21992
rect 20958 21936 23428 21992
rect 20897 21934 23428 21936
rect 20897 21931 20963 21934
rect 23422 21932 23428 21934
rect 23492 21932 23498 21996
rect 25221 21994 25287 21997
rect 26325 21994 26391 21997
rect 25221 21992 26391 21994
rect 25221 21936 25226 21992
rect 25282 21936 26330 21992
rect 26386 21936 26391 21992
rect 25221 21934 26391 21936
rect 25221 21931 25287 21934
rect 26325 21931 26391 21934
rect 37825 21994 37891 21997
rect 38142 21994 38148 21996
rect 37825 21992 38148 21994
rect 37825 21936 37830 21992
rect 37886 21936 38148 21992
rect 37825 21934 38148 21936
rect 37825 21931 37891 21934
rect 38142 21932 38148 21934
rect 38212 21932 38218 21996
rect 22737 21858 22803 21861
rect 20670 21856 22803 21858
rect 20670 21800 22742 21856
rect 22798 21800 22803 21856
rect 20670 21798 22803 21800
rect 22737 21795 22803 21798
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 11513 21586 11579 21589
rect 27613 21586 27679 21589
rect 11513 21584 27679 21586
rect 11513 21528 11518 21584
rect 11574 21528 27618 21584
rect 27674 21528 27679 21584
rect 11513 21526 27679 21528
rect 11513 21523 11579 21526
rect 27613 21523 27679 21526
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1761 21178 1827 21181
rect 200 21176 1827 21178
rect 200 21120 1766 21176
rect 1822 21120 1827 21176
rect 200 21118 1827 21120
rect 200 21088 800 21118
rect 1761 21115 1827 21118
rect 25037 21042 25103 21045
rect 28441 21042 28507 21045
rect 25037 21040 28507 21042
rect 25037 20984 25042 21040
rect 25098 20984 28446 21040
rect 28502 20984 28507 21040
rect 25037 20982 28507 20984
rect 25037 20979 25103 20982
rect 28441 20979 28507 20982
rect 32949 21042 33015 21045
rect 37273 21042 37339 21045
rect 32949 21040 37339 21042
rect 32949 20984 32954 21040
rect 33010 20984 37278 21040
rect 37334 20984 37339 21040
rect 32949 20982 37339 20984
rect 32949 20979 33015 20982
rect 37273 20979 37339 20982
rect 22645 20906 22711 20909
rect 25773 20906 25839 20909
rect 26693 20906 26759 20909
rect 27061 20906 27127 20909
rect 22645 20904 27127 20906
rect 22645 20848 22650 20904
rect 22706 20848 25778 20904
rect 25834 20848 26698 20904
rect 26754 20848 27066 20904
rect 27122 20848 27127 20904
rect 22645 20846 27127 20848
rect 22645 20843 22711 20846
rect 25773 20843 25839 20846
rect 26693 20843 26759 20846
rect 27061 20843 27127 20846
rect 27705 20770 27771 20773
rect 26742 20768 27771 20770
rect 26742 20712 27710 20768
rect 27766 20712 27771 20768
rect 26742 20710 27771 20712
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 21265 20634 21331 20637
rect 21398 20634 21404 20636
rect 21265 20632 21404 20634
rect 21265 20576 21270 20632
rect 21326 20576 21404 20632
rect 21265 20574 21404 20576
rect 21265 20571 21331 20574
rect 21398 20572 21404 20574
rect 21468 20572 21474 20636
rect 26601 20634 26667 20637
rect 26742 20634 26802 20710
rect 27705 20707 27771 20710
rect 26601 20632 26802 20634
rect 26601 20576 26606 20632
rect 26662 20576 26802 20632
rect 26601 20574 26802 20576
rect 26601 20571 26667 20574
rect 31150 20572 31156 20636
rect 31220 20634 31226 20636
rect 32581 20634 32647 20637
rect 31220 20632 32647 20634
rect 31220 20576 32586 20632
rect 32642 20576 32647 20632
rect 31220 20574 32647 20576
rect 31220 20572 31226 20574
rect 32581 20571 32647 20574
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 14917 20498 14983 20501
rect 30741 20500 30807 20501
rect 30741 20498 30788 20500
rect 14917 20496 30788 20498
rect 30852 20498 30858 20500
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 14917 20440 14922 20496
rect 14978 20440 30746 20496
rect 14917 20438 30788 20440
rect 14917 20435 14983 20438
rect 30741 20436 30788 20438
rect 30852 20438 30934 20498
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 30852 20436 30858 20438
rect 30741 20435 30807 20436
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 38193 20364 38259 20365
rect 38142 20300 38148 20364
rect 38212 20362 38259 20364
rect 38212 20360 38304 20362
rect 38254 20304 38304 20360
rect 38212 20302 38304 20304
rect 38212 20300 38259 20302
rect 38193 20299 38259 20300
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 21725 20090 21791 20093
rect 27153 20090 27219 20093
rect 21725 20088 27219 20090
rect 21725 20032 21730 20088
rect 21786 20032 27158 20088
rect 27214 20032 27219 20088
rect 21725 20030 27219 20032
rect 21725 20027 21791 20030
rect 27153 20027 27219 20030
rect 20621 19954 20687 19957
rect 30414 19954 30420 19956
rect 20621 19952 30420 19954
rect 20621 19896 20626 19952
rect 20682 19896 30420 19952
rect 20621 19894 30420 19896
rect 20621 19891 20687 19894
rect 30414 19892 30420 19894
rect 30484 19892 30490 19956
rect 33869 19954 33935 19957
rect 34646 19954 34652 19956
rect 33869 19952 34652 19954
rect 33869 19896 33874 19952
rect 33930 19896 34652 19952
rect 33869 19894 34652 19896
rect 33869 19891 33935 19894
rect 34646 19892 34652 19894
rect 34716 19892 34722 19956
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 26693 19546 26759 19549
rect 27981 19546 28047 19549
rect 26693 19544 28047 19546
rect 26693 19488 26698 19544
rect 26754 19488 27986 19544
rect 28042 19488 28047 19544
rect 26693 19486 28047 19488
rect 26693 19483 26759 19486
rect 27981 19483 28047 19486
rect 32305 19546 32371 19549
rect 34789 19546 34855 19549
rect 35433 19546 35499 19549
rect 32305 19544 35499 19546
rect 32305 19488 32310 19544
rect 32366 19488 34794 19544
rect 34850 19488 35438 19544
rect 35494 19488 35499 19544
rect 32305 19486 35499 19488
rect 32305 19483 32371 19486
rect 34789 19483 34855 19486
rect 35433 19483 35499 19486
rect 23606 19348 23612 19412
rect 23676 19410 23682 19412
rect 34973 19410 35039 19413
rect 23676 19408 36554 19410
rect 23676 19352 34978 19408
rect 35034 19352 36554 19408
rect 23676 19350 36554 19352
rect 23676 19348 23682 19350
rect 34973 19347 35039 19350
rect 33685 19274 33751 19277
rect 36302 19274 36308 19276
rect 33685 19272 36308 19274
rect 33685 19216 33690 19272
rect 33746 19216 36308 19272
rect 33685 19214 36308 19216
rect 33685 19211 33751 19214
rect 36302 19212 36308 19214
rect 36372 19212 36378 19276
rect 200 19138 800 19168
rect 1577 19138 1643 19141
rect 200 19136 1643 19138
rect 200 19080 1582 19136
rect 1638 19080 1643 19136
rect 200 19078 1643 19080
rect 200 19048 800 19078
rect 1577 19075 1643 19078
rect 29545 19138 29611 19141
rect 30046 19138 30052 19140
rect 29545 19136 30052 19138
rect 29545 19080 29550 19136
rect 29606 19080 30052 19136
rect 29545 19078 30052 19080
rect 29545 19075 29611 19078
rect 30046 19076 30052 19078
rect 30116 19076 30122 19140
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 31201 19002 31267 19005
rect 32397 19002 32463 19005
rect 31201 19000 32463 19002
rect 31201 18944 31206 19000
rect 31262 18944 32402 19000
rect 32458 18944 32463 19000
rect 31201 18942 32463 18944
rect 36494 19002 36554 19350
rect 37457 19138 37523 19141
rect 39200 19138 39800 19168
rect 37457 19136 39800 19138
rect 37457 19080 37462 19136
rect 37518 19080 39800 19136
rect 37457 19078 39800 19080
rect 37457 19075 37523 19078
rect 39200 19048 39800 19078
rect 37457 19002 37523 19005
rect 36494 19000 37523 19002
rect 36494 18944 37462 19000
rect 37518 18944 37523 19000
rect 36494 18942 37523 18944
rect 31201 18939 31267 18942
rect 32397 18939 32463 18942
rect 37457 18939 37523 18942
rect 24761 18866 24827 18869
rect 26049 18866 26115 18869
rect 27838 18866 27844 18868
rect 24761 18864 27844 18866
rect 24761 18808 24766 18864
rect 24822 18808 26054 18864
rect 26110 18808 27844 18864
rect 24761 18806 27844 18808
rect 24761 18803 24827 18806
rect 26049 18803 26115 18806
rect 27838 18804 27844 18806
rect 27908 18804 27914 18868
rect 31569 18866 31635 18869
rect 35985 18866 36051 18869
rect 31569 18864 36051 18866
rect 31569 18808 31574 18864
rect 31630 18808 35990 18864
rect 36046 18808 36051 18864
rect 31569 18806 36051 18808
rect 31569 18803 31635 18806
rect 35985 18803 36051 18806
rect 30925 18730 30991 18733
rect 32581 18730 32647 18733
rect 30925 18728 32647 18730
rect 30925 18672 30930 18728
rect 30986 18672 32586 18728
rect 32642 18672 32647 18728
rect 30925 18670 32647 18672
rect 30925 18667 30991 18670
rect 32581 18667 32647 18670
rect 30373 18594 30439 18597
rect 33225 18594 33291 18597
rect 30373 18592 33291 18594
rect 30373 18536 30378 18592
rect 30434 18536 33230 18592
rect 33286 18536 33291 18592
rect 30373 18534 33291 18536
rect 30373 18531 30439 18534
rect 33225 18531 33291 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 39200 18368 39800 18488
rect 23565 18322 23631 18325
rect 27521 18322 27587 18325
rect 23565 18320 27587 18322
rect 23565 18264 23570 18320
rect 23626 18264 27526 18320
rect 27582 18264 27587 18320
rect 23565 18262 27587 18264
rect 23565 18259 23631 18262
rect 27521 18259 27587 18262
rect 18965 18186 19031 18189
rect 25630 18186 25636 18188
rect 18965 18184 25636 18186
rect 18965 18128 18970 18184
rect 19026 18128 25636 18184
rect 18965 18126 25636 18128
rect 18965 18123 19031 18126
rect 25630 18124 25636 18126
rect 25700 18186 25706 18188
rect 32949 18186 33015 18189
rect 25700 18184 33015 18186
rect 25700 18128 32954 18184
rect 33010 18128 33015 18184
rect 25700 18126 33015 18128
rect 25700 18124 25706 18126
rect 32949 18123 33015 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 28758 17852 28764 17916
rect 28828 17914 28834 17916
rect 30373 17914 30439 17917
rect 28828 17912 30439 17914
rect 28828 17856 30378 17912
rect 30434 17856 30439 17912
rect 28828 17854 30439 17856
rect 28828 17852 28834 17854
rect 30373 17851 30439 17854
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 23289 17778 23355 17781
rect 28533 17778 28599 17781
rect 23289 17776 28599 17778
rect 23289 17720 23294 17776
rect 23350 17720 28538 17776
rect 28594 17720 28599 17776
rect 23289 17718 28599 17720
rect 23289 17715 23355 17718
rect 28533 17715 28599 17718
rect 29177 17778 29243 17781
rect 33041 17778 33107 17781
rect 29177 17776 33107 17778
rect 29177 17720 29182 17776
rect 29238 17720 33046 17776
rect 33102 17720 33107 17776
rect 29177 17718 33107 17720
rect 29177 17715 29243 17718
rect 33041 17715 33107 17718
rect 29453 17642 29519 17645
rect 31017 17642 31083 17645
rect 36169 17644 36235 17645
rect 29453 17640 31083 17642
rect 29453 17584 29458 17640
rect 29514 17584 31022 17640
rect 31078 17584 31083 17640
rect 29453 17582 31083 17584
rect 29453 17579 29519 17582
rect 31017 17579 31083 17582
rect 35566 17580 35572 17644
rect 35636 17642 35642 17644
rect 36118 17642 36124 17644
rect 35636 17582 36124 17642
rect 36188 17642 36235 17644
rect 36188 17640 36280 17642
rect 36230 17584 36280 17640
rect 35636 17580 35642 17582
rect 36118 17580 36124 17582
rect 36188 17582 36280 17584
rect 36188 17580 36235 17582
rect 36169 17579 36235 17580
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 25446 17308 25452 17372
rect 25516 17370 25522 17372
rect 27245 17370 27311 17373
rect 25516 17368 27311 17370
rect 25516 17312 27250 17368
rect 27306 17312 27311 17368
rect 25516 17310 27311 17312
rect 25516 17308 25522 17310
rect 27245 17307 27311 17310
rect 35934 17172 35940 17236
rect 36004 17234 36010 17236
rect 38285 17234 38351 17237
rect 36004 17232 38351 17234
rect 36004 17176 38290 17232
rect 38346 17176 38351 17232
rect 36004 17174 38351 17176
rect 36004 17172 36010 17174
rect 38285 17171 38351 17174
rect 200 17098 800 17128
rect 1577 17098 1643 17101
rect 200 17096 1643 17098
rect 200 17040 1582 17096
rect 1638 17040 1643 17096
rect 200 17038 1643 17040
rect 200 17008 800 17038
rect 1577 17035 1643 17038
rect 27061 17098 27127 17101
rect 28533 17098 28599 17101
rect 27061 17096 28599 17098
rect 27061 17040 27066 17096
rect 27122 17040 28538 17096
rect 28594 17040 28599 17096
rect 27061 17038 28599 17040
rect 27061 17035 27127 17038
rect 28533 17035 28599 17038
rect 36905 17098 36971 17101
rect 39200 17098 39800 17128
rect 36905 17096 39800 17098
rect 36905 17040 36910 17096
rect 36966 17040 39800 17096
rect 36905 17038 39800 17040
rect 36905 17035 36971 17038
rect 39200 17008 39800 17038
rect 25221 16962 25287 16965
rect 31753 16962 31819 16965
rect 25221 16960 31819 16962
rect 25221 16904 25226 16960
rect 25282 16904 31758 16960
rect 31814 16904 31819 16960
rect 25221 16902 31819 16904
rect 25221 16899 25287 16902
rect 31753 16899 31819 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 20805 16826 20871 16829
rect 24894 16826 24900 16828
rect 20805 16824 24900 16826
rect 20805 16768 20810 16824
rect 20866 16768 24900 16824
rect 20805 16766 24900 16768
rect 20805 16763 20871 16766
rect 24894 16764 24900 16766
rect 24964 16764 24970 16828
rect 30925 16826 30991 16829
rect 33225 16826 33291 16829
rect 30925 16824 33291 16826
rect 30925 16768 30930 16824
rect 30986 16768 33230 16824
rect 33286 16768 33291 16824
rect 30925 16766 33291 16768
rect 30925 16763 30991 16766
rect 33225 16763 33291 16766
rect 30782 16628 30788 16692
rect 30852 16690 30858 16692
rect 33317 16690 33383 16693
rect 30852 16688 33383 16690
rect 30852 16632 33322 16688
rect 33378 16632 33383 16688
rect 30852 16630 33383 16632
rect 30852 16628 30858 16630
rect 33317 16627 33383 16630
rect 29126 16492 29132 16556
rect 29196 16554 29202 16556
rect 31109 16554 31175 16557
rect 29196 16552 31175 16554
rect 29196 16496 31114 16552
rect 31170 16496 31175 16552
rect 29196 16494 31175 16496
rect 29196 16492 29202 16494
rect 31109 16491 31175 16494
rect 31886 16492 31892 16556
rect 31956 16554 31962 16556
rect 35249 16554 35315 16557
rect 31956 16552 35315 16554
rect 31956 16496 35254 16552
rect 35310 16496 35315 16552
rect 31956 16494 35315 16496
rect 31956 16492 31962 16494
rect 35249 16491 35315 16494
rect 30230 16356 30236 16420
rect 30300 16418 30306 16420
rect 34973 16418 35039 16421
rect 30300 16416 35039 16418
rect 30300 16360 34978 16416
rect 35034 16360 35039 16416
rect 30300 16358 35039 16360
rect 30300 16356 30306 16358
rect 34973 16355 35039 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 32254 16220 32260 16284
rect 32324 16282 32330 16284
rect 36445 16282 36511 16285
rect 32324 16280 36511 16282
rect 32324 16224 36450 16280
rect 36506 16224 36511 16280
rect 32324 16222 36511 16224
rect 32324 16220 32330 16222
rect 36445 16219 36511 16222
rect 20621 16146 20687 16149
rect 22645 16146 22711 16149
rect 20621 16144 22711 16146
rect 20621 16088 20626 16144
rect 20682 16088 22650 16144
rect 22706 16088 22711 16144
rect 20621 16086 22711 16088
rect 20621 16083 20687 16086
rect 22645 16083 22711 16086
rect 31017 16146 31083 16149
rect 36629 16146 36695 16149
rect 31017 16144 36695 16146
rect 31017 16088 31022 16144
rect 31078 16088 36634 16144
rect 36690 16088 36695 16144
rect 31017 16086 36695 16088
rect 31017 16083 31083 16086
rect 36629 16083 36695 16086
rect 22645 16010 22711 16013
rect 27981 16010 28047 16013
rect 22645 16008 28047 16010
rect 22645 15952 22650 16008
rect 22706 15952 27986 16008
rect 28042 15952 28047 16008
rect 22645 15950 28047 15952
rect 22645 15947 22711 15950
rect 27981 15947 28047 15950
rect 30741 16010 30807 16013
rect 33501 16010 33567 16013
rect 30741 16008 33567 16010
rect 30741 15952 30746 16008
rect 30802 15952 33506 16008
rect 33562 15952 33567 16008
rect 30741 15950 33567 15952
rect 30741 15947 30807 15950
rect 33501 15947 33567 15950
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 27654 15676 27660 15740
rect 27724 15738 27730 15740
rect 30925 15738 30991 15741
rect 27724 15736 30991 15738
rect 27724 15680 30930 15736
rect 30986 15680 30991 15736
rect 27724 15678 30991 15680
rect 27724 15676 27730 15678
rect 30925 15675 30991 15678
rect 35433 15738 35499 15741
rect 39200 15738 39800 15768
rect 35433 15736 39800 15738
rect 35433 15680 35438 15736
rect 35494 15680 39800 15736
rect 35433 15678 39800 15680
rect 35433 15675 35499 15678
rect 39200 15648 39800 15678
rect 34881 15602 34947 15605
rect 35750 15602 35756 15604
rect 34881 15600 35756 15602
rect 34881 15544 34886 15600
rect 34942 15544 35756 15600
rect 34881 15542 35756 15544
rect 34881 15539 34947 15542
rect 35750 15540 35756 15542
rect 35820 15540 35826 15604
rect 24710 15268 24716 15332
rect 24780 15330 24786 15332
rect 26509 15330 26575 15333
rect 24780 15328 26575 15330
rect 24780 15272 26514 15328
rect 26570 15272 26575 15328
rect 24780 15270 26575 15272
rect 24780 15268 24786 15270
rect 26509 15267 26575 15270
rect 31334 15268 31340 15332
rect 31404 15330 31410 15332
rect 33041 15330 33107 15333
rect 31404 15328 33107 15330
rect 31404 15272 33046 15328
rect 33102 15272 33107 15328
rect 31404 15270 33107 15272
rect 31404 15268 31410 15270
rect 33041 15267 33107 15270
rect 34646 15268 34652 15332
rect 34716 15330 34722 15332
rect 38009 15330 38075 15333
rect 34716 15328 38075 15330
rect 34716 15272 38014 15328
rect 38070 15272 38075 15328
rect 34716 15270 38075 15272
rect 34716 15268 34722 15270
rect 38009 15267 38075 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 34881 15194 34947 15197
rect 36302 15194 36308 15196
rect 34881 15192 36308 15194
rect 34881 15136 34886 15192
rect 34942 15136 36308 15192
rect 34881 15134 36308 15136
rect 34881 15131 34947 15134
rect 36302 15132 36308 15134
rect 36372 15194 36378 15196
rect 38929 15194 38995 15197
rect 36372 15192 38995 15194
rect 36372 15136 38934 15192
rect 38990 15136 38995 15192
rect 36372 15134 38995 15136
rect 36372 15132 36378 15134
rect 38929 15131 38995 15134
rect 38193 15058 38259 15061
rect 39200 15058 39800 15088
rect 38193 15056 39800 15058
rect 38193 15000 38198 15056
rect 38254 15000 39800 15056
rect 38193 14998 39800 15000
rect 38193 14995 38259 14998
rect 39200 14968 39800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 18505 14378 18571 14381
rect 34646 14378 34652 14380
rect 18505 14376 34652 14378
rect 18505 14320 18510 14376
rect 18566 14320 34652 14376
rect 18505 14318 34652 14320
rect 18505 14315 18571 14318
rect 34646 14316 34652 14318
rect 34716 14316 34722 14380
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 31518 13636 31524 13700
rect 31588 13698 31594 13700
rect 33685 13698 33751 13701
rect 39200 13698 39800 13728
rect 31588 13696 33751 13698
rect 31588 13640 33690 13696
rect 33746 13640 33751 13696
rect 31588 13638 33751 13640
rect 31588 13636 31594 13638
rect 33685 13635 33751 13638
rect 35390 13638 39800 13698
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 32857 13562 32923 13565
rect 32990 13562 32996 13564
rect 32857 13560 32996 13562
rect 32857 13504 32862 13560
rect 32918 13504 32996 13560
rect 32857 13502 32996 13504
rect 32857 13499 32923 13502
rect 32990 13500 32996 13502
rect 33060 13500 33066 13564
rect 32489 13426 32555 13429
rect 35390 13426 35450 13638
rect 39200 13608 39800 13638
rect 36169 13562 36235 13565
rect 36302 13562 36308 13564
rect 36169 13560 36308 13562
rect 36169 13504 36174 13560
rect 36230 13504 36308 13560
rect 36169 13502 36308 13504
rect 36169 13499 36235 13502
rect 36302 13500 36308 13502
rect 36372 13500 36378 13564
rect 32489 13424 35450 13426
rect 32489 13368 32494 13424
rect 32550 13368 35450 13424
rect 32489 13366 35450 13368
rect 32489 13363 32555 13366
rect 33133 13290 33199 13293
rect 36118 13290 36124 13292
rect 33133 13288 36124 13290
rect 33133 13232 33138 13288
rect 33194 13232 36124 13288
rect 33133 13230 36124 13232
rect 33133 13227 33199 13230
rect 36118 13228 36124 13230
rect 36188 13228 36194 13292
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 25998 12684 26004 12748
rect 26068 12746 26074 12748
rect 33685 12746 33751 12749
rect 26068 12744 33751 12746
rect 26068 12688 33690 12744
rect 33746 12688 33751 12744
rect 26068 12686 33751 12688
rect 26068 12684 26074 12686
rect 33685 12683 33751 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 36353 12474 36419 12477
rect 37457 12474 37523 12477
rect 36353 12472 37523 12474
rect 36353 12416 36358 12472
rect 36414 12416 37462 12472
rect 37518 12416 37523 12472
rect 36353 12414 37523 12416
rect 36353 12411 36419 12414
rect 37457 12411 37523 12414
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 32438 12276 32444 12340
rect 32508 12338 32514 12340
rect 33409 12338 33475 12341
rect 32508 12336 33475 12338
rect 32508 12280 33414 12336
rect 33470 12280 33475 12336
rect 32508 12278 33475 12280
rect 32508 12276 32514 12278
rect 33409 12275 33475 12278
rect 33910 12276 33916 12340
rect 33980 12338 33986 12340
rect 36261 12338 36327 12341
rect 33980 12336 36327 12338
rect 33980 12280 36266 12336
rect 36322 12280 36327 12336
rect 33980 12278 36327 12280
rect 33980 12276 33986 12278
rect 36261 12275 36327 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 34646 11868 34652 11932
rect 34716 11930 34722 11932
rect 37549 11930 37615 11933
rect 34716 11928 37615 11930
rect 34716 11872 37554 11928
rect 37610 11872 37615 11928
rect 34716 11870 37615 11872
rect 34716 11868 34722 11870
rect 37549 11867 37615 11870
rect 33726 11596 33732 11660
rect 33796 11658 33802 11660
rect 36261 11658 36327 11661
rect 33796 11656 36327 11658
rect 33796 11600 36266 11656
rect 36322 11600 36327 11656
rect 33796 11598 36327 11600
rect 33796 11596 33802 11598
rect 36261 11595 36327 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 31150 10916 31156 10980
rect 31220 10978 31226 10980
rect 34421 10978 34487 10981
rect 31220 10976 34487 10978
rect 31220 10920 34426 10976
rect 34482 10920 34487 10976
rect 31220 10918 34487 10920
rect 31220 10916 31226 10918
rect 34421 10915 34487 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 33174 10508 33180 10572
rect 33244 10570 33250 10572
rect 36721 10570 36787 10573
rect 33244 10568 36787 10570
rect 33244 10512 36726 10568
rect 36782 10512 36787 10568
rect 33244 10510 36787 10512
rect 33244 10508 33250 10510
rect 36721 10507 36787 10510
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1761 8938 1827 8941
rect 200 8936 1827 8938
rect 200 8880 1766 8936
rect 1822 8880 1827 8936
rect 200 8878 1827 8880
rect 200 8848 800 8878
rect 1761 8875 1827 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 38193 7578 38259 7581
rect 39200 7578 39800 7608
rect 38193 7576 39800 7578
rect 38193 7520 38198 7576
rect 38254 7520 39800 7576
rect 38193 7518 39800 7520
rect 38193 7515 38259 7518
rect 39200 7488 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1577 5538 1643 5541
rect 200 5536 1643 5538
rect 200 5480 1582 5536
rect 1638 5480 1643 5536
rect 200 5478 1643 5480
rect 200 5448 800 5478
rect 1577 5475 1643 5478
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 200 4178 800 4208
rect 1761 4178 1827 4181
rect 200 4176 1827 4178
rect 200 4120 1766 4176
rect 1822 4120 1827 4176
rect 200 4118 1827 4120
rect 200 4088 800 4118
rect 1761 4115 1827 4118
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 37457 3498 37523 3501
rect 39200 3498 39800 3528
rect 37457 3496 39800 3498
rect 37457 3440 37462 3496
rect 37518 3440 39800 3496
rect 37457 3438 39800 3440
rect 37457 3435 37523 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 35893 2684 35959 2685
rect 35893 2680 35940 2684
rect 36004 2682 36010 2684
rect 35893 2624 35898 2680
rect 35893 2620 35940 2624
rect 36004 2622 36050 2682
rect 36004 2620 36010 2622
rect 35893 2619 35959 2620
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 3141 2138 3207 2141
rect 200 2136 3207 2138
rect 200 2080 3146 2136
rect 3202 2080 3207 2136
rect 200 2078 3207 2080
rect 200 2048 800 2078
rect 3141 2075 3207 2078
rect 36813 2138 36879 2141
rect 39200 2138 39800 2168
rect 36813 2136 39800 2138
rect 36813 2080 36818 2136
rect 36874 2080 39800 2136
rect 36813 2078 39800 2080
rect 36813 2075 36879 2078
rect 39200 2048 39800 2078
rect 200 778 800 808
rect 1393 778 1459 781
rect 200 776 1459 778
rect 200 720 1398 776
rect 1454 720 1459 776
rect 200 718 1459 720
rect 200 688 800 718
rect 1393 715 1459 718
rect 38193 778 38259 781
rect 39200 778 39800 808
rect 38193 776 39800 778
rect 38193 720 38198 776
rect 38254 720 39800 776
rect 38193 718 39800 720
rect 38193 715 38259 718
rect 39200 688 39800 718
rect 37181 98 37247 101
rect 39200 98 39800 128
rect 37181 96 39800 98
rect 37181 40 37186 96
rect 37242 40 39800 96
rect 37181 38 39800 40
rect 37181 35 37247 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 35572 37300 35636 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 9444 36484 9508 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 33180 36544 33244 36548
rect 33180 36488 33194 36544
rect 33194 36488 33244 36544
rect 33180 36484 33244 36488
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 32444 36348 32508 36412
rect 29132 35940 29196 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 15700 34580 15764 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 33916 33764 33980 33828
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 34652 33356 34716 33420
rect 27660 33280 27724 33284
rect 27660 33224 27674 33280
rect 27674 33224 27724 33280
rect 27660 33220 27724 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 25452 32328 25516 32332
rect 25452 32272 25502 32328
rect 25502 32272 25516 32328
rect 25452 32268 25516 32272
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 25636 31996 25700 32060
rect 36308 31784 36372 31788
rect 36308 31728 36322 31784
rect 36322 31728 36372 31784
rect 36308 31724 36372 31728
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 34652 30968 34716 30972
rect 34652 30912 34666 30968
rect 34666 30912 34716 30968
rect 34652 30908 34716 30912
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 19380 30364 19444 30428
rect 24716 30364 24780 30428
rect 28764 30364 28828 30428
rect 30236 30364 30300 30428
rect 31892 30364 31956 30428
rect 21404 30228 21468 30292
rect 31524 29956 31588 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 9444 29820 9508 29884
rect 19380 29472 19444 29476
rect 19380 29416 19430 29472
rect 19430 29416 19444 29472
rect 19380 29412 19444 29416
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 26004 29140 26068 29204
rect 31340 29064 31404 29068
rect 31340 29008 31354 29064
rect 31354 29008 31404 29064
rect 31340 29004 31404 29008
rect 32260 29064 32324 29068
rect 32260 29008 32274 29064
rect 32274 29008 32324 29064
rect 32260 29004 32324 29008
rect 32996 29004 33060 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 34468 26344 34532 26348
rect 34468 26288 34482 26344
rect 34482 26288 34532 26344
rect 34468 26284 34532 26288
rect 23428 26148 23492 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 24900 25740 24964 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19380 25196 19444 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 30420 24924 30484 24988
rect 33732 24984 33796 24988
rect 33732 24928 33746 24984
rect 33746 24928 33796 24984
rect 33732 24924 33796 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 27844 23428 27908 23492
rect 35756 23428 35820 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 30052 23020 30116 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 15700 22612 15764 22676
rect 23612 22612 23676 22676
rect 19380 22400 19444 22404
rect 19380 22344 19394 22400
rect 19394 22344 19444 22400
rect 19380 22340 19444 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 23428 21932 23492 21996
rect 38148 21932 38212 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 21404 20572 21468 20636
rect 31156 20572 31220 20636
rect 30788 20496 30852 20500
rect 30788 20440 30802 20496
rect 30802 20440 30852 20496
rect 30788 20436 30852 20440
rect 38148 20360 38212 20364
rect 38148 20304 38198 20360
rect 38198 20304 38212 20360
rect 38148 20300 38212 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 30420 19892 30484 19956
rect 34652 19892 34716 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 23612 19348 23676 19412
rect 36308 19212 36372 19276
rect 30052 19076 30116 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 27844 18804 27908 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 25636 18124 25700 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 28764 17852 28828 17916
rect 35572 17580 35636 17644
rect 36124 17640 36188 17644
rect 36124 17584 36174 17640
rect 36174 17584 36188 17640
rect 36124 17580 36188 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 25452 17308 25516 17372
rect 35940 17172 36004 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 24900 16764 24964 16828
rect 30788 16628 30852 16692
rect 29132 16492 29196 16556
rect 31892 16492 31956 16556
rect 30236 16356 30300 16420
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 32260 16220 32324 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 27660 15676 27724 15740
rect 35756 15540 35820 15604
rect 24716 15268 24780 15332
rect 31340 15268 31404 15332
rect 34652 15268 34716 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 36308 15132 36372 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 34652 14316 34716 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 31524 13636 31588 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 32996 13500 33060 13564
rect 36308 13500 36372 13564
rect 36124 13228 36188 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 26004 12684 26068 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 32444 12276 32508 12340
rect 33916 12276 33980 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 34652 11868 34716 11932
rect 33732 11596 33796 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 31156 10916 31220 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 33180 10508 33244 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 35940 2680 36004 2684
rect 35940 2624 35954 2680
rect 35954 2624 36004 2680
rect 35940 2620 36004 2624
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 9443 36548 9509 36549
rect 9443 36484 9444 36548
rect 9508 36484 9509 36548
rect 9443 36483 9509 36484
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 9446 29885 9506 36483
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 33179 36548 33245 36549
rect 33179 36484 33180 36548
rect 33244 36484 33245 36548
rect 33179 36483 33245 36484
rect 32443 36412 32509 36413
rect 32443 36348 32444 36412
rect 32508 36348 32509 36412
rect 32443 36347 32509 36348
rect 29131 36004 29197 36005
rect 29131 35940 29132 36004
rect 29196 35940 29197 36004
rect 29131 35939 29197 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 15699 34644 15765 34645
rect 15699 34580 15700 34644
rect 15764 34580 15765 34644
rect 15699 34579 15765 34580
rect 9443 29884 9509 29885
rect 9443 29820 9444 29884
rect 9508 29820 9509 29884
rect 9443 29819 9509 29820
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 15702 22677 15762 34579
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 27659 33284 27725 33285
rect 27659 33220 27660 33284
rect 27724 33220 27725 33284
rect 27659 33219 27725 33220
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 25451 32332 25517 32333
rect 25451 32268 25452 32332
rect 25516 32268 25517 32332
rect 25451 32267 25517 32268
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19379 30428 19445 30429
rect 19379 30364 19380 30428
rect 19444 30364 19445 30428
rect 19379 30363 19445 30364
rect 19382 29477 19442 30363
rect 19379 29476 19445 29477
rect 19379 29412 19380 29476
rect 19444 29412 19445 29476
rect 19379 29411 19445 29412
rect 19568 29408 19888 30432
rect 24715 30428 24781 30429
rect 24715 30364 24716 30428
rect 24780 30364 24781 30428
rect 24715 30363 24781 30364
rect 21403 30292 21469 30293
rect 21403 30228 21404 30292
rect 21468 30228 21469 30292
rect 21403 30227 21469 30228
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19379 25260 19445 25261
rect 19379 25196 19380 25260
rect 19444 25196 19445 25260
rect 19379 25195 19445 25196
rect 15699 22676 15765 22677
rect 15699 22612 15700 22676
rect 15764 22612 15765 22676
rect 15699 22611 15765 22612
rect 19382 22405 19442 25195
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19379 22404 19445 22405
rect 19379 22340 19380 22404
rect 19444 22340 19445 22404
rect 19379 22339 19445 22340
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 21406 20637 21466 30227
rect 23427 26212 23493 26213
rect 23427 26148 23428 26212
rect 23492 26148 23493 26212
rect 23427 26147 23493 26148
rect 23430 21997 23490 26147
rect 23611 22676 23677 22677
rect 23611 22612 23612 22676
rect 23676 22612 23677 22676
rect 23611 22611 23677 22612
rect 23427 21996 23493 21997
rect 23427 21932 23428 21996
rect 23492 21932 23493 21996
rect 23427 21931 23493 21932
rect 21403 20636 21469 20637
rect 21403 20572 21404 20636
rect 21468 20572 21469 20636
rect 21403 20571 21469 20572
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 23614 19413 23674 22611
rect 23611 19412 23677 19413
rect 23611 19348 23612 19412
rect 23676 19348 23677 19412
rect 23611 19347 23677 19348
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 24718 15333 24778 30363
rect 24899 25804 24965 25805
rect 24899 25740 24900 25804
rect 24964 25740 24965 25804
rect 24899 25739 24965 25740
rect 24902 16829 24962 25739
rect 25454 17373 25514 32267
rect 25635 32060 25701 32061
rect 25635 31996 25636 32060
rect 25700 31996 25701 32060
rect 25635 31995 25701 31996
rect 25638 18189 25698 31995
rect 26003 29204 26069 29205
rect 26003 29140 26004 29204
rect 26068 29140 26069 29204
rect 26003 29139 26069 29140
rect 25635 18188 25701 18189
rect 25635 18124 25636 18188
rect 25700 18124 25701 18188
rect 25635 18123 25701 18124
rect 25451 17372 25517 17373
rect 25451 17308 25452 17372
rect 25516 17308 25517 17372
rect 25451 17307 25517 17308
rect 24899 16828 24965 16829
rect 24899 16764 24900 16828
rect 24964 16764 24965 16828
rect 24899 16763 24965 16764
rect 24715 15332 24781 15333
rect 24715 15268 24716 15332
rect 24780 15268 24781 15332
rect 24715 15267 24781 15268
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 26006 12749 26066 29139
rect 27662 15741 27722 33219
rect 28763 30428 28829 30429
rect 28763 30364 28764 30428
rect 28828 30364 28829 30428
rect 28763 30363 28829 30364
rect 27843 23492 27909 23493
rect 27843 23428 27844 23492
rect 27908 23428 27909 23492
rect 27843 23427 27909 23428
rect 27846 18869 27906 23427
rect 27843 18868 27909 18869
rect 27843 18804 27844 18868
rect 27908 18804 27909 18868
rect 27843 18803 27909 18804
rect 28766 17917 28826 30363
rect 28763 17916 28829 17917
rect 28763 17852 28764 17916
rect 28828 17852 28829 17916
rect 28763 17851 28829 17852
rect 29134 16557 29194 35939
rect 30235 30428 30301 30429
rect 30235 30364 30236 30428
rect 30300 30364 30301 30428
rect 30235 30363 30301 30364
rect 31891 30428 31957 30429
rect 31891 30364 31892 30428
rect 31956 30364 31957 30428
rect 31891 30363 31957 30364
rect 30051 23084 30117 23085
rect 30051 23020 30052 23084
rect 30116 23020 30117 23084
rect 30051 23019 30117 23020
rect 30054 19141 30114 23019
rect 30051 19140 30117 19141
rect 30051 19076 30052 19140
rect 30116 19076 30117 19140
rect 30051 19075 30117 19076
rect 29131 16556 29197 16557
rect 29131 16492 29132 16556
rect 29196 16492 29197 16556
rect 29131 16491 29197 16492
rect 30238 16421 30298 30363
rect 31523 30020 31589 30021
rect 31523 29956 31524 30020
rect 31588 29956 31589 30020
rect 31523 29955 31589 29956
rect 31339 29068 31405 29069
rect 31339 29004 31340 29068
rect 31404 29004 31405 29068
rect 31339 29003 31405 29004
rect 30419 24988 30485 24989
rect 30419 24924 30420 24988
rect 30484 24924 30485 24988
rect 30419 24923 30485 24924
rect 30422 19957 30482 24923
rect 31155 20636 31221 20637
rect 31155 20572 31156 20636
rect 31220 20572 31221 20636
rect 31155 20571 31221 20572
rect 30787 20500 30853 20501
rect 30787 20436 30788 20500
rect 30852 20436 30853 20500
rect 30787 20435 30853 20436
rect 30419 19956 30485 19957
rect 30419 19892 30420 19956
rect 30484 19892 30485 19956
rect 30419 19891 30485 19892
rect 30790 16693 30850 20435
rect 30787 16692 30853 16693
rect 30787 16628 30788 16692
rect 30852 16628 30853 16692
rect 30787 16627 30853 16628
rect 30235 16420 30301 16421
rect 30235 16356 30236 16420
rect 30300 16356 30301 16420
rect 30235 16355 30301 16356
rect 27659 15740 27725 15741
rect 27659 15676 27660 15740
rect 27724 15676 27725 15740
rect 27659 15675 27725 15676
rect 26003 12748 26069 12749
rect 26003 12684 26004 12748
rect 26068 12684 26069 12748
rect 26003 12683 26069 12684
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 31158 10981 31218 20571
rect 31342 15333 31402 29003
rect 31339 15332 31405 15333
rect 31339 15268 31340 15332
rect 31404 15268 31405 15332
rect 31339 15267 31405 15268
rect 31526 13701 31586 29955
rect 31894 16557 31954 30363
rect 32259 29068 32325 29069
rect 32259 29004 32260 29068
rect 32324 29004 32325 29068
rect 32259 29003 32325 29004
rect 31891 16556 31957 16557
rect 31891 16492 31892 16556
rect 31956 16492 31957 16556
rect 31891 16491 31957 16492
rect 32262 16285 32322 29003
rect 32259 16284 32325 16285
rect 32259 16220 32260 16284
rect 32324 16220 32325 16284
rect 32259 16219 32325 16220
rect 31523 13700 31589 13701
rect 31523 13636 31524 13700
rect 31588 13636 31589 13700
rect 31523 13635 31589 13636
rect 32446 12341 32506 36347
rect 32995 29068 33061 29069
rect 32995 29004 32996 29068
rect 33060 29004 33061 29068
rect 32995 29003 33061 29004
rect 32998 13565 33058 29003
rect 32995 13564 33061 13565
rect 32995 13500 32996 13564
rect 33060 13500 33061 13564
rect 32995 13499 33061 13500
rect 32443 12340 32509 12341
rect 32443 12276 32444 12340
rect 32508 12276 32509 12340
rect 32443 12275 32509 12276
rect 31155 10980 31221 10981
rect 31155 10916 31156 10980
rect 31220 10916 31221 10980
rect 31155 10915 31221 10916
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 33182 10573 33242 36483
rect 34928 36480 35248 37504
rect 35571 37364 35637 37365
rect 35571 37300 35572 37364
rect 35636 37300 35637 37364
rect 35571 37299 35637 37300
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 33915 33828 33981 33829
rect 33915 33764 33916 33828
rect 33980 33764 33981 33828
rect 33915 33763 33981 33764
rect 33731 24988 33797 24989
rect 33731 24924 33732 24988
rect 33796 24924 33797 24988
rect 33731 24923 33797 24924
rect 33734 11661 33794 24923
rect 33918 12341 33978 33763
rect 34651 33420 34717 33421
rect 34651 33356 34652 33420
rect 34716 33356 34717 33420
rect 34651 33355 34717 33356
rect 34654 30973 34714 33355
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34651 30972 34717 30973
rect 34651 30908 34652 30972
rect 34716 30908 34717 30972
rect 34651 30907 34717 30908
rect 34467 26348 34533 26349
rect 34467 26284 34468 26348
rect 34532 26284 34533 26348
rect 34467 26283 34533 26284
rect 34470 12450 34530 26283
rect 34654 19957 34714 30907
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34651 19956 34717 19957
rect 34651 19892 34652 19956
rect 34716 19892 34717 19956
rect 34651 19891 34717 19892
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 35574 17645 35634 37299
rect 36307 31788 36373 31789
rect 36307 31724 36308 31788
rect 36372 31724 36373 31788
rect 36307 31723 36373 31724
rect 35755 23492 35821 23493
rect 35755 23428 35756 23492
rect 35820 23428 35821 23492
rect 35755 23427 35821 23428
rect 35571 17644 35637 17645
rect 35571 17580 35572 17644
rect 35636 17580 35637 17644
rect 35571 17579 35637 17580
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34651 15332 34717 15333
rect 34651 15268 34652 15332
rect 34716 15268 34717 15332
rect 34651 15267 34717 15268
rect 34654 14381 34714 15267
rect 34928 14720 35248 15744
rect 35758 15605 35818 23427
rect 36310 19277 36370 31723
rect 38147 21996 38213 21997
rect 38147 21932 38148 21996
rect 38212 21932 38213 21996
rect 38147 21931 38213 21932
rect 38150 20365 38210 21931
rect 38147 20364 38213 20365
rect 38147 20300 38148 20364
rect 38212 20300 38213 20364
rect 38147 20299 38213 20300
rect 36307 19276 36373 19277
rect 36307 19212 36308 19276
rect 36372 19212 36373 19276
rect 36307 19211 36373 19212
rect 36123 17644 36189 17645
rect 36123 17580 36124 17644
rect 36188 17580 36189 17644
rect 36123 17579 36189 17580
rect 35939 17236 36005 17237
rect 35939 17172 35940 17236
rect 36004 17172 36005 17236
rect 35939 17171 36005 17172
rect 35755 15604 35821 15605
rect 35755 15540 35756 15604
rect 35820 15540 35821 15604
rect 35755 15539 35821 15540
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34651 14380 34717 14381
rect 34651 14316 34652 14380
rect 34716 14316 34717 14380
rect 34651 14315 34717 14316
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34470 12390 34714 12450
rect 33915 12340 33981 12341
rect 33915 12276 33916 12340
rect 33980 12276 33981 12340
rect 33915 12275 33981 12276
rect 34654 11933 34714 12390
rect 34651 11932 34717 11933
rect 34651 11868 34652 11932
rect 34716 11868 34717 11932
rect 34651 11867 34717 11868
rect 33731 11660 33797 11661
rect 33731 11596 33732 11660
rect 33796 11596 33797 11660
rect 33731 11595 33797 11596
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 33179 10572 33245 10573
rect 33179 10508 33180 10572
rect 33244 10508 33245 10572
rect 33179 10507 33245 10508
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35942 2685 36002 17171
rect 36126 13293 36186 17579
rect 36307 15196 36373 15197
rect 36307 15132 36308 15196
rect 36372 15132 36373 15196
rect 36307 15131 36373 15132
rect 36310 13565 36370 15131
rect 36307 13564 36373 13565
rect 36307 13500 36308 13564
rect 36372 13500 36373 13564
rect 36307 13499 36373 13500
rect 36123 13292 36189 13293
rect 36123 13228 36124 13292
rect 36188 13228 36189 13292
rect 36123 13227 36189 13228
rect 35939 2684 36005 2685
rect 35939 2620 35940 2684
rect 36004 2620 36005 2684
rect 35939 2619 36005 2620
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 37628 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 16744 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1667941163
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1667941163
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1667941163
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1667941163
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_20
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_28
timestamp 1667941163
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1667941163
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1667941163
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_186
timestamp 1667941163
transform 1 0 18216 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_198
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_210
timestamp 1667941163
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_348
timestamp 1667941163
transform 1 0 33120 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_360
timestamp 1667941163
transform 1 0 34224 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_372
timestamp 1667941163
transform 1 0 35328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_377
timestamp 1667941163
transform 1 0 35788 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_399
timestamp 1667941163
transform 1 0 37812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_16
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_385
timestamp 1667941163
transform 1 0 36524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1667941163
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1667941163
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1667941163
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_8
timestamp 1667941163
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1667941163
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_339
timestamp 1667941163
transform 1 0 32292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_343
timestamp 1667941163
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1667941163
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1667941163
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_314
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 1667941163
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 1667941163
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1667941163
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_75
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_87
timestamp 1667941163
transform 1 0 9108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1667941163
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1667941163
transform 1 0 17388 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_182
timestamp 1667941163
transform 1 0 17848 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_194
timestamp 1667941163
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_206
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_345
timestamp 1667941163
transform 1 0 32844 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1667941163
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_66
timestamp 1667941163
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_78
timestamp 1667941163
transform 1 0 8280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1667941163
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1667941163
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_200
timestamp 1667941163
transform 1 0 19504 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_212
timestamp 1667941163
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_264
timestamp 1667941163
transform 1 0 25392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1667941163
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_398
timestamp 1667941163
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1667941163
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1667941163
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1667941163
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_213
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1667941163
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1667941163
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_294
timestamp 1667941163
transform 1 0 28152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1667941163
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1667941163
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_66
timestamp 1667941163
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1667941163
transform 1 0 8280 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1667941163
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_101
timestamp 1667941163
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1667941163
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_197
timestamp 1667941163
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_209
timestamp 1667941163
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 1667941163
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_242
timestamp 1667941163
transform 1 0 23368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_254
timestamp 1667941163
transform 1 0 24472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_262
timestamp 1667941163
transform 1 0 25208 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_266
timestamp 1667941163
transform 1 0 25576 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1667941163
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1667941163
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_289
timestamp 1667941163
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_301
timestamp 1667941163
transform 1 0 28796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_313
timestamp 1667941163
transform 1 0 29900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1667941163
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_402
timestamp 1667941163
transform 1 0 38088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1667941163
transform 1 0 38456 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1667941163
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_94
timestamp 1667941163
transform 1 0 9752 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_106
timestamp 1667941163
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_118
timestamp 1667941163
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp 1667941163
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1667941163
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1667941163
transform 1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_213
timestamp 1667941163
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1667941163
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_223
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1667941163
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1667941163
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1667941163
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_271
timestamp 1667941163
transform 1 0 26036 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_283
timestamp 1667941163
transform 1 0 27140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_295
timestamp 1667941163
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_382
timestamp 1667941163
transform 1 0 36248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_397
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1667941163
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_140
timestamp 1667941163
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_152
timestamp 1667941163
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1667941163
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_180
timestamp 1667941163
transform 1 0 17664 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_204
timestamp 1667941163
transform 1 0 19872 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1667941163
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_263
timestamp 1667941163
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1667941163
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_304
timestamp 1667941163
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_316
timestamp 1667941163
transform 1 0 30176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1667941163
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_344
timestamp 1667941163
transform 1 0 32752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_356
timestamp 1667941163
transform 1 0 33856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_365
timestamp 1667941163
transform 1 0 34684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_374
timestamp 1667941163
transform 1 0 35512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_381
timestamp 1667941163
transform 1 0 36156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1667941163
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1667941163
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_90
timestamp 1667941163
transform 1 0 9384 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_102
timestamp 1667941163
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_114
timestamp 1667941163
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_126
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_169
timestamp 1667941163
transform 1 0 16652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_179
timestamp 1667941163
transform 1 0 17572 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1667941163
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_208
timestamp 1667941163
transform 1 0 20240 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_216
timestamp 1667941163
transform 1 0 20976 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1667941163
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_227
timestamp 1667941163
transform 1 0 21988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_235
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1667941163
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_339
timestamp 1667941163
transform 1 0 32292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_351
timestamp 1667941163
transform 1 0 33396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1667941163
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_371
timestamp 1667941163
transform 1 0 35236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_375
timestamp 1667941163
transform 1 0 35604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_382
timestamp 1667941163
transform 1 0 36248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_397
timestamp 1667941163
transform 1 0 37628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_94
timestamp 1667941163
transform 1 0 9752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1667941163
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1667941163
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_150
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1667941163
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1667941163
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_202
timestamp 1667941163
transform 1 0 19688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1667941163
transform 1 0 22540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1667941163
transform 1 0 24840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_269
timestamp 1667941163
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1667941163
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_355
timestamp 1667941163
transform 1 0 33764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_362
timestamp 1667941163
transform 1 0 34408 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_369
timestamp 1667941163
transform 1 0 35052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_376
timestamp 1667941163
transform 1 0 35696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_380
timestamp 1667941163
transform 1 0 36064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_398
timestamp 1667941163
transform 1 0 37720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_115
timestamp 1667941163
transform 1 0 11684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1667941163
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_126
timestamp 1667941163
transform 1 0 12696 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1667941163
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_208
timestamp 1667941163
transform 1 0 20240 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_220
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_232
timestamp 1667941163
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1667941163
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1667941163
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_287
timestamp 1667941163
transform 1 0 27508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_293
timestamp 1667941163
transform 1 0 28060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_297
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1667941163
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_353
timestamp 1667941163
transform 1 0 33580 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1667941163
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_374
timestamp 1667941163
transform 1 0 35512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_381
timestamp 1667941163
transform 1 0 36156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_388
timestamp 1667941163
transform 1 0 36800 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1667941163
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_66
timestamp 1667941163
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 1667941163
transform 1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1667941163
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_91
timestamp 1667941163
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_128
timestamp 1667941163
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1667941163
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1667941163
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1667941163
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_210
timestamp 1667941163
transform 1 0 20424 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1667941163
transform 1 0 22540 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_238
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_250
timestamp 1667941163
transform 1 0 24104 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1667941163
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_274
timestamp 1667941163
transform 1 0 26312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1667941163
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_356
timestamp 1667941163
transform 1 0 33856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_363
timestamp 1667941163
transform 1 0 34500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1667941163
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_377
timestamp 1667941163
transform 1 0 35788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1667941163
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_124
timestamp 1667941163
transform 1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1667941163
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_154
timestamp 1667941163
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1667941163
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_178
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1667941163
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_214
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_226
timestamp 1667941163
transform 1 0 21896 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_275
timestamp 1667941163
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_282
timestamp 1667941163
transform 1 0 27048 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_340
timestamp 1667941163
transform 1 0 32384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_347
timestamp 1667941163
transform 1 0 33028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_354
timestamp 1667941163
transform 1 0 33672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1667941163
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_370
timestamp 1667941163
transform 1 0 35144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_378
timestamp 1667941163
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_388
timestamp 1667941163
transform 1 0 36800 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_395
timestamp 1667941163
transform 1 0 37444 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1667941163
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1667941163
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1667941163
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1667941163
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_101
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1667941163
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_186
timestamp 1667941163
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_213
timestamp 1667941163
transform 1 0 20700 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_231
timestamp 1667941163
transform 1 0 22356 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_239
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_254
timestamp 1667941163
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_291
timestamp 1667941163
transform 1 0 27876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_297
timestamp 1667941163
transform 1 0 28428 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1667941163
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_310
timestamp 1667941163
transform 1 0 29624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_314
timestamp 1667941163
transform 1 0 29992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_320
timestamp 1667941163
transform 1 0 30544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1667941163
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_342
timestamp 1667941163
transform 1 0 32568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_351
timestamp 1667941163
transform 1 0 33396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_364
timestamp 1667941163
transform 1 0 34592 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_398
timestamp 1667941163
transform 1 0 37720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1667941163
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_185
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1667941163
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_229
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_235
timestamp 1667941163
transform 1 0 22724 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_272
timestamp 1667941163
transform 1 0 26128 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_293
timestamp 1667941163
transform 1 0 28060 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1667941163
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1667941163
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_340
timestamp 1667941163
transform 1 0 32384 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_348
timestamp 1667941163
transform 1 0 33120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_370
timestamp 1667941163
transform 1 0 35144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_378
timestamp 1667941163
transform 1 0 35880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1667941163
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_394
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_89
timestamp 1667941163
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_103
timestamp 1667941163
transform 1 0 10580 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_118
timestamp 1667941163
transform 1 0 11960 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1667941163
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_151
timestamp 1667941163
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_179
timestamp 1667941163
transform 1 0 17572 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_191
timestamp 1667941163
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_203
timestamp 1667941163
transform 1 0 19780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_234
timestamp 1667941163
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_248
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_296
timestamp 1667941163
transform 1 0 28336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_302
timestamp 1667941163
transform 1 0 28888 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1667941163
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1667941163
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1667941163
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1667941163
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_355
timestamp 1667941163
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_362
timestamp 1667941163
transform 1 0 34408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_366
timestamp 1667941163
transform 1 0 34776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_370
timestamp 1667941163
transform 1 0 35144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_377
timestamp 1667941163
transform 1 0 35788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_384
timestamp 1667941163
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_398
timestamp 1667941163
transform 1 0 37720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_114
timestamp 1667941163
transform 1 0 11592 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1667941163
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1667941163
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_146
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_170
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_182
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_206
timestamp 1667941163
transform 1 0 20056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_222
timestamp 1667941163
transform 1 0 21528 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_234
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1667941163
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_259
timestamp 1667941163
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_278
timestamp 1667941163
transform 1 0 26680 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_290
timestamp 1667941163
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1667941163
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_319
timestamp 1667941163
transform 1 0 30452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_326
timestamp 1667941163
transform 1 0 31096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_341
timestamp 1667941163
transform 1 0 32476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_351
timestamp 1667941163
transform 1 0 33396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1667941163
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_370
timestamp 1667941163
transform 1 0 35144 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_376
timestamp 1667941163
transform 1 0 35696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_386
timestamp 1667941163
transform 1 0 36616 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_397
timestamp 1667941163
transform 1 0 37628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_102
timestamp 1667941163
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1667941163
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1667941163
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_135
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_141
timestamp 1667941163
transform 1 0 14076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_192
timestamp 1667941163
transform 1 0 18768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_198
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1667941163
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_209
timestamp 1667941163
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1667941163
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_242
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_266
timestamp 1667941163
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1667941163
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1667941163
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_319
timestamp 1667941163
transform 1 0 30452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_325
timestamp 1667941163
transform 1 0 31004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_352
timestamp 1667941163
transform 1 0 33488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_365
timestamp 1667941163
transform 1 0 34684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_372
timestamp 1667941163
transform 1 0 35328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_379
timestamp 1667941163
transform 1 0 35972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1667941163
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_101
timestamp 1667941163
transform 1 0 10396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_113
timestamp 1667941163
transform 1 0 11500 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_126
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1667941163
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_180
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1667941163
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1667941163
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_223
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1667941163
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1667941163
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_261
timestamp 1667941163
transform 1 0 25116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_284
timestamp 1667941163
transform 1 0 27232 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_314
timestamp 1667941163
transform 1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_328
timestamp 1667941163
transform 1 0 31280 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_335
timestamp 1667941163
transform 1 0 31924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_342
timestamp 1667941163
transform 1 0 32568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_349
timestamp 1667941163
transform 1 0 33212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 1667941163
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_370
timestamp 1667941163
transform 1 0 35144 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_393
timestamp 1667941163
transform 1 0 37260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_397
timestamp 1667941163
transform 1 0 37628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1667941163
transform 1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_90
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1667941163
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 1667941163
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_145
timestamp 1667941163
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1667941163
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_192
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_209
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_231
timestamp 1667941163
transform 1 0 22356 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_239
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1667941163
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_292
timestamp 1667941163
transform 1 0 27968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1667941163
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_319
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_326
timestamp 1667941163
transform 1 0 31096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1667941163
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_354
timestamp 1667941163
transform 1 0 33672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_371
timestamp 1667941163
transform 1 0 35236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1667941163
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_404
timestamp 1667941163
transform 1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_35
timestamp 1667941163
transform 1 0 4324 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_47
timestamp 1667941163
transform 1 0 5428 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_59
timestamp 1667941163
transform 1 0 6532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_71
timestamp 1667941163
transform 1 0 7636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1667941163
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_111
timestamp 1667941163
transform 1 0 11316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_117
timestamp 1667941163
transform 1 0 11868 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_127
timestamp 1667941163
transform 1 0 12788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_223
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_231
timestamp 1667941163
transform 1 0 22356 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_281
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_329
timestamp 1667941163
transform 1 0 31372 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_343
timestamp 1667941163
transform 1 0 32660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1667941163
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_370
timestamp 1667941163
transform 1 0 35144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_384
timestamp 1667941163
transform 1 0 36432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_391
timestamp 1667941163
transform 1 0 37076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_398
timestamp 1667941163
transform 1 0 37720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_405
timestamp 1667941163
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1667941163
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1667941163
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1667941163
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_192
timestamp 1667941163
transform 1 0 18768 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_255
timestamp 1667941163
transform 1 0 24564 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_265
timestamp 1667941163
transform 1 0 25484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1667941163
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_299
timestamp 1667941163
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_306
timestamp 1667941163
transform 1 0 29256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_312
timestamp 1667941163
transform 1 0 29808 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_326
timestamp 1667941163
transform 1 0 31096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1667941163
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_356
timestamp 1667941163
transform 1 0 33856 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_363
timestamp 1667941163
transform 1 0 34500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_370
timestamp 1667941163
transform 1 0 35144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_377
timestamp 1667941163
transform 1 0 35788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_384
timestamp 1667941163
transform 1 0 36432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_398
timestamp 1667941163
transform 1 0 37720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_10
timestamp 1667941163
transform 1 0 2024 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1667941163
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1667941163
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1667941163
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_119
timestamp 1667941163
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_131
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_154
timestamp 1667941163
transform 1 0 15272 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_180
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_186
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1667941163
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_202
timestamp 1667941163
transform 1 0 19688 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_214
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_238
timestamp 1667941163
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_281
timestamp 1667941163
transform 1 0 26956 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1667941163
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_314
timestamp 1667941163
transform 1 0 29992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_328
timestamp 1667941163
transform 1 0 31280 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_335
timestamp 1667941163
transform 1 0 31924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_342
timestamp 1667941163
transform 1 0 32568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_349
timestamp 1667941163
transform 1 0 33212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1667941163
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_384
timestamp 1667941163
transform 1 0 36432 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_391
timestamp 1667941163
transform 1 0 37076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_398
timestamp 1667941163
transform 1 0 37720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 1667941163
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1667941163
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_138
timestamp 1667941163
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_150
timestamp 1667941163
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1667941163
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_180
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_192
timestamp 1667941163
transform 1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_236
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_248
timestamp 1667941163
transform 1 0 23920 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 1667941163
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_264
timestamp 1667941163
transform 1 0 25392 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_268
timestamp 1667941163
transform 1 0 25760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1667941163
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_298
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_308
timestamp 1667941163
transform 1 0 29440 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1667941163
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1667941163
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_360
timestamp 1667941163
transform 1 0 34224 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_377
timestamp 1667941163
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1667941163
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_128
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1667941163
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_182
timestamp 1667941163
transform 1 0 17848 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_225
timestamp 1667941163
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_274
timestamp 1667941163
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1667941163
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_332
timestamp 1667941163
transform 1 0 31648 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_376
timestamp 1667941163
transform 1 0 35696 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1667941163
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_63
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_70
timestamp 1667941163
transform 1 0 7544 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_82
timestamp 1667941163
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_94
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1667941163
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_191
timestamp 1667941163
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_215
timestamp 1667941163
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_242
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_257
timestamp 1667941163
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_262
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_270
timestamp 1667941163
transform 1 0 25944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1667941163
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_297
timestamp 1667941163
transform 1 0 28428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1667941163
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_311
timestamp 1667941163
transform 1 0 29716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_319
timestamp 1667941163
transform 1 0 30452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1667941163
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_342
timestamp 1667941163
transform 1 0 32568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_355
timestamp 1667941163
transform 1 0 33764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_369
timestamp 1667941163
transform 1 0 35052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_376
timestamp 1667941163
transform 1 0 35696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_383
timestamp 1667941163
transform 1 0 36340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1667941163
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1667941163
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1667941163
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_264
timestamp 1667941163
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1667941163
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_278
timestamp 1667941163
transform 1 0 26680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1667941163
transform 1 0 27600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_292
timestamp 1667941163
transform 1 0 27968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_329
timestamp 1667941163
transform 1 0 31372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_340
timestamp 1667941163
transform 1 0 32384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_348
timestamp 1667941163
transform 1 0 33120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_352
timestamp 1667941163
transform 1 0 33488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1667941163
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1667941163
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_373
timestamp 1667941163
transform 1 0 35420 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_380
timestamp 1667941163
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_387
timestamp 1667941163
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_391
timestamp 1667941163
transform 1 0 37076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_80
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_92
timestamp 1667941163
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1667941163
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1667941163
transform 1 0 23644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1667941163
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_263
timestamp 1667941163
transform 1 0 25300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_270
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1667941163
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 1667941163
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_309
timestamp 1667941163
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_321
timestamp 1667941163
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1667941163
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1667941163
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_398
timestamp 1667941163
transform 1 0 37720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_10
timestamp 1667941163
transform 1 0 2024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1667941163
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1667941163
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_90
timestamp 1667941163
transform 1 0 9384 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_122
timestamp 1667941163
transform 1 0 12328 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1667941163
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_156
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_175
timestamp 1667941163
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_257
timestamp 1667941163
transform 1 0 24748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_261
timestamp 1667941163
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1667941163
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_341
timestamp 1667941163
transform 1 0 32476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_387
timestamp 1667941163
transform 1 0 36708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_393
timestamp 1667941163
transform 1 0 37260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1667941163
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1667941163
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_77
timestamp 1667941163
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_102
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_106
timestamp 1667941163
transform 1 0 10856 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1667941163
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_151
timestamp 1667941163
transform 1 0 14996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_159
timestamp 1667941163
transform 1 0 15732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_255
timestamp 1667941163
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1667941163
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_270
timestamp 1667941163
transform 1 0 25944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_303
timestamp 1667941163
transform 1 0 28980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_311
timestamp 1667941163
transform 1 0 29716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1667941163
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_362
timestamp 1667941163
transform 1 0 34408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1667941163
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_95
timestamp 1667941163
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_107
timestamp 1667941163
transform 1 0 10948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_116
timestamp 1667941163
transform 1 0 11776 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1667941163
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_160
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_172
timestamp 1667941163
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_230
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_283
timestamp 1667941163
transform 1 0 27140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_295
timestamp 1667941163
transform 1 0 28244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_322
timestamp 1667941163
transform 1 0 30728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1667941163
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1667941163
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_388
timestamp 1667941163
transform 1 0 36800 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_399
timestamp 1667941163
transform 1 0 37812 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_124
timestamp 1667941163
transform 1 0 12512 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_132
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_136
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_148
timestamp 1667941163
transform 1 0 14720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1667941163
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1667941163
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_241
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_265
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_308
timestamp 1667941163
transform 1 0 29440 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1667941163
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_398
timestamp 1667941163
transform 1 0 37720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1667941163
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_68
timestamp 1667941163
transform 1 0 7360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_95
timestamp 1667941163
transform 1 0 9844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_107
timestamp 1667941163
transform 1 0 10948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_111
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1667941163
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_122
timestamp 1667941163
transform 1 0 12328 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_129
timestamp 1667941163
transform 1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1667941163
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1667941163
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_158
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_170
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_182
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_205
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1667941163
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_238
timestamp 1667941163
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_264
timestamp 1667941163
transform 1 0 25392 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_276
timestamp 1667941163
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_288
timestamp 1667941163
transform 1 0 27600 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_300
timestamp 1667941163
transform 1 0 28704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_315
timestamp 1667941163
transform 1 0 30084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_336
timestamp 1667941163
transform 1 0 32016 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1667941163
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_387
timestamp 1667941163
transform 1 0 36708 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1667941163
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_95
timestamp 1667941163
transform 1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_99
timestamp 1667941163
transform 1 0 10212 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1667941163
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1667941163
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_154
timestamp 1667941163
transform 1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_233
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1667941163
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1667941163
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_304
timestamp 1667941163
transform 1 0 29072 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1667941163
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_359
timestamp 1667941163
transform 1 0 34132 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_371
timestamp 1667941163
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_383
timestamp 1667941163
transform 1 0 36340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_61
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 1667941163
transform 1 0 7176 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_95
timestamp 1667941163
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_122
timestamp 1667941163
transform 1 0 12328 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1667941163
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1667941163
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1667941163
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1667941163
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_222
timestamp 1667941163
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_275
timestamp 1667941163
transform 1 0 26404 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_287
timestamp 1667941163
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1667941163
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1667941163
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1667941163
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_396
timestamp 1667941163
transform 1 0 37536 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_399
timestamp 1667941163
transform 1 0 37812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1667941163
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1667941163
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_77
timestamp 1667941163
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1667941163
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_133
timestamp 1667941163
transform 1 0 13340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1667941163
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_153
timestamp 1667941163
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1667941163
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_194
timestamp 1667941163
transform 1 0 18952 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1667941163
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_238
timestamp 1667941163
transform 1 0 23000 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_250
timestamp 1667941163
transform 1 0 24104 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_262
timestamp 1667941163
transform 1 0 25208 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1667941163
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_299
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_323
timestamp 1667941163
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_359
timestamp 1667941163
transform 1 0 34132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_401
timestamp 1667941163
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1667941163
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_112
timestamp 1667941163
transform 1 0 11408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_124
timestamp 1667941163
transform 1 0 12512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_132
timestamp 1667941163
transform 1 0 13248 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_152
timestamp 1667941163
transform 1 0 15088 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_171
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1667941163
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_226
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_230
timestamp 1667941163
transform 1 0 22264 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_278
timestamp 1667941163
transform 1 0 26680 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_290
timestamp 1667941163
transform 1 0 27784 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_302
timestamp 1667941163
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1667941163
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_340
timestamp 1667941163
transform 1 0 32384 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_352
timestamp 1667941163
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_387
timestamp 1667941163
transform 1 0 36708 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_404
timestamp 1667941163
transform 1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_87
timestamp 1667941163
transform 1 0 9108 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_91
timestamp 1667941163
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1667941163
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1667941163
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_128
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_139
timestamp 1667941163
transform 1 0 13892 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_151
timestamp 1667941163
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_208
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1667941163
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_250
timestamp 1667941163
transform 1 0 24104 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1667941163
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_304
timestamp 1667941163
transform 1 0 29072 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1667941163
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_365
timestamp 1667941163
transform 1 0 34684 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_377
timestamp 1667941163
transform 1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1667941163
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1667941163
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_103
timestamp 1667941163
transform 1 0 10580 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_115
timestamp 1667941163
transform 1 0 11684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_125
timestamp 1667941163
transform 1 0 12604 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_146
timestamp 1667941163
transform 1 0 14536 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_155
timestamp 1667941163
transform 1 0 15364 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_172
timestamp 1667941163
transform 1 0 16928 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_184
timestamp 1667941163
transform 1 0 18032 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1667941163
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_331
timestamp 1667941163
transform 1 0 31556 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1667941163
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_387
timestamp 1667941163
transform 1 0 36708 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_395
timestamp 1667941163
transform 1 0 37444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_399
timestamp 1667941163
transform 1 0 37812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1667941163
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_65
timestamp 1667941163
transform 1 0 7084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_72
timestamp 1667941163
transform 1 0 7728 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_79
timestamp 1667941163
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_91
timestamp 1667941163
transform 1 0 9476 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_101
timestamp 1667941163
transform 1 0 10396 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_128
timestamp 1667941163
transform 1 0 12880 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_132
timestamp 1667941163
transform 1 0 13248 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1667941163
transform 1 0 13616 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_185
timestamp 1667941163
transform 1 0 18124 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_209
timestamp 1667941163
transform 1 0 20332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1667941163
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_233
timestamp 1667941163
transform 1 0 22540 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_257
timestamp 1667941163
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1667941163
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1667941163
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_287
timestamp 1667941163
transform 1 0 27508 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_308
timestamp 1667941163
transform 1 0 29440 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_320
timestamp 1667941163
transform 1 0 30544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1667941163
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_397
timestamp 1667941163
transform 1 0 37628 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_401
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_59
timestamp 1667941163
transform 1 0 6532 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_63
timestamp 1667941163
transform 1 0 6900 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_71
timestamp 1667941163
transform 1 0 7636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1667941163
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_90
timestamp 1667941163
transform 1 0 9384 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_98
timestamp 1667941163
transform 1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_104
timestamp 1667941163
transform 1 0 10672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_116
timestamp 1667941163
transform 1 0 11776 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1667941163
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1667941163
transform 1 0 13064 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_134
timestamp 1667941163
transform 1 0 13432 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_161
timestamp 1667941163
transform 1 0 15916 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_183
timestamp 1667941163
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_236
timestamp 1667941163
transform 1 0 22816 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1667941163
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_276
timestamp 1667941163
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1667941163
transform 1 0 27600 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_292
timestamp 1667941163
transform 1 0 27968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1667941163
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_325
timestamp 1667941163
transform 1 0 31004 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_346
timestamp 1667941163
transform 1 0 32936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1667941163
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_388
timestamp 1667941163
transform 1 0 36800 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_394
timestamp 1667941163
transform 1 0 37352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_398
timestamp 1667941163
transform 1 0 37720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1667941163
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_96
timestamp 1667941163
transform 1 0 9936 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_103
timestamp 1667941163
transform 1 0 10580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_124
timestamp 1667941163
transform 1 0 12512 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_131
timestamp 1667941163
transform 1 0 13156 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1667941163
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_142
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1667941163
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_207
timestamp 1667941163
transform 1 0 20148 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_259
timestamp 1667941163
transform 1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1667941163
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1667941163
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_69
timestamp 1667941163
transform 1 0 7452 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1667941163
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_92
timestamp 1667941163
transform 1 0 9568 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_104
timestamp 1667941163
transform 1 0 10672 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1667941163
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_151
timestamp 1667941163
transform 1 0 14996 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_164
timestamp 1667941163
transform 1 0 16192 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_176
timestamp 1667941163
transform 1 0 17296 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1667941163
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_219
timestamp 1667941163
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_231
timestamp 1667941163
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1667941163
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_275
timestamp 1667941163
transform 1 0 26404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_322
timestamp 1667941163
transform 1 0 30728 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_328
timestamp 1667941163
transform 1 0 31280 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_349
timestamp 1667941163
transform 1 0 33212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 1667941163
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_387
timestamp 1667941163
transform 1 0 36708 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_394
timestamp 1667941163
transform 1 0 37352 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_400
timestamp 1667941163
transform 1 0 37904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_96
timestamp 1667941163
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_119
timestamp 1667941163
transform 1 0 12052 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_126
timestamp 1667941163
transform 1 0 12696 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_130
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_134
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_174
timestamp 1667941163
transform 1 0 17112 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_207
timestamp 1667941163
transform 1 0 20148 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1667941163
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1667941163
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_303
timestamp 1667941163
transform 1 0 28980 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_311
timestamp 1667941163
transform 1 0 29716 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_353
timestamp 1667941163
transform 1 0 33580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1667941163
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_73
timestamp 1667941163
transform 1 0 7820 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_100
timestamp 1667941163
transform 1 0 10304 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_113
timestamp 1667941163
transform 1 0 11500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_120
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_154
timestamp 1667941163
transform 1 0 15272 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_168
timestamp 1667941163
transform 1 0 16560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_172
timestamp 1667941163
transform 1 0 16928 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_215
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_239
timestamp 1667941163
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_276
timestamp 1667941163
transform 1 0 26496 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_284
timestamp 1667941163
transform 1 0 27232 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1667941163
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_342
timestamp 1667941163
transform 1 0 32568 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_350
timestamp 1667941163
transform 1 0 33304 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1667941163
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_387
timestamp 1667941163
transform 1 0 36708 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1667941163
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_77
timestamp 1667941163
transform 1 0 8188 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_82
timestamp 1667941163
transform 1 0 8648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_89
timestamp 1667941163
transform 1 0 9292 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_96
timestamp 1667941163
transform 1 0 9936 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_103
timestamp 1667941163
transform 1 0 10580 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_118
timestamp 1667941163
transform 1 0 11960 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_126
timestamp 1667941163
transform 1 0 12696 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_131
timestamp 1667941163
transform 1 0 13156 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_138
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_155
timestamp 1667941163
transform 1 0 15364 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_185
timestamp 1667941163
transform 1 0 18124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_207
timestamp 1667941163
transform 1 0 20148 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_260
timestamp 1667941163
transform 1 0 25024 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_267
timestamp 1667941163
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_304
timestamp 1667941163
transform 1 0 29072 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1667941163
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_360
timestamp 1667941163
transform 1 0 34224 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_372
timestamp 1667941163
transform 1 0 35328 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_384
timestamp 1667941163
transform 1 0 36432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1667941163
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_399
timestamp 1667941163
transform 1 0 37812 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_62
timestamp 1667941163
transform 1 0 6808 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_70
timestamp 1667941163
transform 1 0 7544 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_74
timestamp 1667941163
transform 1 0 7912 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1667941163
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_92
timestamp 1667941163
transform 1 0 9568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1667941163
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_103
timestamp 1667941163
transform 1 0 10580 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_107
timestamp 1667941163
transform 1 0 10948 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_114
timestamp 1667941163
transform 1 0 11592 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_127
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1667941163
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_150
timestamp 1667941163
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1667941163
transform 1 0 15272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1667941163
transform 1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_171
timestamp 1667941163
transform 1 0 16836 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_175
timestamp 1667941163
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_187
timestamp 1667941163
transform 1 0 18308 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1667941163
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_224
timestamp 1667941163
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_276
timestamp 1667941163
transform 1 0 26496 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_291
timestamp 1667941163
transform 1 0 27876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1667941163
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_383
timestamp 1667941163
transform 1 0 36340 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_85
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_89
timestamp 1667941163
transform 1 0 9292 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1667941163
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_124
timestamp 1667941163
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_131
timestamp 1667941163
transform 1 0 13156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_139
timestamp 1667941163
transform 1 0 13892 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_143
timestamp 1667941163
transform 1 0 14260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_153
timestamp 1667941163
transform 1 0 15180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1667941163
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_210
timestamp 1667941163
transform 1 0 20424 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1667941163
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_233
timestamp 1667941163
transform 1 0 22540 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_238
timestamp 1667941163
transform 1 0 23000 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1667941163
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1667941163
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_288
timestamp 1667941163
transform 1 0 27600 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_300
timestamp 1667941163
transform 1 0 28704 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_312
timestamp 1667941163
transform 1 0 29808 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_324
timestamp 1667941163
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_346
timestamp 1667941163
transform 1 0 32936 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_358
timestamp 1667941163
transform 1 0 34040 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_366
timestamp 1667941163
transform 1 0 34776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1667941163
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1667941163
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_69
timestamp 1667941163
transform 1 0 7452 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_91
timestamp 1667941163
transform 1 0 9476 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_98
timestamp 1667941163
transform 1 0 10120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_105
timestamp 1667941163
transform 1 0 10764 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_112
timestamp 1667941163
transform 1 0 11408 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_129
timestamp 1667941163
transform 1 0 12972 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1667941163
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_154
timestamp 1667941163
transform 1 0 15272 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_160
timestamp 1667941163
transform 1 0 15824 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_170
timestamp 1667941163
transform 1 0 16744 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_219
timestamp 1667941163
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_231
timestamp 1667941163
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1667941163
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_276
timestamp 1667941163
transform 1 0 26496 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_288
timestamp 1667941163
transform 1 0 27600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1667941163
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1667941163
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1667941163
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_358
timestamp 1667941163
transform 1 0 34040 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1667941163
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_387
timestamp 1667941163
transform 1 0 36708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_393
timestamp 1667941163
transform 1 0 37260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_397
timestamp 1667941163
transform 1 0 37628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_64
timestamp 1667941163
transform 1 0 6992 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_76
timestamp 1667941163
transform 1 0 8096 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_83
timestamp 1667941163
transform 1 0 8740 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_94
timestamp 1667941163
transform 1 0 9752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_101
timestamp 1667941163
transform 1 0 10396 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1667941163
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_124
timestamp 1667941163
transform 1 0 12512 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_133
timestamp 1667941163
transform 1 0 13340 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_146
timestamp 1667941163
transform 1 0 14536 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1667941163
transform 1 0 15180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1667941163
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_176
timestamp 1667941163
transform 1 0 17296 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_184
timestamp 1667941163
transform 1 0 18032 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_206
timestamp 1667941163
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1667941163
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_257
timestamp 1667941163
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1667941163
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_342
timestamp 1667941163
transform 1 0 32568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_366
timestamp 1667941163
transform 1 0 34776 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_377
timestamp 1667941163
transform 1 0 35788 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_384
timestamp 1667941163
transform 1 0 36432 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_94
timestamp 1667941163
transform 1 0 9752 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_101
timestamp 1667941163
transform 1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_108
timestamp 1667941163
transform 1 0 11040 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_115
timestamp 1667941163
transform 1 0 11684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_128
timestamp 1667941163
transform 1 0 12880 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_137
timestamp 1667941163
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1667941163
transform 1 0 14444 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_149
timestamp 1667941163
transform 1 0 14812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_162
timestamp 1667941163
transform 1 0 16008 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_169
timestamp 1667941163
transform 1 0 16652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_181
timestamp 1667941163
transform 1 0 17756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1667941163
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_229
timestamp 1667941163
transform 1 0 22172 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1667941163
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1667941163
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1667941163
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_325
timestamp 1667941163
transform 1 0 31004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_335
timestamp 1667941163
transform 1 0 31924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_343
timestamp 1667941163
transform 1 0 32660 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_355
timestamp 1667941163
transform 1 0 33764 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1667941163
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_380
timestamp 1667941163
transform 1 0 36064 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_395
timestamp 1667941163
transform 1 0 37444 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_399
timestamp 1667941163
transform 1 0 37812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_16
timestamp 1667941163
transform 1 0 2576 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_28
timestamp 1667941163
transform 1 0 3680 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_40
timestamp 1667941163
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1667941163
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_77
timestamp 1667941163
transform 1 0 8188 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_89
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_98
timestamp 1667941163
transform 1 0 10120 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_106
timestamp 1667941163
transform 1 0 10856 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1667941163
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_124
timestamp 1667941163
transform 1 0 12512 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_132
timestamp 1667941163
transform 1 0 13248 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1667941163
transform 1 0 14168 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_178
timestamp 1667941163
transform 1 0 17480 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_190
timestamp 1667941163
transform 1 0 18584 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_248
timestamp 1667941163
transform 1 0 23920 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_347
timestamp 1667941163
transform 1 0 33028 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1667941163
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_379
timestamp 1667941163
transform 1 0 35972 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_383
timestamp 1667941163
transform 1 0 36340 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1667941163
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_8
timestamp 1667941163
transform 1 0 1840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1667941163
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_36
timestamp 1667941163
transform 1 0 4416 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_48
timestamp 1667941163
transform 1 0 5520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_56
timestamp 1667941163
transform 1 0 6256 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_62
timestamp 1667941163
transform 1 0 6808 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_73
timestamp 1667941163
transform 1 0 7820 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_95
timestamp 1667941163
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_102
timestamp 1667941163
transform 1 0 10488 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_106
timestamp 1667941163
transform 1 0 10856 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_110
timestamp 1667941163
transform 1 0 11224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_117
timestamp 1667941163
transform 1 0 11868 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_124
timestamp 1667941163
transform 1 0 12512 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_131
timestamp 1667941163
transform 1 0 13156 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_158
timestamp 1667941163
transform 1 0 15640 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1667941163
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_227
timestamp 1667941163
transform 1 0 21988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_239
timestamp 1667941163
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_279
timestamp 1667941163
transform 1 0 26772 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_294
timestamp 1667941163
transform 1 0 28152 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1667941163
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_322
timestamp 1667941163
transform 1 0 30728 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_328
timestamp 1667941163
transform 1 0 31280 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_338
timestamp 1667941163
transform 1 0 32200 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1667941163
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_370
timestamp 1667941163
transform 1 0 35144 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_378
timestamp 1667941163
transform 1 0 35880 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_383
timestamp 1667941163
transform 1 0 36340 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_390
timestamp 1667941163
transform 1 0 36984 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_18
timestamp 1667941163
transform 1 0 2760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_22
timestamp 1667941163
transform 1 0 3128 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_26
timestamp 1667941163
transform 1 0 3496 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_38
timestamp 1667941163
transform 1 0 4600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_50
timestamp 1667941163
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_63
timestamp 1667941163
transform 1 0 6900 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_67
timestamp 1667941163
transform 1 0 7268 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_84
timestamp 1667941163
transform 1 0 8832 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_92
timestamp 1667941163
transform 1 0 9568 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_97
timestamp 1667941163
transform 1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1667941163
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_119
timestamp 1667941163
transform 1 0 12052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_131
timestamp 1667941163
transform 1 0 13156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_139
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_144
timestamp 1667941163
transform 1 0 14352 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_151
timestamp 1667941163
transform 1 0 14996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_158
timestamp 1667941163
transform 1 0 15640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_162
timestamp 1667941163
transform 1 0 16008 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_180
timestamp 1667941163
transform 1 0 17664 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_184
timestamp 1667941163
transform 1 0 18032 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_206
timestamp 1667941163
transform 1 0 20056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1667941163
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_257
timestamp 1667941163
transform 1 0 24748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1667941163
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_288
timestamp 1667941163
transform 1 0 27600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_313
timestamp 1667941163
transform 1 0 29900 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_320
timestamp 1667941163
transform 1 0 30544 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_324
timestamp 1667941163
transform 1 0 30912 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1667941163
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_342
timestamp 1667941163
transform 1 0 32568 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_354
timestamp 1667941163
transform 1 0 33672 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_366
timestamp 1667941163
transform 1 0 34776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_370
timestamp 1667941163
transform 1 0 35144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_377
timestamp 1667941163
transform 1 0 35788 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_12
timestamp 1667941163
transform 1 0 2208 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_34
timestamp 1667941163
transform 1 0 4232 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_46
timestamp 1667941163
transform 1 0 5336 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_50
timestamp 1667941163
transform 1 0 5704 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_54
timestamp 1667941163
transform 1 0 6072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_61
timestamp 1667941163
transform 1 0 6716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_68
timestamp 1667941163
transform 1 0 7360 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_75
timestamp 1667941163
transform 1 0 8004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_92
timestamp 1667941163
transform 1 0 9568 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_96
timestamp 1667941163
transform 1 0 9936 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_100
timestamp 1667941163
transform 1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_117
timestamp 1667941163
transform 1 0 11868 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_125
timestamp 1667941163
transform 1 0 12604 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_135
timestamp 1667941163
transform 1 0 13524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_152
timestamp 1667941163
transform 1 0 15088 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_182
timestamp 1667941163
transform 1 0 17848 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1667941163
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_223
timestamp 1667941163
transform 1 0 21620 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1667941163
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_275
timestamp 1667941163
transform 1 0 26404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_299
timestamp 1667941163
transform 1 0 28612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1667941163
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_334
timestamp 1667941163
transform 1 0 31832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_358
timestamp 1667941163
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1667941163
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_392
timestamp 1667941163
transform 1 0 37168 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_18
timestamp 1667941163
transform 1 0 2760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_32
timestamp 1667941163
transform 1 0 4048 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_36
timestamp 1667941163
transform 1 0 4416 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_40
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_63
timestamp 1667941163
transform 1 0 6900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_67
timestamp 1667941163
transform 1 0 7268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_74
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_82
timestamp 1667941163
transform 1 0 8648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_89
timestamp 1667941163
transform 1 0 9292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_96
timestamp 1667941163
transform 1 0 9936 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_103
timestamp 1667941163
transform 1 0 10580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_123
timestamp 1667941163
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_135
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_140
timestamp 1667941163
transform 1 0 13984 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_148
timestamp 1667941163
transform 1 0 14720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1667941163
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1667941163
transform 1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_271
timestamp 1667941163
transform 1 0 26036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1667941163
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1667941163
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_311
timestamp 1667941163
transform 1 0 29716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_318
timestamp 1667941163
transform 1 0 30360 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_327
timestamp 1667941163
transform 1 0 31188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_343
timestamp 1667941163
transform 1 0 32660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_351
timestamp 1667941163
transform 1 0 33396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_358
timestamp 1667941163
transform 1 0 34040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_383
timestamp 1667941163
transform 1 0 36340 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1667941163
transform 1 0 9936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_103
timestamp 1667941163
transform 1 0 10580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_152
timestamp 1667941163
transform 1 0 15088 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_184
timestamp 1667941163
transform 1 0 18032 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_190
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 1667941163
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1667941163
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1667941163
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_257
timestamp 1667941163
transform 1 0 24748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1667941163
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 28980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 30176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0399_
timestamp 1667941163
transform 1 0 30360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0400_
timestamp 1667941163
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 22724 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 17020 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0403_
timestamp 1667941163
transform 1 0 32292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 26680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0406_
timestamp 1667941163
transform 1 0 31464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 10304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 11684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0412_
timestamp 1667941163
transform 1 0 10120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0413_
timestamp 1667941163
transform 1 0 8464 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 9752 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0415_
timestamp 1667941163
transform 1 0 14536 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 10672 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0418_
timestamp 1667941163
transform 1 0 10212 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0419_
timestamp 1667941163
transform 1 0 9476 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0420_
timestamp 1667941163
transform 1 0 31464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0421_
timestamp 1667941163
transform 1 0 12144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 25392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 11500 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0424_
timestamp 1667941163
transform 1 0 19872 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0425_
timestamp 1667941163
transform 1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0426_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 35512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0430_
timestamp 1667941163
transform 1 0 14904 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 32936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 35144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0433_
timestamp 1667941163
transform 1 0 25116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 34132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0437_
timestamp 1667941163
transform 1 0 36064 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0438_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0439_
timestamp 1667941163
transform 1 0 32292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0442_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0443_
timestamp 1667941163
transform 1 0 32292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1667941163
transform 1 0 15640 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 14904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1667941163
transform 1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 29532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 22264 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1667941163
transform 1 0 29808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 3220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 2300 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 6716 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1667941163
transform 1 0 33212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 35052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0459_
timestamp 1667941163
transform 1 0 32292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462_
timestamp 1667941163
transform 1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0464_
timestamp 1667941163
transform 1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0465_
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 31648 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 17112 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1667941163
transform 1 0 13340 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1667941163
transform 1 0 20516 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 16376 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 9016 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1667941163
transform 1 0 9292 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 7728 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 18216 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 14904 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 32660 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 26956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 25024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 28244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 14720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 14904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 21160 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 13800 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 15732 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 10304 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 12420 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 6808 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 8280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0508_
timestamp 1667941163
transform 1 0 6900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0509_
timestamp 1667941163
transform 1 0 8464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 6624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 27968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0515_
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0520_
timestamp 1667941163
transform 1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 8372 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 8280 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 4508 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 6532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 9016 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 12880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0529_
timestamp 1667941163
transform 1 0 9200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 11776 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 19780 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform 1 0 12420 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 12788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0538_
timestamp 1667941163
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 19780 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 28520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 15548 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 14996 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 8372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 11040 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1667941163
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 8280 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 36708 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 34132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform 1 0 33396 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 34040 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 37076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 37444 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 32936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1667941163
transform 1 0 31464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform 1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 34776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 34132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 35328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 35880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 34132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 34132 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 33764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 36800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 15456 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 36156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 35512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 13524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 12880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 13432 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 35972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 34408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 10948 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 14996 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 25484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 34040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 34224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 9844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 7176 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 37720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 32292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 36156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 32476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 33488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 32016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 37352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0631_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 28796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 7820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 9200 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 9108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 6440 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 11040 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0648_
timestamp 1667941163
transform 1 0 12788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 16928 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 34132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 35236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 33856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 8372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 36156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 7636 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 36156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 35236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 37720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 27324 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 25760 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 36708 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 10304 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 25300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 36708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 37076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 8372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 36616 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 6992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 13064 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 11408 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 17204 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 7544 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 35512 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 9752 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0703_
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 13524 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0713_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0714_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25392 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0715_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 35512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 35696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 30360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 10948 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 13524 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 33580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 37168 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 36708 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0726_
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 35512 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 10948 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 30084 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 32752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 36616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 31556 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0737_
timestamp 1667941163
transform 1 0 27968 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 33580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 28336 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 37720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 36340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 37444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 36616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0748_
timestamp 1667941163
transform 1 0 28060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 26404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 33580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 22908 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 30360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 26036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 23736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 23552 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0759_
timestamp 1667941163
transform 1 0 21160 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 15364 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 12880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 14352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 21988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 11592 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 12880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 13524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0770_
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 15088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 32936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 32108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 26128 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 12788 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 14352 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0781_
timestamp 1667941163
transform 1 0 27508 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 11868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 31004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 33304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 37444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 36432 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 36064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0792_
timestamp 1667941163
transform 1 0 22540 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 32936 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 32292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 13524 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 14996 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0803_
timestamp 1667941163
transform 1 0 28888 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 38088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 34224 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 37444 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 37352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 38088 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 37352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 37536 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0814_
timestamp 1667941163
transform 1 0 12420 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 10396 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 10304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 13524 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 14720 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 14076 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0825_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26680 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 13984 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 28980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 36800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 37444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 24380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 25760 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0844_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29900 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0845_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30728 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 27232 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0847_
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0848_
timestamp 1667941163
transform 1 0 18124 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0849_
timestamp 1667941163
transform 1 0 18216 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0850_
timestamp 1667941163
transform 1 0 32476 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 32384 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 32568 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0854_
timestamp 1667941163
transform 1 0 34868 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 34408 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0856_
timestamp 1667941163
transform 1 0 21712 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0857_
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0858_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34684 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 32292 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 34684 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 32844 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 32936 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0863_
timestamp 1667941163
transform 1 0 30728 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0864_
timestamp 1667941163
transform 1 0 34868 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0865_
timestamp 1667941163
transform 1 0 31096 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0866_
timestamp 1667941163
transform 1 0 24840 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 23184 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 32292 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 32568 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0870_
timestamp 1667941163
transform 1 0 31372 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0871_
timestamp 1667941163
transform 1 0 34868 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0872_
timestamp 1667941163
transform 1 0 32384 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0873_
timestamp 1667941163
transform 1 0 34868 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0874_
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0875_
timestamp 1667941163
transform 1 0 34868 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0878_
timestamp 1667941163
transform 1 0 22816 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0879_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0881_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 23000 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0883_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 19412 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0885_
timestamp 1667941163
transform 1 0 18216 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0887_
timestamp 1667941163
transform 1 0 20976 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0888_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0889_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 19412 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 21804 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0893_
timestamp 1667941163
transform 1 0 20700 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0894_
timestamp 1667941163
transform 1 0 18124 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 24196 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform 1 0 27600 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0897_
timestamp 1667941163
transform 1 0 29440 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 25852 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0899_
timestamp 1667941163
transform 1 0 25208 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0900_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 31464 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 24932 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0903_
timestamp 1667941163
transform 1 0 18124 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 27600 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0906_
timestamp 1667941163
transform 1 0 29716 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 29256 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0908_
timestamp 1667941163
transform 1 0 28704 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0909_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 30176 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 32292 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0912_
timestamp 1667941163
transform 1 0 23368 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 19228 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 29440 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 27600 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 27140 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 26772 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0918_
timestamp 1667941163
transform 1 0 21988 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0919_
timestamp 1667941163
transform 1 0 18308 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 18216 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 32200 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 29808 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 32384 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform 1 0 29900 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform 1 0 34408 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 34868 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 34776 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 34868 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 34868 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0935_
timestamp 1667941163
transform 1 0 18216 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0936_
timestamp 1667941163
transform 1 0 23736 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0937_
timestamp 1667941163
transform 1 0 27968 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 24840 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 22264 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 19688 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0942_
timestamp 1667941163
transform 1 0 24288 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0943_
timestamp 1667941163
transform 1 0 18124 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 17112 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1667941163
transform 1 0 24656 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1667941163
transform 1 0 24840 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 27416 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 31924 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0950_
timestamp 1667941163
transform 1 0 29808 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 30544 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1667941163
transform 1 0 27324 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0953_
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 19136 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform 1 0 20424 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 22264 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 20056 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0958_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0961_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0989_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 35880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1667941163
transform 1 0 27324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 5796 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 32936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0996_
timestamp 1667941163
transform 1 0 20516 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 36708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 10304 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 37444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 8372 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 35972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 37812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1667941163
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 36156 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 25024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 14904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 30912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 33764 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1667941163
transform 1 0 10028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 27876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 4140 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 28980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 38088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1029_
timestamp 1667941163
transform 1 0 28612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 6624 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 37352 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 32384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 37352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 37444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 9292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1667941163
transform 1 0 33396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1667941163
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1044_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28704 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1045__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 33764 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11040 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1047_
timestamp 1667941163
transform 1 0 27232 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 12052 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1049_
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1051_
timestamp 1667941163
transform 1 0 11776 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1052_
timestamp 1667941163
transform 1 0 11960 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1053_
timestamp 1667941163
transform 1 0 31096 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 36156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1055_
timestamp 1667941163
transform 1 0 37536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1055__143
timestamp 1667941163
transform 1 0 37720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1056_
timestamp 1667941163
transform 1 0 34592 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1057_
timestamp 1667941163
transform 1 0 37168 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1058_
timestamp 1667941163
transform 1 0 31372 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1059_
timestamp 1667941163
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 14444 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1061_
timestamp 1667941163
transform 1 0 12512 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1062__144
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1062_
timestamp 1667941163
transform 1 0 12972 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 35604 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 35696 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1065_
timestamp 1667941163
transform 1 0 15364 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 35236 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 15364 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1068__145
timestamp 1667941163
transform 1 0 38088 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 37168 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 32292 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 30636 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1072_
timestamp 1667941163
transform 1 0 12328 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1073_
timestamp 1667941163
transform 1 0 37536 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1073__146
timestamp 1667941163
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1074_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 35972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1077__147
timestamp 1667941163
transform 1 0 33488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 31648 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1080_
timestamp 1667941163
transform 1 0 14260 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1081_
timestamp 1667941163
transform 1 0 37444 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1081__148
timestamp 1667941163
transform 1 0 37536 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 32292 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 37444 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1084_
timestamp 1667941163
transform 1 0 34684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1085__149
timestamp 1667941163
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 10212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 14260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 20332 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1089__150
timestamp 1667941163
transform 1 0 8372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 9844 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1093_
timestamp 1667941163
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1093__151
timestamp 1667941163
transform 1 0 13248 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1094_
timestamp 1667941163
transform 1 0 14904 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1095_
timestamp 1667941163
transform 1 0 14168 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1097__152
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 22724 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1099_
timestamp 1667941163
transform 1 0 21712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 22632 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1101_
timestamp 1667941163
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1102_
timestamp 1667941163
transform 1 0 12144 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1102__153
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1103_
timestamp 1667941163
transform 1 0 22540 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 11960 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1105_
timestamp 1667941163
transform 1 0 14536 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1106_
timestamp 1667941163
transform 1 0 11500 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1107_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1108__154
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1108_
timestamp 1667941163
transform 1 0 9936 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1111_
timestamp 1667941163
transform 1 0 11040 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 9384 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1113_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1114_
timestamp 1667941163
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1114__155
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform 1 0 28520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1117_
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1120__156
timestamp 1667941163
transform 1 0 8280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 8924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 7728 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 9108 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 7544 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1125_
timestamp 1667941163
transform 1 0 15548 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 13984 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 11500 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 11684 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1128__157
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 9936 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 11776 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 15640 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 14444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 25576 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 24932 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1140__158
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 25024 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 14444 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 27324 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 27968 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 26680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 26864 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 15456 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1152__159
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 12788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1153_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1154_
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 23736 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 12420 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1159_
timestamp 1667941163
transform 1 0 37076 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 15456 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 30544 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 10488 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1164__160
timestamp 1667941163
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 32568 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1167_
timestamp 1667941163
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 33856 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 12512 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 20792 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1173_
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1174_
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1175__161
timestamp 1667941163
transform 1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1175_
timestamp 1667941163
transform 1 0 29256 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1176_
timestamp 1667941163
transform 1 0 17112 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1177_
timestamp 1667941163
transform 1 0 2300 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1178_
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1179_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 15916 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1182_
timestamp 1667941163
transform 1 0 15732 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1183_
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 10304 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1185_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1186_
timestamp 1667941163
transform 1 0 16008 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1187__162
timestamp 1667941163
transform 1 0 37536 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1187_
timestamp 1667941163
transform 1 0 36432 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1188_
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1189_
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1190_
timestamp 1667941163
transform 1 0 18216 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1191_
timestamp 1667941163
transform 1 0 33212 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1192_
timestamp 1667941163
transform 1 0 34040 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1193_
timestamp 1667941163
transform 1 0 22724 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1194_
timestamp 1667941163
transform 1 0 36248 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1195_
timestamp 1667941163
transform 1 0 30636 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1196_
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1197_
timestamp 1667941163
transform 1 0 33856 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1198_
timestamp 1667941163
transform 1 0 30176 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1199_
timestamp 1667941163
transform 1 0 35328 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1199__163
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1200_
timestamp 1667941163
transform 1 0 33028 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1201_
timestamp 1667941163
transform 1 0 15180 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1202_
timestamp 1667941163
transform 1 0 10028 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1203_
timestamp 1667941163
transform 1 0 15824 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1204_
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1205_
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1206_
timestamp 1667941163
transform 1 0 30452 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1207_
timestamp 1667941163
transform 1 0 9108 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1208_
timestamp 1667941163
transform 1 0 12144 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1209_
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1210_
timestamp 1667941163
transform 1 0 10672 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1211__164
timestamp 1667941163
transform 1 0 6992 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1211_
timestamp 1667941163
transform 1 0 7636 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1212_
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1213_
timestamp 1667941163
transform 1 0 10396 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 10672 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1215_
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1216_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1217_
timestamp 1667941163
transform 1 0 14168 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1218_
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 13340 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1220_
timestamp 1667941163
transform 1 0 10212 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1667941163
transform 1 0 32016 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1667941163
transform 1 0 16376 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1223__165
timestamp 1667941163
transform 1 0 25392 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1224_
timestamp 1667941163
transform 1 0 22908 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1225_
timestamp 1667941163
transform 1 0 32476 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1226_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1227_
timestamp 1667941163
transform 1 0 16468 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1228_
timestamp 1667941163
transform 1 0 29900 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1229_
timestamp 1667941163
transform 1 0 28980 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1231_
timestamp 1667941163
transform 1 0 31464 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1232_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1233_
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1234_
timestamp 1667941163
transform 1 0 12788 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1235__166
timestamp 1667941163
transform 1 0 14628 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1235_
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1236_
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1237_
timestamp 1667941163
transform 1 0 23276 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1238_
timestamp 1667941163
transform 1 0 16836 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1239_
timestamp 1667941163
transform 1 0 16928 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1240_
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1241_
timestamp 1667941163
transform 1 0 24932 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1242_
timestamp 1667941163
transform 1 0 19044 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1243_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1244_
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26956 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 21988 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 20516 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 25300 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 20516 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 20976 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 26864 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 27140 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 28060 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 33304 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 29716 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 33396 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 32752 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1667941163
transform 1 0 5152 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 35512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform 1 0 25760 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 7636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform 1 0 20332 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 31004 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1667941163
transform 1 0 15456 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 32292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform 1 0 37444 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 26404 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 37444 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 36800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 32108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 16100 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1667941163
transform 1 0 37444 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 3128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 3772 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 36064 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 8372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1667941163
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 5152 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 14720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 18216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 13616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 37996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  sb_1__0__141
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 3 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 4 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 5 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 6 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 7 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 8 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 9 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 10 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 11 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 12 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 13 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 14 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 15 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 16 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 17 nsew signal input
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 18 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 19 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 20 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 21 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 22 nsew signal tristate
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 23 nsew signal tristate
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 24 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 25 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 26 nsew signal tristate
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 27 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 28 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 29 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 30 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 32 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 33 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 34 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 35 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 36 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 38 nsew signal tristate
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 39 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 40 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 41 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 42 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 43 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 44 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 45 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 46 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 47 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 48 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 49 nsew signal input
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 50 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 51 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 52 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 53 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 54 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 55 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 56 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 57 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 58 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 59 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 60 nsew signal tristate
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 61 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 62 nsew signal tristate
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 63 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 64 nsew signal tristate
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 65 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 66 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 67 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 68 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 69 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 70 nsew signal tristate
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 71 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 72 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 73 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 74 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 75 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 76 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 77 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 78 nsew signal input
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 79 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 80 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_in[12]
port 81 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chany_top_in[13]
port 82 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[14]
port 83 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 84 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 85 nsew signal input
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_top_in[17]
port 86 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_top_in[18]
port 87 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_in[1]
port 88 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 89 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_top_in[3]
port 90 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[4]
port 91 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_top_in[5]
port 92 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 93 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 94 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_top_in[8]
port 95 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 96 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_top_out[0]
port 97 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 98 nsew signal tristate
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 99 nsew signal tristate
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 100 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 101 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_out[14]
port 102 nsew signal tristate
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_out[15]
port 103 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_out[16]
port 104 nsew signal tristate
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 105 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_out[18]
port 106 nsew signal tristate
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_out[2]
port 108 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[3]
port 109 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[4]
port 110 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 111 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[6]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[7]
port 113 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_top_out[8]
port 114 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_top_out[9]
port 115 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 116 nsew signal input
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 117 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 118 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 119 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 120 nsew signal input
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 121 nsew signal input
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 122 nsew signal input
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 123 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 124 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 125 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 pReset
port 126 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 prog_clk
port 127 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 131 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 132 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 136 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 137 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 138 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 139 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 140 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 141 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 vssd1
port 143 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 26542 22542 26542 22542 0 _0000_
rlabel metal1 21567 30634 21567 30634 0 _0001_
rlabel via2 14490 32827 14490 32827 0 _0002_
rlabel metal2 22218 25738 22218 25738 0 _0003_
rlabel metal1 12650 35224 12650 35224 0 _0004_
rlabel metal1 14490 34952 14490 34952 0 _0005_
rlabel metal2 13662 31161 13662 31161 0 _0006_
rlabel metal1 13294 30056 13294 30056 0 _0007_
rlabel metal1 17059 27030 17059 27030 0 _0008_
rlabel metal1 14398 27608 14398 27608 0 _0009_
rlabel metal1 31740 20570 31740 20570 0 _0010_
rlabel metal1 31556 21114 31556 21114 0 _0011_
rlabel metal1 28658 18938 28658 18938 0 _0012_
rlabel metal1 28198 20026 28198 20026 0 _0013_
rlabel metal1 26181 26282 26181 26282 0 _0014_
rlabel metal1 35466 20570 35466 20570 0 _0015_
rlabel metal2 12926 28118 12926 28118 0 _0016_
rlabel metal1 14674 18326 14674 18326 0 _0017_
rlabel metal1 14582 25704 14582 25704 0 _0018_
rlabel via2 31142 16541 31142 16541 0 _0019_
rlabel metal1 17250 26792 17250 26792 0 _0020_
rlabel metal1 31149 34646 31149 34646 0 _0021_
rlabel metal1 29946 17850 29946 17850 0 _0022_
rlabel metal1 37076 15130 37076 15130 0 _0023_
rlabel metal1 34132 20978 34132 20978 0 _0024_
rlabel metal1 36156 20570 36156 20570 0 _0025_
rlabel metal2 28198 21828 28198 21828 0 _0026_
rlabel metal1 23000 21658 23000 21658 0 _0027_
rlabel metal2 31004 22080 31004 22080 0 _0028_
rlabel metal2 31280 22916 31280 22916 0 _0029_
rlabel metal2 28612 27132 28612 27132 0 _0030_
rlabel via2 11086 31195 11086 31195 0 _0031_
rlabel metal1 12742 35088 12742 35088 0 _0032_
rlabel metal1 18354 32538 18354 32538 0 _0033_
rlabel metal1 17066 32742 17066 32742 0 _0034_
rlabel via2 12926 34085 12926 34085 0 _0035_
rlabel metal1 34139 36074 34139 36074 0 _0036_
rlabel via2 35006 16405 35006 16405 0 _0037_
rlabel metal1 38042 16490 38042 16490 0 _0038_
rlabel metal1 36248 18122 36248 18122 0 _0039_
rlabel metal1 33120 21386 33120 21386 0 _0040_
rlabel metal1 37950 18938 37950 18938 0 _0041_
rlabel metal1 37674 17850 37674 17850 0 _0042_
rlabel metal1 37260 22202 37260 22202 0 _0043_
rlabel metal1 37720 17714 37720 17714 0 _0044_
rlabel metal1 38502 16422 38502 16422 0 _0045_
rlabel metal1 36853 21590 36853 21590 0 _0046_
rlabel metal1 30820 18938 30820 18938 0 _0047_
rlabel metal2 13202 29954 13202 29954 0 _0048_
rlabel metal1 18485 29206 18485 29206 0 _0049_
rlabel metal1 20746 33048 20746 33048 0 _0050_
rlabel via2 13662 35275 13662 35275 0 _0051_
rlabel metal2 12650 35275 12650 35275 0 _0052_
rlabel metal2 10166 35853 10166 35853 0 _0053_
rlabel metal2 14858 35088 14858 35088 0 _0054_
rlabel metal1 15456 35598 15456 35598 0 _0055_
rlabel metal1 18124 34102 18124 34102 0 _0056_
rlabel metal1 19550 33449 19550 33449 0 _0057_
rlabel metal1 17066 32334 17066 32334 0 _0058_
rlabel metal2 29118 18768 29118 18768 0 _0059_
rlabel metal2 15134 33303 15134 33303 0 _0060_
rlabel metal1 28060 14586 28060 14586 0 _0061_
rlabel metal2 33718 16320 33718 16320 0 _0062_
rlabel metal1 33771 27370 33771 27370 0 _0063_
rlabel metal2 36938 21386 36938 21386 0 _0064_
rlabel metal1 38272 18870 38272 18870 0 _0065_
rlabel metal1 29401 27370 29401 27370 0 _0066_
rlabel metal2 30958 15657 30958 15657 0 _0067_
rlabel metal1 24472 21658 24472 21658 0 _0068_
rlabel metal1 25484 21114 25484 21114 0 _0069_
rlabel metal1 24840 20570 24840 20570 0 _0070_
rlabel metal1 24886 21590 24886 21590 0 _0071_
rlabel metal1 21029 22678 21029 22678 0 _0072_
rlabel metal1 18446 23623 18446 23623 0 _0073_
rlabel metal1 21114 26391 21114 26391 0 _0074_
rlabel via2 27278 17323 27278 17323 0 _0075_
rlabel metal1 34362 15130 34362 15130 0 _0076_
rlabel metal1 35558 16218 35558 16218 0 _0077_
rlabel metal1 30452 17782 30452 17782 0 _0078_
rlabel metal1 15042 31960 15042 31960 0 _0079_
rlabel metal1 16100 33558 16100 33558 0 _0080_
rlabel metal1 14306 31926 14306 31926 0 _0081_
rlabel via2 33718 12699 33718 12699 0 _0082_
rlabel metal1 38272 13498 38272 13498 0 _0083_
rlabel metal1 35282 20230 35282 20230 0 _0084_
rlabel metal2 36846 34850 36846 34850 0 _0085_
rlabel metal2 36846 36312 36846 36312 0 _0086_
rlabel metal1 35696 35802 35696 35802 0 _0087_
rlabel metal2 20654 36057 20654 36057 0 _0088_
rlabel metal1 29854 36822 29854 36822 0 _0089_
rlabel via2 32890 13515 32890 13515 0 _0090_
rlabel via3 33741 24956 33741 24956 0 _0091_
rlabel metal1 36892 12410 36892 12410 0 _0092_
rlabel via2 37582 11883 37582 11883 0 _0093_
rlabel metal1 34868 35462 34868 35462 0 _0094_
rlabel metal2 31694 34680 31694 34680 0 _0095_
rlabel metal2 37582 25602 37582 25602 0 _0096_
rlabel metal1 32844 18326 32844 18326 0 _0097_
rlabel metal1 27508 18394 27508 18394 0 _0098_
rlabel metal2 26542 15215 26542 15215 0 _0099_
rlabel metal1 38180 15130 38180 15130 0 _0100_
rlabel metal1 38870 14586 38870 14586 0 _0101_
rlabel via2 36478 16235 36478 16235 0 _0102_
rlabel metal1 38134 13974 38134 13974 0 _0103_
rlabel metal2 36754 10387 36754 10387 0 _0104_
rlabel metal1 37497 32810 37497 32810 0 _0105_
rlabel metal1 26496 21114 26496 21114 0 _0106_
rlabel via3 36317 31756 36317 31756 0 _0107_
rlabel metal1 23138 20026 23138 20026 0 _0108_
rlabel metal1 20884 26010 20884 26010 0 _0109_
rlabel metal2 26128 20502 26128 20502 0 _0110_
rlabel metal1 30498 18632 30498 18632 0 _0111_
rlabel metal1 27600 19414 27600 19414 0 _0112_
rlabel metal1 26082 20026 26082 20026 0 _0113_
rlabel metal2 23874 24888 23874 24888 0 _0114_
rlabel metal1 23736 20026 23736 20026 0 _0115_
rlabel metal2 15502 35292 15502 35292 0 _0116_
rlabel metal2 19504 28084 19504 28084 0 _0117_
rlabel metal1 26542 20910 26542 20910 0 _0118_
rlabel via2 19826 30277 19826 30277 0 _0119_
rlabel metal2 14398 18428 14398 18428 0 _0120_
rlabel metal2 17250 21726 17250 21726 0 _0121_
rlabel metal1 34178 35190 34178 35190 0 _0122_
rlabel metal1 34270 18224 34270 18224 0 _0123_
rlabel metal1 13708 35054 13708 35054 0 _0124_
rlabel metal2 14030 32708 14030 32708 0 _0125_
rlabel metal1 8510 31824 8510 31824 0 _0126_
rlabel metal2 8694 25092 8694 25092 0 _0127_
rlabel metal1 7498 20502 7498 20502 0 _0128_
rlabel metal2 22310 16796 22310 16796 0 _0129_
rlabel metal2 26450 13124 26450 13124 0 _0130_
rlabel metal2 21022 10812 21022 10812 0 _0131_
rlabel metal1 6210 35054 6210 35054 0 _0132_
rlabel metal1 9154 31450 9154 31450 0 _0133_
rlabel metal2 9246 27268 9246 27268 0 _0134_
rlabel metal2 19826 15878 19826 15878 0 _0135_
rlabel metal2 13018 16218 13018 16218 0 _0136_
rlabel metal1 12650 12172 12650 12172 0 _0137_
rlabel metal1 22908 12614 22908 12614 0 _0138_
rlabel metal1 20654 8908 20654 8908 0 _0139_
rlabel metal1 15824 22202 15824 22202 0 _0140_
rlabel metal1 15226 13940 15226 13940 0 _0141_
rlabel metal2 11270 17476 11270 17476 0 _0142_
rlabel metal2 7774 25670 7774 25670 0 _0143_
rlabel metal2 19642 13498 19642 13498 0 _0144_
rlabel metal1 11638 15130 11638 15130 0 _0145_
rlabel metal1 34270 34612 34270 34612 0 _0146_
rlabel metal2 37674 29002 37674 29002 0 _0147_
rlabel metal2 13570 26758 13570 26758 0 _0148_
rlabel metal2 31418 15164 31418 15164 0 _0149_
rlabel metal2 36110 10948 36110 10948 0 _0150_
rlabel metal2 34362 11322 34362 11322 0 _0151_
rlabel metal2 19274 19839 19274 19839 0 _0152_
rlabel metal2 27462 17952 27462 17952 0 _0153_
rlabel metal1 36754 34612 36754 34612 0 _0154_
rlabel metal1 36754 36720 36754 36720 0 _0155_
rlabel metal1 38962 14994 38962 14994 0 _0156_
rlabel metal2 28934 21080 28934 21080 0 _0157_
rlabel metal1 34086 13498 34086 13498 0 _0158_
rlabel metal2 11270 29818 11270 29818 0 _0159_
rlabel metal1 25806 19414 25806 19414 0 _0160_
rlabel metal1 9614 33524 9614 33524 0 _0161_
rlabel metal1 15272 31994 15272 31994 0 _0162_
rlabel metal1 22816 21114 22816 21114 0 _0163_
rlabel metal2 12006 33048 12006 33048 0 _0164_
rlabel metal1 11822 31722 11822 31722 0 _0165_
rlabel metal2 32430 33728 32430 33728 0 _0166_
rlabel metal2 36386 11254 36386 11254 0 _0167_
rlabel metal1 36938 11050 36938 11050 0 _0168_
rlabel metal1 34914 18394 34914 18394 0 _0169_
rlabel metal1 37260 12138 37260 12138 0 _0170_
rlabel metal1 31556 33626 31556 33626 0 _0171_
rlabel metal1 37030 10778 37030 10778 0 _0172_
rlabel metal1 13616 34170 13616 34170 0 _0173_
rlabel metal1 12880 32198 12880 32198 0 _0174_
rlabel metal1 13432 29274 13432 29274 0 _0175_
rlabel metal1 35190 12954 35190 12954 0 _0176_
rlabel metal1 35788 12954 35788 12954 0 _0177_
rlabel metal2 15594 28050 15594 28050 0 _0178_
rlabel metal2 36294 18530 36294 18530 0 _0179_
rlabel metal1 16836 30294 16836 30294 0 _0180_
rlabel metal1 37168 17850 37168 17850 0 _0181_
rlabel metal2 14030 23358 14030 23358 0 _0182_
rlabel metal1 33856 15674 33856 15674 0 _0183_
rlabel metal2 30866 20638 30866 20638 0 _0184_
rlabel metal1 12650 16150 12650 16150 0 _0185_
rlabel metal1 34454 11322 34454 11322 0 _0186_
rlabel metal1 35972 10778 35972 10778 0 _0187_
rlabel metal1 34776 11866 34776 11866 0 _0188_
rlabel metal1 35236 14450 35236 14450 0 _0189_
rlabel metal2 31878 14620 31878 14620 0 _0190_
rlabel metal1 13938 27098 13938 27098 0 _0191_
rlabel metal2 31326 16286 31326 16286 0 _0192_
rlabel metal1 13708 28730 13708 28730 0 _0193_
rlabel metal1 37536 28730 37536 28730 0 _0194_
rlabel metal1 33304 34510 33304 34510 0 _0195_
rlabel metal1 37260 32402 37260 32402 0 _0196_
rlabel metal1 34546 34170 34546 34170 0 _0197_
rlabel metal1 10442 15572 10442 15572 0 _0198_
rlabel metal2 19458 13668 19458 13668 0 _0199_
rlabel metal2 14398 14756 14398 14756 0 _0200_
rlabel metal1 20700 14994 20700 14994 0 _0201_
rlabel metal1 8832 26010 8832 26010 0 _0202_
rlabel metal1 10074 17544 10074 17544 0 _0203_
rlabel metal1 8924 25330 8924 25330 0 _0204_
rlabel metal2 17066 16286 17066 16286 0 _0205_
rlabel metal1 13800 13974 13800 13974 0 _0206_
rlabel metal1 15364 23290 15364 23290 0 _0207_
rlabel metal2 14398 15912 14398 15912 0 _0208_
rlabel metal2 27370 18462 27370 18462 0 _0209_
rlabel metal2 20470 9316 20470 9316 0 _0210_
rlabel metal2 22862 11492 22862 11492 0 _0211_
rlabel metal2 22126 9826 22126 9826 0 _0212_
rlabel metal1 22908 12274 22908 12274 0 _0213_
rlabel metal2 13294 15198 13294 15198 0 _0214_
rlabel metal1 12420 12750 12420 12750 0 _0215_
rlabel metal1 22724 16150 22724 16150 0 _0216_
rlabel metal2 12190 18088 12190 18088 0 _0217_
rlabel metal2 15042 13124 15042 13124 0 _0218_
rlabel metal1 11730 21896 11730 21896 0 _0219_
rlabel metal1 11408 32470 11408 32470 0 _0220_
rlabel metal2 9706 28594 9706 28594 0 _0221_
rlabel metal1 9338 35156 9338 35156 0 _0222_
rlabel metal2 8510 34408 8510 34408 0 _0223_
rlabel metal2 13018 28764 13018 28764 0 _0224_
rlabel metal1 9016 34578 9016 34578 0 _0225_
rlabel metal1 27094 13498 27094 13498 0 _0226_
rlabel metal1 20884 10778 20884 10778 0 _0227_
rlabel metal1 23506 17068 23506 17068 0 _0228_
rlabel metal1 28888 13906 28888 13906 0 _0229_
rlabel metal1 20608 13362 20608 13362 0 _0230_
rlabel metal1 29026 15538 29026 15538 0 _0231_
rlabel metal2 9338 24412 9338 24412 0 _0232_
rlabel metal1 8234 22610 8234 22610 0 _0233_
rlabel metal2 8326 31212 8326 31212 0 _0234_
rlabel metal1 7774 28186 7774 28186 0 _0235_
rlabel metal1 9292 22202 9292 22202 0 _0236_
rlabel metal1 7360 28118 7360 28118 0 _0237_
rlabel metal1 15640 32470 15640 32470 0 _0238_
rlabel metal1 14306 28730 14306 28730 0 _0239_
rlabel metal1 11776 24378 11776 24378 0 _0240_
rlabel metal2 12466 23528 12466 23528 0 _0241_
rlabel metal1 10626 21590 10626 21590 0 _0242_
rlabel metal2 12006 28696 12006 28696 0 _0243_
rlabel metal1 21758 19822 21758 19822 0 _0244_
rlabel metal2 23690 20706 23690 20706 0 _0245_
rlabel metal1 15364 29818 15364 29818 0 _0246_
rlabel metal2 13938 25534 13938 25534 0 _0247_
rlabel metal1 11178 33558 11178 33558 0 _0248_
rlabel metal2 14674 25262 14674 25262 0 _0249_
rlabel metal1 26082 13974 26082 13974 0 _0250_
rlabel metal2 25162 15640 25162 15640 0 _0251_
rlabel metal2 19642 11322 19642 11322 0 _0252_
rlabel metal2 24794 10200 24794 10200 0 _0253_
rlabel metal2 17066 10880 17066 10880 0 _0254_
rlabel metal1 25806 11798 25806 11798 0 _0255_
rlabel metal1 15364 18394 15364 18394 0 _0256_
rlabel metal1 27048 16762 27048 16762 0 _0257_
rlabel metal1 28612 16218 28612 16218 0 _0258_
rlabel metal1 27232 13158 27232 13158 0 _0259_
rlabel metal1 26680 13430 26680 13430 0 _0260_
rlabel metal1 19366 18938 19366 18938 0 _0261_
rlabel metal2 17066 35870 17066 35870 0 _0262_
rlabel metal1 16100 34170 16100 34170 0 _0263_
rlabel metal1 8832 36278 8832 36278 0 _0264_
rlabel metal2 10626 35955 10626 35955 0 _0265_
rlabel metal1 33120 32538 33120 32538 0 _0266_
rlabel metal1 15686 33626 15686 33626 0 _0267_
rlabel metal1 21298 21114 21298 21114 0 _0268_
rlabel metal2 21390 21046 21390 21046 0 _0269_
rlabel metal1 17388 32946 17388 32946 0 _0270_
rlabel metal2 11178 36210 11178 36210 0 _0271_
rlabel metal2 37030 25840 37030 25840 0 _0272_
rlabel metal1 14582 27914 14582 27914 0 _0273_
rlabel metal2 29578 20706 29578 20706 0 _0274_
rlabel metal2 20746 19550 20746 19550 0 _0275_
rlabel metal2 11086 18258 11086 18258 0 _0276_
rlabel metal1 19366 17510 19366 17510 0 _0277_
rlabel metal1 32798 15368 32798 15368 0 _0278_
rlabel metal1 29532 16762 29532 16762 0 _0279_
rlabel metal2 32522 15742 32522 15742 0 _0280_
rlabel metal1 34638 16150 34638 16150 0 _0281_
rlabel metal1 35144 19754 35144 19754 0 _0282_
rlabel metal1 14306 24310 14306 24310 0 _0283_
rlabel metal2 21390 17442 21390 17442 0 _0284_
rlabel metal2 19642 19992 19642 19992 0 _0285_
rlabel metal1 29486 19414 29486 19414 0 _0286_
rlabel metal1 22586 16762 22586 16762 0 _0287_
rlabel metal1 29578 16218 29578 16218 0 _0288_
rlabel metal1 16652 22406 16652 22406 0 _0289_
rlabel metal1 4692 33626 4692 33626 0 _0290_
rlabel metal1 2116 34714 2116 34714 0 _0291_
rlabel metal1 11500 29206 11500 29206 0 _0292_
rlabel metal1 11362 25942 11362 25942 0 _0293_
rlabel metal1 15594 32538 15594 32538 0 _0294_
rlabel metal1 15870 24786 15870 24786 0 _0295_
rlabel metal1 1794 36856 1794 36856 0 _0296_
rlabel metal2 12742 25704 12742 25704 0 _0297_
rlabel metal2 32522 19754 32522 19754 0 _0298_
rlabel metal1 16606 28594 16606 28594 0 _0299_
rlabel metal1 36340 31790 36340 31790 0 _0300_
rlabel metal1 28704 11050 28704 11050 0 _0301_
rlabel metal1 15824 25466 15824 25466 0 _0302_
rlabel metal1 19274 12886 19274 12886 0 _0303_
rlabel metal2 33442 14552 33442 14552 0 _0304_
rlabel metal1 34914 15674 34914 15674 0 _0305_
rlabel metal1 22540 15062 22540 15062 0 _0306_
rlabel metal1 36156 19890 36156 19890 0 _0307_
rlabel metal2 30866 14382 30866 14382 0 _0308_
rlabel metal1 25990 18632 25990 18632 0 _0309_
rlabel metal2 35650 19448 35650 19448 0 _0310_
rlabel metal1 30452 14246 30452 14246 0 _0311_
rlabel metal1 35282 13498 35282 13498 0 _0312_
rlabel metal2 33258 17816 33258 17816 0 _0313_
rlabel metal1 15226 28730 15226 28730 0 _0314_
rlabel metal1 12282 17238 12282 17238 0 _0315_
rlabel metal2 16974 16643 16974 16643 0 _0316_
rlabel metal1 11776 22950 11776 22950 0 _0317_
rlabel metal2 25622 16728 25622 16728 0 _0318_
rlabel metal1 31142 18394 31142 18394 0 _0319_
rlabel metal1 9706 30634 9706 30634 0 _0320_
rlabel metal2 12374 26622 12374 26622 0 _0321_
rlabel metal1 14720 34578 14720 34578 0 _0322_
rlabel metal1 10442 35530 10442 35530 0 _0323_
rlabel metal2 8602 34680 8602 34680 0 _0324_
rlabel metal1 13938 33592 13938 33592 0 _0325_
rlabel metal2 10350 35496 10350 35496 0 _0326_
rlabel metal2 10902 31144 10902 31144 0 _0327_
rlabel metal2 9890 32878 9890 32878 0 _0328_
rlabel metal1 11500 28118 11500 28118 0 _0329_
rlabel metal1 13110 31382 13110 31382 0 _0330_
rlabel metal1 15364 36822 15364 36822 0 _0331_
rlabel metal1 13018 34578 13018 34578 0 _0332_
rlabel metal2 10442 26792 10442 26792 0 _0333_
rlabel metal1 32338 18394 32338 18394 0 _0334_
rlabel metal1 16882 33626 16882 33626 0 _0335_
rlabel metal1 24242 31926 24242 31926 0 _0336_
rlabel metal2 20746 17034 20746 17034 0 _0337_
rlabel metal1 32154 17238 32154 17238 0 _0338_
rlabel metal2 27370 15198 27370 15198 0 _0339_
rlabel metal2 17526 18530 17526 18530 0 _0340_
rlabel metal2 30498 17442 30498 17442 0 _0341_
rlabel metal2 29210 15470 29210 15470 0 _0342_
rlabel metal2 29946 20876 29946 20876 0 _0343_
rlabel metal1 31694 17544 31694 17544 0 _0344_
rlabel metal1 18400 18938 18400 18938 0 _0345_
rlabel metal2 20194 17816 20194 17816 0 _0346_
rlabel metal1 13386 10710 13386 10710 0 _0347_
rlabel metal1 14950 19754 14950 19754 0 _0348_
rlabel metal1 17756 13974 17756 13974 0 _0349_
rlabel metal2 23414 14739 23414 14739 0 _0350_
rlabel metal1 18308 11866 18308 11866 0 _0351_
rlabel metal2 17158 14552 17158 14552 0 _0352_
rlabel metal1 15870 17306 15870 17306 0 _0353_
rlabel metal1 23736 14042 23736 14042 0 _0354_
rlabel metal1 19918 19414 19918 19414 0 _0355_
rlabel metal1 15364 21658 15364 21658 0 _0356_
rlabel metal1 13616 22746 13616 22746 0 _0357_
rlabel metal3 1142 19108 1142 19108 0 ccff_head
rlabel metal3 1234 7548 1234 7548 0 ccff_tail
rlabel metal2 5198 38260 5198 38260 0 chanx_left_in[0]
rlabel metal3 1142 5508 1142 5508 0 chanx_left_in[10]
rlabel metal2 35466 1860 35466 1860 0 chanx_left_in[11]
rlabel metal2 25806 1588 25806 1588 0 chanx_left_in[12]
rlabel metal3 1188 22508 1188 22508 0 chanx_left_in[13]
rlabel metal3 1142 6868 1142 6868 0 chanx_left_in[14]
rlabel metal1 17388 36754 17388 36754 0 chanx_left_in[15]
rlabel metal3 1142 38828 1142 38828 0 chanx_left_in[16]
rlabel metal2 12926 1588 12926 1588 0 chanx_left_in[17]
rlabel metal2 29026 1588 29026 1588 0 chanx_left_in[18]
rlabel metal1 27692 37230 27692 37230 0 chanx_left_in[1]
rlabel metal1 6210 37298 6210 37298 0 chanx_left_in[2]
rlabel metal2 24518 1588 24518 1588 0 chanx_left_in[3]
rlabel metal1 7866 36788 7866 36788 0 chanx_left_in[4]
rlabel metal2 20010 1588 20010 1588 0 chanx_left_in[5]
rlabel metal3 1142 17068 1142 17068 0 chanx_left_in[6]
rlabel metal3 1924 2108 1924 2108 0 chanx_left_in[7]
rlabel metal1 28750 37196 28750 37196 0 chanx_left_in[8]
rlabel metal2 11638 1588 11638 1588 0 chanx_left_in[9]
rlabel metal2 38226 32385 38226 32385 0 chanx_left_out[0]
rlabel via2 38226 27285 38226 27285 0 chanx_left_out[10]
rlabel metal2 9706 1520 9706 1520 0 chanx_left_out[11]
rlabel metal3 1050 748 1050 748 0 chanx_left_out[12]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[13]
rlabel metal1 14904 37094 14904 37094 0 chanx_left_out[14]
rlabel metal2 38226 30515 38226 30515 0 chanx_left_out[15]
rlabel metal2 38226 28815 38226 28815 0 chanx_left_out[16]
rlabel metal1 32430 36890 32430 36890 0 chanx_left_out[17]
rlabel metal2 18078 1520 18078 1520 0 chanx_left_out[18]
rlabel metal1 36248 37094 36248 37094 0 chanx_left_out[1]
rlabel metal3 38740 12308 38740 12308 0 chanx_left_out[2]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[3]
rlabel metal3 1234 30668 1234 30668 0 chanx_left_out[4]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[5]
rlabel metal2 36846 2193 36846 2193 0 chanx_left_out[6]
rlabel metal2 20010 38158 20010 38158 0 chanx_left_out[7]
rlabel via2 38226 35445 38226 35445 0 chanx_left_out[8]
rlabel metal1 36662 2550 36662 2550 0 chanx_left_out[9]
rlabel metal2 20378 37196 20378 37196 0 chanx_right_in[0]
rlabel metal2 34178 1554 34178 1554 0 chanx_right_in[10]
rlabel metal1 31096 35666 31096 35666 0 chanx_right_in[11]
rlabel metal1 34776 37230 34776 37230 0 chanx_right_in[12]
rlabel metal1 37306 36142 37306 36142 0 chanx_right_in[13]
rlabel metal1 15824 37298 15824 37298 0 chanx_right_in[14]
rlabel metal2 38318 9707 38318 9707 0 chanx_right_in[15]
rlabel metal2 32522 13107 32522 13107 0 chanx_right_in[16]
rlabel metal2 37490 19193 37490 19193 0 chanx_right_in[17]
rlabel metal2 27738 1588 27738 1588 0 chanx_right_in[18]
rlabel metal2 37490 38063 37490 38063 0 chanx_right_in[1]
rlabel metal2 38134 33099 38134 33099 0 chanx_right_in[2]
rlabel metal1 26634 36720 26634 36720 0 chanx_right_in[3]
rlabel metal1 12328 37298 12328 37298 0 chanx_right_in[4]
rlabel metal2 37490 24021 37490 24021 0 chanx_right_in[5]
rlabel metal1 6026 36720 6026 36720 0 chanx_right_in[6]
rlabel metal1 9890 37196 9890 37196 0 chanx_right_in[7]
rlabel metal1 22678 37230 22678 37230 0 chanx_right_in[8]
rlabel metal2 10350 1588 10350 1588 0 chanx_right_in[9]
rlabel metal2 2622 38209 2622 38209 0 chanx_right_out[0]
rlabel metal2 38226 15181 38226 15181 0 chanx_right_out[10]
rlabel metal1 4048 37094 4048 37094 0 chanx_right_out[11]
rlabel metal2 38226 2329 38226 2329 0 chanx_right_out[12]
rlabel metal3 1234 14348 1234 14348 0 chanx_right_out[13]
rlabel metal2 38226 7633 38226 7633 0 chanx_right_out[14]
rlabel metal3 1234 28628 1234 28628 0 chanx_right_out[15]
rlabel metal2 16790 1520 16790 1520 0 chanx_right_out[16]
rlabel metal3 1234 21148 1234 21148 0 chanx_right_out[17]
rlabel metal2 16146 1520 16146 1520 0 chanx_right_out[18]
rlabel metal3 1234 24548 1234 24548 0 chanx_right_out[1]
rlabel metal1 33074 36890 33074 36890 0 chanx_right_out[2]
rlabel metal3 1234 32708 1234 32708 0 chanx_right_out[3]
rlabel metal2 30314 1520 30314 1520 0 chanx_right_out[4]
rlabel metal2 38226 25177 38226 25177 0 chanx_right_out[5]
rlabel via2 38226 5525 38226 5525 0 chanx_right_out[6]
rlabel metal1 27370 37128 27370 37128 0 chanx_right_out[7]
rlabel metal1 38778 35258 38778 35258 0 chanx_right_out[8]
rlabel metal1 37536 36890 37536 36890 0 chanx_right_out[9]
rlabel metal2 690 2438 690 2438 0 chany_top_in[0]
rlabel metal2 5198 1588 5198 1588 0 chany_top_in[10]
rlabel metal2 38686 2098 38686 2098 0 chany_top_in[11]
rlabel metal3 1234 13668 1234 13668 0 chany_top_in[12]
rlabel metal2 38318 21913 38318 21913 0 chany_top_in[13]
rlabel metal1 32338 13328 32338 13328 0 chany_top_in[14]
rlabel metal1 16560 35666 16560 35666 0 chany_top_in[15]
rlabel metal2 3266 1588 3266 1588 0 chany_top_in[16]
rlabel via2 37490 3485 37490 3485 0 chany_top_in[17]
rlabel metal1 37628 11526 37628 11526 0 chany_top_in[18]
rlabel metal3 1234 27268 1234 27268 0 chany_top_in[1]
rlabel metal2 2346 38029 2346 38029 0 chany_top_in[2]
rlabel metal3 1234 25908 1234 25908 0 chany_top_in[3]
rlabel metal3 1234 20468 1234 20468 0 chany_top_in[4]
rlabel metal2 3450 38131 3450 38131 0 chany_top_in[5]
rlabel metal1 37490 34510 37490 34510 0 chany_top_in[6]
rlabel metal2 8418 1588 8418 1588 0 chany_top_in[7]
rlabel metal3 1234 17748 1234 17748 0 chany_top_in[8]
rlabel metal2 23230 1588 23230 1588 0 chany_top_in[9]
rlabel metal2 37398 1792 37398 1792 0 chany_top_out[0]
rlabel metal1 13708 36890 13708 36890 0 chany_top_out[10]
rlabel metal2 30958 1520 30958 1520 0 chany_top_out[11]
rlabel metal2 3910 1792 3910 1792 0 chany_top_out[12]
rlabel metal2 14858 1520 14858 1520 0 chany_top_out[13]
rlabel metal2 38226 29393 38226 29393 0 chany_top_out[15]
rlabel metal2 38226 20519 38226 20519 0 chany_top_out[16]
rlabel metal2 32246 1520 32246 1520 0 chany_top_out[17]
rlabel metal3 1234 23868 1234 23868 0 chany_top_out[18]
rlabel metal2 38226 10353 38226 10353 0 chany_top_out[1]
rlabel metal3 1234 32028 1234 32028 0 chany_top_out[2]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[3]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[4]
rlabel metal2 36754 823 36754 823 0 chany_top_out[5]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[6]
rlabel metal3 1234 12308 1234 12308 0 chany_top_out[7]
rlabel metal3 1234 34068 1234 34068 0 chany_top_out[8]
rlabel metal3 1234 3468 1234 3468 0 chany_top_out[9]
rlabel metal1 33396 28118 33396 28118 0 clknet_0_prog_clk
rlabel metal2 19366 25568 19366 25568 0 clknet_4_0_0_prog_clk
rlabel metal1 32476 22066 32476 22066 0 clknet_4_10_0_prog_clk
rlabel metal1 34868 27506 34868 27506 0 clknet_4_11_0_prog_clk
rlabel metal2 29946 29920 29946 29920 0 clknet_4_12_0_prog_clk
rlabel metal2 30590 33966 30590 33966 0 clknet_4_13_0_prog_clk
rlabel metal1 32476 29138 32476 29138 0 clknet_4_14_0_prog_clk
rlabel metal1 32338 37230 32338 37230 0 clknet_4_15_0_prog_clk
rlabel metal1 18216 27982 18216 27982 0 clknet_4_1_0_prog_clk
rlabel metal1 25024 23086 25024 23086 0 clknet_4_2_0_prog_clk
rlabel metal1 22034 27030 22034 27030 0 clknet_4_3_0_prog_clk
rlabel metal1 18308 32334 18308 32334 0 clknet_4_4_0_prog_clk
rlabel metal2 22034 34238 22034 34238 0 clknet_4_5_0_prog_clk
rlabel metal2 24610 31926 24610 31926 0 clknet_4_6_0_prog_clk
rlabel metal2 26634 34510 26634 34510 0 clknet_4_7_0_prog_clk
rlabel metal1 27416 23698 27416 23698 0 clknet_4_8_0_prog_clk
rlabel metal1 24656 27438 24656 27438 0 clknet_4_9_0_prog_clk
rlabel metal2 46 2098 46 2098 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1234 4148 1234 4148 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 2898 36261 2898 36261 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 9200 37230 9200 37230 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 23414 37230 23414 37230 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal3 1234 29308 1234 29308 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 6486 1588 6486 1588 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 1978 1588 1978 1588 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 1234 8908 1234 8908 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 21298 38226 21298 38226 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal1 26634 18258 26634 18258 0 mem_left_track_1.DFFR_0_.D
rlabel metal1 17933 30906 17933 30906 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 9522 34000 9522 34000 0 mem_left_track_1.DFFR_1_.Q
rlabel via2 19918 33371 19918 33371 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 18814 35241 18814 35241 0 mem_left_track_1.DFFR_3_.Q
rlabel metal2 21206 36805 21206 36805 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 16054 34476 16054 34476 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 13018 34952 13018 34952 0 mem_left_track_1.DFFR_6_.Q
rlabel metal1 19734 33558 19734 33558 0 mem_left_track_1.DFFR_7_.Q
rlabel metal1 21666 34102 21666 34102 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 18354 18564 18354 18564 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 19458 17850 19458 17850 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 30406 16592 30406 16592 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 30222 16286 30222 16286 0 mem_left_track_17.DFFR_3_.Q
rlabel metal1 32062 27540 32062 27540 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 31832 18258 31832 18258 0 mem_left_track_17.DFFR_5_.Q
rlabel metal2 20010 33728 20010 33728 0 mem_left_track_17.DFFR_6_.Q
rlabel metal1 25760 32946 25760 32946 0 mem_left_track_17.DFFR_7_.Q
rlabel metal1 14996 21522 14996 21522 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 18124 15470 18124 15470 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 17710 17170 17710 17170 0 mem_left_track_25.DFFR_2_.Q
rlabel metal1 20056 11730 20056 11730 0 mem_left_track_25.DFFR_3_.Q
rlabel metal1 20884 19346 20884 19346 0 mem_left_track_25.DFFR_4_.Q
rlabel metal1 20470 17170 20470 17170 0 mem_left_track_25.DFFR_5_.Q
rlabel metal1 19182 17714 19182 17714 0 mem_left_track_25.DFFR_6_.Q
rlabel metal1 19504 23766 19504 23766 0 mem_left_track_25.DFFR_7_.Q
rlabel metal1 21160 17170 21160 17170 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 17710 17442 17710 17442 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 20102 17714 20102 17714 0 mem_left_track_33.DFFR_2_.Q
rlabel metal1 32890 20910 32890 20910 0 mem_left_track_33.DFFR_3_.Q
rlabel metal1 29302 20434 29302 20434 0 mem_left_track_33.DFFR_4_.Q
rlabel metal1 13386 27982 13386 27982 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 32246 32402 32246 32402 0 mem_left_track_9.DFFR_1_.Q
rlabel metal3 21367 20604 21367 20604 0 mem_left_track_9.DFFR_2_.Q
rlabel metal2 18446 34782 18446 34782 0 mem_left_track_9.DFFR_3_.Q
rlabel metal2 18262 36346 18262 36346 0 mem_left_track_9.DFFR_4_.Q
rlabel metal2 24840 31756 24840 31756 0 mem_right_track_0.DFFR_0_.D
rlabel metal1 18814 26894 18814 26894 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 18630 22950 18630 22950 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 12972 28492 12972 28492 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 14766 29648 14766 29648 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 19596 32810 19596 32810 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 21298 33082 21298 33082 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 32706 23001 32706 23001 0 mem_right_track_16.DFFR_0_.D
rlabel metal1 33672 22066 33672 22066 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 33718 14994 33718 14994 0 mem_right_track_16.DFFR_1_.Q
rlabel metal3 35351 15572 35351 15572 0 mem_right_track_16.DFFR_2_.Q
rlabel metal1 22034 15062 22034 15062 0 mem_right_track_16.DFFR_3_.Q
rlabel metal1 34684 20910 34684 20910 0 mem_right_track_16.DFFR_4_.Q
rlabel metal1 32384 20434 32384 20434 0 mem_right_track_16.DFFR_5_.Q
rlabel metal1 32522 36040 32522 36040 0 mem_right_track_16.DFFR_6_.Q
rlabel metal1 35995 35054 35995 35054 0 mem_right_track_16.DFFR_7_.Q
rlabel metal1 12650 32232 12650 32232 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 19918 16626 19918 16626 0 mem_right_track_24.DFFR_1_.Q
rlabel metal2 20010 28730 20010 28730 0 mem_right_track_24.DFFR_2_.Q
rlabel metal1 18170 17000 18170 17000 0 mem_right_track_24.DFFR_3_.Q
rlabel metal2 31418 19856 31418 19856 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 36662 19822 36662 19822 0 mem_right_track_24.DFFR_5_.Q
rlabel metal1 35282 22542 35282 22542 0 mem_right_track_24.DFFR_6_.Q
rlabel metal1 35374 13294 35374 13294 0 mem_right_track_24.DFFR_7_.Q
rlabel metal1 33534 23222 33534 23222 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 18814 11662 18814 11662 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 26266 11186 26266 11186 0 mem_right_track_32.DFFR_2_.Q
rlabel metal1 28842 16082 28842 16082 0 mem_right_track_32.DFFR_3_.Q
rlabel metal1 28428 23630 28428 23630 0 mem_right_track_32.DFFR_4_.Q
rlabel metal2 12834 30872 12834 30872 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 15226 28220 15226 28220 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 8326 32963 8326 32963 0 mem_right_track_8.DFFR_2_.Q
rlabel metal2 14950 32708 14950 32708 0 mem_right_track_8.DFFR_3_.Q
rlabel metal2 20654 29546 20654 29546 0 mem_right_track_8.DFFR_4_.Q
rlabel metal1 29762 19346 29762 19346 0 mem_right_track_8.DFFR_5_.Q
rlabel via1 29394 26894 29394 26894 0 mem_right_track_8.DFFR_6_.Q
rlabel metal1 18492 35734 18492 35734 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 19504 32538 19504 32538 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 20378 31858 20378 31858 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 22172 20910 22172 20910 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 29026 20502 29026 20502 0 mem_top_track_0.DFFR_4_.Q
rlabel metal2 34730 36210 34730 36210 0 mem_top_track_0.DFFR_5_.Q
rlabel metal1 34224 11730 34224 11730 0 mem_top_track_10.DFFR_0_.D
rlabel metal1 32798 28424 32798 28424 0 mem_top_track_10.DFFR_0_.Q
rlabel metal1 34178 32810 34178 32810 0 mem_top_track_10.DFFR_1_.Q
rlabel metal1 33396 37298 33396 37298 0 mem_top_track_12.DFFR_0_.Q
rlabel metal2 34178 36487 34178 36487 0 mem_top_track_12.DFFR_1_.Q
rlabel metal1 36708 32334 36708 32334 0 mem_top_track_14.DFFR_0_.Q
rlabel metal2 11914 14722 11914 14722 0 mem_top_track_14.DFFR_1_.Q
rlabel metal1 17434 16592 17434 16592 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 8418 25228 8418 25228 0 mem_top_track_16.DFFR_1_.Q
rlabel metal1 11178 21998 11178 21998 0 mem_top_track_18.DFFR_0_.Q
rlabel metal1 11822 18802 11822 18802 0 mem_top_track_18.DFFR_1_.Q
rlabel metal2 35926 36057 35926 36057 0 mem_top_track_2.DFFR_0_.Q
rlabel metal1 36340 36006 36340 36006 0 mem_top_track_2.DFFR_1_.Q
rlabel metal1 32568 19210 32568 19210 0 mem_top_track_2.DFFR_2_.Q
rlabel metal1 37536 10710 37536 10710 0 mem_top_track_2.DFFR_3_.Q
rlabel metal3 32821 10948 32821 10948 0 mem_top_track_2.DFFR_4_.Q
rlabel metal1 35949 11118 35949 11118 0 mem_top_track_2.DFFR_5_.Q
rlabel metal1 20148 36006 20148 36006 0 mem_top_track_20.DFFR_0_.Q
rlabel metal2 21298 30498 21298 30498 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 23000 30634 23000 30634 0 mem_top_track_22.DFFR_0_.Q
rlabel metal1 29348 14382 29348 14382 0 mem_top_track_22.DFFR_1_.Q
rlabel metal1 16054 21964 16054 21964 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 14398 15470 14398 15470 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 23460 13294 23460 13294 0 mem_top_track_26.DFFR_0_.Q
rlabel metal1 20010 8976 20010 8976 0 mem_top_track_26.DFFR_1_.Q
rlabel metal2 6854 21148 6854 21148 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 34868 25942 34868 25942 0 mem_top_track_4.DFFR_0_.Q
rlabel metal1 36662 25670 36662 25670 0 mem_top_track_4.DFFR_1_.Q
rlabel metal1 34822 30158 34822 30158 0 mem_top_track_4.DFFR_2_.Q
rlabel metal1 21022 26452 21022 26452 0 mem_top_track_4.DFFR_3_.Q
rlabel metal1 21988 36074 21988 36074 0 mem_top_track_4.DFFR_4_.Q
rlabel metal1 20102 30124 20102 30124 0 mem_top_track_4.DFFR_5_.Q
rlabel metal1 19182 23732 19182 23732 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 13938 24276 13938 24276 0 mem_top_track_6.DFFR_1_.Q
rlabel metal1 33350 15538 33350 15538 0 mem_top_track_6.DFFR_2_.Q
rlabel metal2 36662 27200 36662 27200 0 mem_top_track_6.DFFR_3_.Q
rlabel metal1 32430 32742 32430 32742 0 mem_top_track_6.DFFR_4_.Q
rlabel metal1 34638 33286 34638 33286 0 mem_top_track_6.DFFR_5_.Q
rlabel metal1 33902 12206 33902 12206 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 10028 11866 10028 11866 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 9614 31994 9614 31994 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 9936 12954 9936 12954 0 mux_left_track_1.INVTX1_2_.out
rlabel metal1 16560 32946 16560 32946 0 mux_left_track_1.INVTX1_3_.out
rlabel metal1 13524 34510 13524 34510 0 mux_left_track_1.INVTX1_4_.out
rlabel metal1 13524 33286 13524 33286 0 mux_left_track_1.INVTX1_5_.out
rlabel metal1 9016 35122 9016 35122 0 mux_left_track_1.INVTX1_6_.out
rlabel metal1 10166 16490 10166 16490 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 7774 35258 7774 35258 0 mux_left_track_1.INVTX1_8_.out
rlabel metal2 12466 27132 12466 27132 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 14582 34646 14582 34646 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 36271 33966 36271 33966 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36386 33660 36386 33660 0 mux_left_track_1.out
rlabel metal2 16974 20910 16974 20910 0 mux_left_track_17.INVTX1_0_.out
rlabel metal2 12374 19074 12374 19074 0 mux_left_track_17.INVTX1_1_.out
rlabel metal1 30038 18360 30038 18360 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 33626 14586 33626 14586 0 mux_left_track_17.INVTX1_3_.out
rlabel metal2 35742 17408 35742 17408 0 mux_left_track_17.INVTX1_4_.out
rlabel metal1 19780 16218 19780 16218 0 mux_left_track_17.INVTX1_5_.out
rlabel metal2 31878 16609 31878 16609 0 mux_left_track_17.INVTX1_6_.out
rlabel metal1 18308 8330 18308 8330 0 mux_left_track_17.INVTX1_7_.out
rlabel metal2 14904 33388 14904 33388 0 mux_left_track_17.INVTX1_8_.out
rlabel metal1 18538 20366 18538 20366 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 31970 16558 31970 16558 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 35558 33439 35558 33439 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36478 34340 36478 34340 0 mux_left_track_17.out
rlabel metal1 12098 24718 12098 24718 0 mux_left_track_25.INVTX1_0_.out
rlabel metal1 15732 11866 15732 11866 0 mux_left_track_25.INVTX1_1_.out
rlabel metal1 12098 18326 12098 18326 0 mux_left_track_25.INVTX1_2_.out
rlabel metal1 25070 14280 25070 14280 0 mux_left_track_25.INVTX1_3_.out
rlabel metal2 14398 20434 14398 20434 0 mux_left_track_25.INVTX1_4_.out
rlabel metal1 17296 11322 17296 11322 0 mux_left_track_25.INVTX1_5_.out
rlabel metal1 22632 12274 22632 12274 0 mux_left_track_25.INVTX1_6_.out
rlabel metal2 16974 11662 16974 11662 0 mux_left_track_25.INVTX1_7_.out
rlabel metal2 10994 9316 10994 9316 0 mux_left_track_25.INVTX1_8_.out
rlabel metal1 19090 19278 19090 19278 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 19366 18326 19366 18326 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 2162 3060 2162 3060 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 2576 3026 2576 3026 0 mux_left_track_25.out
rlabel metal2 10902 21658 10902 21658 0 mux_left_track_33.INVTX1_0_.out
rlabel metal2 33350 15079 33350 15079 0 mux_left_track_33.INVTX1_1_.out
rlabel metal1 33856 16014 33856 16014 0 mux_left_track_33.INVTX1_2_.out
rlabel metal1 18216 12070 18216 12070 0 mux_left_track_33.INVTX1_3_.out
rlabel metal1 35880 14382 35880 14382 0 mux_left_track_33.INVTX1_4_.out
rlabel metal2 36294 17238 36294 17238 0 mux_left_track_33.INVTX1_5_.out
rlabel metal1 8372 31926 8372 31926 0 mux_left_track_33.INVTX1_6_.out
rlabel metal1 9982 18666 9982 18666 0 mux_left_track_33.INVTX1_7_.out
rlabel metal1 35052 16014 35052 16014 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 28474 17204 28474 17204 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 13754 19788 13754 19788 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 25024 19210 25024 19210 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 36202 19414 36202 19414 0 mux_left_track_33.out
rlabel metal1 14720 24718 14720 24718 0 mux_left_track_9.INVTX1_0_.out
rlabel metal2 23966 12143 23966 12143 0 mux_left_track_9.INVTX1_1_.out
rlabel metal2 33994 21216 33994 21216 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 37306 12308 37306 12308 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 34822 34034 34822 34034 0 mux_left_track_9.INVTX1_4_.out
rlabel metal1 17020 31994 17020 31994 0 mux_left_track_9.INVTX1_5_.out
rlabel metal2 12558 35666 12558 35666 0 mux_left_track_9.INVTX1_6_.out
rlabel metal1 10120 36346 10120 36346 0 mux_left_track_9.INVTX1_7_.out
rlabel metal1 15824 34510 15824 34510 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 35466 34816 35466 34816 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 13478 36550 13478 36550 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 16238 34408 16238 34408 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 8602 32844 8602 32844 0 mux_left_track_9.out
rlabel metal1 10534 33422 10534 33422 0 mux_right_track_0.INVTX1_3_.out
rlabel metal1 10120 21454 10120 21454 0 mux_right_track_0.INVTX1_4_.out
rlabel metal2 11178 28526 11178 28526 0 mux_right_track_0.INVTX1_5_.out
rlabel metal2 14398 27200 14398 27200 0 mux_right_track_0.INVTX1_6_.out
rlabel metal2 11638 26860 11638 26860 0 mux_right_track_0.INVTX1_7_.out
rlabel metal1 17020 21998 17020 21998 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11638 21522 11638 21522 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 14582 26418 14582 26418 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14536 32742 14536 32742 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 8924 32742 8924 32742 0 mux_right_track_0.out
rlabel metal1 30314 13838 30314 13838 0 mux_right_track_16.INVTX1_4_.out
rlabel metal2 25438 10336 25438 10336 0 mux_right_track_16.INVTX1_5_.out
rlabel metal1 14214 30770 14214 30770 0 mux_right_track_16.INVTX1_6_.out
rlabel metal1 18262 13498 18262 13498 0 mux_right_track_16.INVTX1_7_.out
rlabel metal1 15042 25160 15042 25160 0 mux_right_track_16.INVTX1_8_.out
rlabel metal1 35604 19414 35604 19414 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 30452 11186 30452 11186 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 38870 31790 38870 31790 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36800 35802 36800 35802 0 mux_right_track_16.out
rlabel metal1 8878 30770 8878 30770 0 mux_right_track_24.INVTX1_4_.out
rlabel metal1 36616 14518 36616 14518 0 mux_right_track_24.INVTX1_5_.out
rlabel metal2 15318 29648 15318 29648 0 mux_right_track_24.INVTX1_6_.out
rlabel metal1 9706 17238 9706 17238 0 mux_right_track_24.INVTX1_7_.out
rlabel metal2 22770 10540 22770 10540 0 mux_right_track_24.INVTX1_8_.out
rlabel metal2 20010 15742 20010 15742 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 12098 17544 12098 17544 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 36616 4114 36616 4114 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36938 3468 36938 3468 0 mux_right_track_24.out
rlabel metal2 16974 10234 16974 10234 0 mux_right_track_32.INVTX1_4_.out
rlabel metal1 25208 8602 25208 8602 0 mux_right_track_32.INVTX1_5_.out
rlabel metal1 27554 12274 27554 12274 0 mux_right_track_32.INVTX1_6_.out
rlabel metal2 17618 11356 17618 11356 0 mux_right_track_32.INVTX1_7_.out
rlabel metal2 15134 19040 15134 19040 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 25392 11662 25392 11662 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 24978 10574 24978 10574 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 22310 10166 22310 10166 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 19458 9180 19458 9180 0 mux_right_track_32.out
rlabel metal2 1702 36873 1702 36873 0 mux_right_track_8.INVTX1_4_.out
rlabel metal1 16882 11866 16882 11866 0 mux_right_track_8.INVTX1_5_.out
rlabel metal2 2438 35819 2438 35819 0 mux_right_track_8.INVTX1_6_.out
rlabel via2 1702 35717 1702 35717 0 mux_right_track_8.INVTX1_7_.out
rlabel metal1 20148 13362 20148 13362 0 mux_right_track_8.INVTX1_8_.out
rlabel metal1 16744 32810 16744 32810 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 2714 36448 2714 36448 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 27324 9554 27324 9554 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 28106 9146 28106 9146 0 mux_right_track_8.out
rlabel metal1 11454 22066 11454 22066 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 12834 35020 12834 35020 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 10948 32810 10948 32810 0 mux_top_track_0.INVTX1_3_.out
rlabel metal1 26634 20366 26634 20366 0 mux_top_track_0.INVTX1_5_.out
rlabel metal2 19918 23154 19918 23154 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11868 32946 11868 32946 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 34178 14042 34178 14042 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 33764 12614 33764 12614 0 mux_top_track_0.out
rlabel metal2 14720 19414 14720 19414 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 32062 15232 32062 15232 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 32568 4590 32568 4590 0 mux_top_track_10.out
rlabel metal2 35926 33422 35926 33422 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 37628 32878 37628 32878 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 37536 33082 37536 33082 0 mux_top_track_12.out
rlabel metal2 19274 14450 19274 14450 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 10902 15198 10902 15198 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 7728 12818 7728 12818 0 mux_top_track_14.out
rlabel metal1 10442 17714 10442 17714 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 9798 27302 9798 27302 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 8234 28322 8234 28322 0 mux_top_track_16.out
rlabel metal2 12098 19890 12098 19890 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13202 13940 13202 13940 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11408 9622 11408 9622 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 7130 8908 7130 8908 0 mux_top_track_18.out
rlabel metal1 29578 15470 29578 15470 0 mux_top_track_2.INVTX1_1_.out
rlabel metal2 31510 35292 31510 35292 0 mux_top_track_2.INVTX1_3_.out
rlabel metal2 36294 12053 36294 12053 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal3 15663 34612 15663 34612 0 mux_top_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 37214 11594 37214 11594 0 mux_top_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 36708 10166 36708 10166 0 mux_top_track_2.out
rlabel metal2 9798 34680 9798 34680 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11776 28730 11776 28730 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13754 35598 13754 35598 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 12466 36924 12466 36924 0 mux_top_track_20.out
rlabel metal2 27278 16320 27278 16320 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21252 11866 21252 11866 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28888 10642 28888 10642 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 29026 9146 29026 9146 0 mux_top_track_22.out
rlabel metal2 16376 18700 16376 18700 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10994 5678 10994 5678 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 8418 6086 8418 6086 0 mux_top_track_24.out
rlabel metal2 23138 10812 23138 10812 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20562 9350 20562 9350 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18308 7378 18308 7378 0 mux_top_track_26.out
rlabel metal1 11132 34510 11132 34510 0 mux_top_track_36.INVTX1_1_.out
rlabel metal1 6854 9622 6854 9622 0 mux_top_track_36.INVTX1_2_.out
rlabel metal2 8234 30192 8234 30192 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9338 23290 9338 23290 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8142 24786 8142 24786 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 7314 24378 7314 24378 0 mux_top_track_36.out
rlabel metal2 36294 14790 36294 14790 0 mux_top_track_4.INVTX1_2_.out
rlabel metal2 15594 20475 15594 20475 0 mux_top_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14858 29750 14858 29750 0 mux_top_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 9522 29818 9522 29818 0 mux_top_track_4.out
rlabel metal1 11132 15130 11132 15130 0 mux_top_track_6.INVTX1_0_.out
rlabel metal1 32522 10778 32522 10778 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 14490 16558 14490 16558 0 mux_top_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 35144 17646 35144 17646 0 mux_top_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 36340 17782 36340 17782 0 mux_top_track_6.out
rlabel metal2 36386 15062 36386 15062 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 36547 11866 36547 11866 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35006 11560 35006 11560 0 mux_top_track_8.out
rlabel metal2 1886 19516 1886 19516 0 net1
rlabel metal2 17066 2550 17066 2550 0 net10
rlabel metal1 37076 8330 37076 8330 0 net100
rlabel metal2 14858 36414 14858 36414 0 net101
rlabel metal1 36800 35258 36800 35258 0 net102
rlabel via3 35949 2652 35949 2652 0 net103
rlabel metal1 5474 36346 5474 36346 0 net104
rlabel metal2 18538 14297 18538 14297 0 net105
rlabel metal1 4048 37230 4048 37230 0 net106
rlabel metal1 37398 3162 37398 3162 0 net107
rlabel metal1 4255 14382 4255 14382 0 net108
rlabel metal1 25645 7854 25645 7854 0 net109
rlabel metal1 29256 2618 29256 2618 0 net11
rlabel metal2 1794 19635 1794 19635 0 net110
rlabel metal1 17480 2414 17480 2414 0 net111
rlabel metal2 1610 21692 1610 21692 0 net112
rlabel metal2 16790 2618 16790 2618 0 net113
rlabel metal2 5014 25228 5014 25228 0 net114
rlabel metal2 33074 36550 33074 36550 0 net115
rlabel metal2 2990 33898 2990 33898 0 net116
rlabel metal1 29164 8806 29164 8806 0 net117
rlabel metal1 13662 26316 13662 26316 0 net118
rlabel metal1 36961 5678 36961 5678 0 net119
rlabel metal1 27784 37094 27784 37094 0 net12
rlabel metal1 14306 27540 14306 27540 0 net120
rlabel metal1 37996 35054 37996 35054 0 net121
rlabel metal1 36018 36584 36018 36584 0 net122
rlabel metal1 37490 2958 37490 2958 0 net123
rlabel metal2 13662 36958 13662 36958 0 net124
rlabel metal1 30590 2482 30590 2482 0 net125
rlabel metal2 5566 4556 5566 4556 0 net126
rlabel metal2 14950 4794 14950 4794 0 net127
rlabel via3 38203 20332 38203 20332 0 net128
rlabel metal1 38088 28390 38088 28390 0 net129
rlabel metal1 6762 37230 6762 37230 0 net13
rlabel metal2 32338 2618 32338 2618 0 net130
rlabel metal1 2185 24174 2185 24174 0 net131
rlabel metal1 37766 10642 37766 10642 0 net132
rlabel metal1 3772 32402 3772 32402 0 net133
rlabel metal1 37536 18394 37536 18394 0 net134
rlabel metal1 38548 34578 38548 34578 0 net135
rlabel metal1 37490 2380 37490 2380 0 net136
rlabel metal1 37720 35258 37720 35258 0 net137
rlabel metal1 6946 12886 6946 12886 0 net138
rlabel metal2 1610 31654 1610 31654 0 net139
rlabel metal1 25208 9894 25208 9894 0 net14
rlabel metal1 3680 3570 3680 3570 0 net140
rlabel metal2 38318 4369 38318 4369 0 net141
rlabel metal1 33534 13838 33534 13838 0 net142
rlabel metal1 37720 11186 37720 11186 0 net143
rlabel metal2 13110 30124 13110 30124 0 net144
rlabel metal1 37306 21046 37306 21046 0 net145
rlabel metal1 37030 9622 37030 9622 0 net146
rlabel metal2 33534 14722 33534 14722 0 net147
rlabel metal2 37490 31008 37490 31008 0 net148
rlabel metal2 10258 15776 10258 15776 0 net149
rlabel metal1 8694 29138 8694 29138 0 net15
rlabel metal1 8786 26350 8786 26350 0 net150
rlabel metal2 13294 13600 13294 13600 0 net151
rlabel metal2 20838 9724 20838 9724 0 net152
rlabel metal2 12190 12988 12190 12988 0 net153
rlabel metal2 9982 29920 9982 29920 0 net154
rlabel metal1 20976 11186 20976 11186 0 net155
rlabel metal1 8648 22542 8648 22542 0 net156
rlabel metal1 11408 23630 11408 23630 0 net157
rlabel metal2 24702 10336 24702 10336 0 net158
rlabel metal2 12558 36380 12558 36380 0 net159
rlabel metal2 23138 2482 23138 2482 0 net16
rlabel metal2 13110 19550 13110 19550 0 net160
rlabel metal1 29394 17272 29394 17272 0 net161
rlabel metal1 36708 31858 36708 31858 0 net162
rlabel metal2 35466 12852 35466 12852 0 net163
rlabel metal1 7406 35598 7406 35598 0 net164
rlabel metal1 25024 30770 25024 30770 0 net165
rlabel metal2 14582 20128 14582 20128 0 net166
rlabel metal2 1886 17476 1886 17476 0 net17
rlabel metal1 3864 2618 3864 2618 0 net18
rlabel metal1 30728 36754 30728 36754 0 net19
rlabel metal1 5336 25874 5336 25874 0 net2
rlabel metal1 12006 2380 12006 2380 0 net20
rlabel metal2 20470 36516 20470 36516 0 net21
rlabel metal2 17894 3264 17894 3264 0 net22
rlabel metal1 32338 35632 32338 35632 0 net23
rlabel metal3 35397 37332 35397 37332 0 net24
rlabel metal2 37582 36533 37582 36533 0 net25
rlabel metal1 16928 31790 16928 31790 0 net26
rlabel metal1 37674 12682 37674 12682 0 net27
rlabel metal1 32844 12206 32844 12206 0 net28
rlabel metal2 21482 17476 21482 17476 0 net29
rlabel metal1 1932 5746 1932 5746 0 net3
rlabel metal1 30176 10574 30176 10574 0 net30
rlabel metal1 38732 37230 38732 37230 0 net31
rlabel metal1 38594 33354 38594 33354 0 net32
rlabel metal2 15318 35870 15318 35870 0 net33
rlabel metal1 13110 18734 13110 18734 0 net34
rlabel metal1 37674 8500 37674 8500 0 net35
rlabel metal1 13110 33524 13110 33524 0 net36
rlabel metal1 9798 32878 9798 32878 0 net37
rlabel metal1 34178 32912 34178 32912 0 net38
rlabel metal1 18561 2550 18561 2550 0 net39
rlabel metal1 34316 3026 34316 3026 0 net4
rlabel metal1 4600 3978 4600 3978 0 net40
rlabel metal1 7268 2550 7268 2550 0 net41
rlabel metal1 35328 3706 35328 3706 0 net42
rlabel metal2 8510 14994 8510 14994 0 net43
rlabel metal1 37996 21862 37996 21862 0 net44
rlabel metal1 32660 13430 32660 13430 0 net45
rlabel metal2 17250 35020 17250 35020 0 net46
rlabel metal1 4462 2482 4462 2482 0 net47
rlabel metal1 33212 3570 33212 3570 0 net48
rlabel metal1 36754 11628 36754 11628 0 net49
rlabel metal1 17710 2278 17710 2278 0 net5
rlabel metal1 7544 21998 7544 21998 0 net50
rlabel metal1 5934 30702 5934 30702 0 net51
rlabel metal1 7498 21522 7498 21522 0 net52
rlabel metal1 5428 21114 5428 21114 0 net53
rlabel metal1 9246 31790 9246 31790 0 net54
rlabel metal2 36156 30396 36156 30396 0 net55
rlabel metal1 11316 2618 11316 2618 0 net56
rlabel metal2 8326 18870 8326 18870 0 net57
rlabel metal1 23598 2618 23598 2618 0 net58
rlabel metal1 4002 3706 4002 3706 0 net59
rlabel metal2 11684 19516 11684 19516 0 net6
rlabel metal1 4646 4794 4646 4794 0 net60
rlabel metal1 1610 34952 1610 34952 0 net61
rlabel metal1 7590 35088 7590 35088 0 net62
rlabel metal1 20102 37128 20102 37128 0 net63
rlabel metal2 9338 30532 9338 30532 0 net64
rlabel metal1 6762 2618 6762 2618 0 net65
rlabel metal1 3588 2550 3588 2550 0 net66
rlabel metal2 1610 12886 1610 12886 0 net67
rlabel metal2 22034 36992 22034 36992 0 net68
rlabel metal1 19826 2618 19826 2618 0 net69
rlabel metal1 1840 18734 1840 18734 0 net7
rlabel metal1 35466 7514 35466 7514 0 net70
rlabel metal1 6164 31314 6164 31314 0 net71
rlabel metal2 9522 10642 9522 10642 0 net72
rlabel metal1 7544 10030 7544 10030 0 net73
rlabel metal1 16790 11730 16790 11730 0 net74
rlabel metal1 22770 2550 22770 2550 0 net75
rlabel metal1 38226 14450 38226 14450 0 net76
rlabel metal1 23920 2278 23920 2278 0 net77
rlabel metal2 6486 36193 6486 36193 0 net78
rlabel metal1 26174 36754 26174 36754 0 net79
rlabel metal1 17434 36686 17434 36686 0 net8
rlabel metal1 6486 32878 6486 32878 0 net80
rlabel metal1 8556 35054 8556 35054 0 net81
rlabel metal1 28244 2550 28244 2550 0 net82
rlabel metal2 8786 12852 8786 12852 0 net83
rlabel metal1 1610 7888 1610 7888 0 net84
rlabel metal2 38042 33082 38042 33082 0 net85
rlabel metal2 20838 16745 20838 16745 0 net86
rlabel metal1 9614 2482 9614 2482 0 net87
rlabel metal2 1610 2618 1610 2618 0 net88
rlabel metal1 38042 13192 38042 13192 0 net89
rlabel metal1 1978 22032 1978 22032 0 net9
rlabel metal1 14766 37162 14766 37162 0 net90
rlabel metal1 37536 30226 37536 30226 0 net91
rlabel metal1 36570 12342 36570 12342 0 net92
rlabel metal3 32407 36380 32407 36380 0 net93
rlabel metal1 19688 2482 19688 2482 0 net94
rlabel metal2 36202 36941 36202 36941 0 net95
rlabel metal1 37950 13294 37950 13294 0 net96
rlabel metal2 36018 6188 36018 6188 0 net97
rlabel metal1 2185 30702 2185 30702 0 net98
rlabel metal2 10810 16252 10810 16252 0 net99
rlabel metal2 19366 1588 19366 1588 0 pReset
rlabel metal2 35466 37551 35466 37551 0 prog_clk
rlabel metal3 38786 6868 38786 6868 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1234 36108 1234 36108 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1234 10948 1234 10948 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7130 1588 7130 1588 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 13570 1588 13570 1588 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel via2 38318 25891 38318 25891 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 22586 1588 22586 1588 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 29716 37298 29716 37298 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 31234 37196 31234 37196 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 690 38294 690 38294 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 5382 36788 5382 36788 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 27094 1588 27094 1588 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal3 1234 10268 1234 10268 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
