magic
tech sky130A
magscale 1 2
timestamp 1674174591
<< viali >>
rect 4248 37417 4282 37451
rect 11069 37417 11103 37451
rect 1869 37281 1903 37315
rect 7021 37281 7055 37315
rect 9597 37281 9631 37315
rect 11989 37281 12023 37315
rect 1593 37213 1627 37247
rect 3985 37213 4019 37247
rect 6745 37213 6779 37247
rect 9321 37213 9355 37247
rect 11713 37213 11747 37247
rect 14289 37213 14323 37247
rect 15577 37213 15611 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 19625 37213 19659 37247
rect 19901 37213 19935 37247
rect 20085 37213 20119 37247
rect 22201 37213 22235 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 26065 37213 26099 37247
rect 27997 37213 28031 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 35081 37213 35115 37247
rect 36921 37213 36955 37247
rect 38025 37213 38059 37247
rect 3341 37077 3375 37111
rect 5733 37077 5767 37111
rect 8493 37077 8527 37111
rect 13461 37077 13495 37111
rect 14473 37077 14507 37111
rect 15761 37077 15795 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 19441 37077 19475 37111
rect 20269 37077 20303 37111
rect 22017 37077 22051 37111
rect 22661 37077 22695 37111
rect 24777 37077 24811 37111
rect 25881 37077 25915 37111
rect 27813 37077 27847 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 34897 37077 34931 37111
rect 36737 37077 36771 37111
rect 38209 37077 38243 37111
rect 5917 36873 5951 36907
rect 15945 36873 15979 36907
rect 16865 36873 16899 36907
rect 14473 36805 14507 36839
rect 1593 36737 1627 36771
rect 4169 36737 4203 36771
rect 17049 36737 17083 36771
rect 17509 36737 17543 36771
rect 18153 36737 18187 36771
rect 18797 36737 18831 36771
rect 19625 36737 19659 36771
rect 37657 36737 37691 36771
rect 38301 36737 38335 36771
rect 1869 36669 1903 36703
rect 3617 36669 3651 36703
rect 4445 36669 4479 36703
rect 7021 36669 7055 36703
rect 7297 36669 7331 36703
rect 8769 36669 8803 36703
rect 9321 36669 9355 36703
rect 9597 36669 9631 36703
rect 11897 36669 11931 36703
rect 12173 36669 12207 36703
rect 14197 36669 14231 36703
rect 18245 36669 18279 36703
rect 18889 36601 18923 36635
rect 38117 36601 38151 36635
rect 11069 36533 11103 36567
rect 13645 36533 13679 36567
rect 17601 36533 17635 36567
rect 19441 36533 19475 36567
rect 37473 36533 37507 36567
rect 10149 36329 10183 36363
rect 15761 36329 15795 36363
rect 17969 36329 18003 36363
rect 14473 36261 14507 36295
rect 1593 36193 1627 36227
rect 1869 36193 1903 36227
rect 4445 36193 4479 36227
rect 6745 36193 6779 36227
rect 8493 36193 8527 36227
rect 10701 36193 10735 36227
rect 9137 36125 9171 36159
rect 9965 36125 9999 36159
rect 13369 36125 13403 36159
rect 14657 36125 14691 36159
rect 15117 36125 15151 36159
rect 15945 36125 15979 36159
rect 16589 36125 16623 36159
rect 17049 36125 17083 36159
rect 17509 36125 17543 36159
rect 18521 36125 18555 36159
rect 38301 36125 38335 36159
rect 4721 36057 4755 36091
rect 7021 36057 7055 36091
rect 10977 36057 11011 36091
rect 17141 36057 17175 36091
rect 3341 35989 3375 36023
rect 6193 35989 6227 36023
rect 9321 35989 9355 36023
rect 12449 35989 12483 36023
rect 13185 35989 13219 36023
rect 15209 35989 15243 36023
rect 16405 35989 16439 36023
rect 17601 35989 17635 36023
rect 18337 35989 18371 36023
rect 38117 35989 38151 36023
rect 5917 35785 5951 35819
rect 14657 35785 14691 35819
rect 15209 35785 15243 35819
rect 1869 35649 1903 35683
rect 5733 35649 5767 35683
rect 6837 35649 6871 35683
rect 14105 35649 14139 35683
rect 14565 35649 14599 35683
rect 15393 35649 15427 35683
rect 15853 35649 15887 35683
rect 16865 35649 16899 35683
rect 17509 35649 17543 35683
rect 2145 35581 2179 35615
rect 3065 35581 3099 35615
rect 3341 35581 3375 35615
rect 7113 35581 7147 35615
rect 8585 35581 8619 35615
rect 9137 35581 9171 35615
rect 9413 35581 9447 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 13461 35581 13495 35615
rect 13921 35513 13955 35547
rect 4813 35445 4847 35479
rect 10885 35445 10919 35479
rect 15945 35445 15979 35479
rect 16957 35445 16991 35479
rect 17601 35445 17635 35479
rect 4708 35241 4742 35275
rect 22753 35241 22787 35275
rect 6193 35173 6227 35207
rect 17417 35173 17451 35207
rect 1593 35105 1627 35139
rect 1869 35105 1903 35139
rect 4445 35105 4479 35139
rect 6653 35105 6687 35139
rect 9137 35105 9171 35139
rect 9413 35105 9447 35139
rect 14289 35105 14323 35139
rect 11529 35037 11563 35071
rect 16497 35037 16531 35071
rect 17601 35037 17635 35071
rect 22937 35037 22971 35071
rect 38025 35037 38059 35071
rect 6929 34969 6963 35003
rect 11805 34969 11839 35003
rect 14565 34969 14599 35003
rect 16589 34969 16623 35003
rect 3341 34901 3375 34935
rect 8401 34901 8435 34935
rect 10885 34901 10919 34935
rect 13277 34901 13311 34935
rect 16037 34901 16071 34935
rect 38209 34901 38243 34935
rect 14841 34697 14875 34731
rect 18245 34697 18279 34731
rect 2145 34629 2179 34663
rect 1869 34561 1903 34595
rect 2789 34561 2823 34595
rect 4169 34561 4203 34595
rect 6561 34561 6595 34595
rect 10333 34561 10367 34595
rect 10793 34561 10827 34595
rect 11713 34561 11747 34595
rect 14197 34561 14231 34595
rect 14749 34561 14783 34595
rect 15393 34561 15427 34595
rect 15485 34561 15519 34595
rect 16037 34561 16071 34595
rect 16865 34561 16899 34595
rect 17509 34561 17543 34595
rect 18153 34561 18187 34595
rect 3065 34493 3099 34527
rect 5917 34493 5951 34527
rect 7849 34493 7883 34527
rect 10885 34493 10919 34527
rect 11989 34493 12023 34527
rect 13461 34493 13495 34527
rect 16957 34493 16991 34527
rect 6745 34425 6779 34459
rect 16129 34425 16163 34459
rect 4432 34357 4466 34391
rect 8112 34357 8146 34391
rect 9597 34357 9631 34391
rect 10149 34357 10183 34391
rect 14197 34357 14231 34391
rect 17601 34357 17635 34391
rect 2881 34153 2915 34187
rect 7100 34153 7134 34187
rect 11792 34153 11826 34187
rect 18061 34153 18095 34187
rect 35909 34153 35943 34187
rect 8585 34085 8619 34119
rect 10885 34085 10919 34119
rect 16773 34085 16807 34119
rect 3985 34017 4019 34051
rect 6009 34017 6043 34051
rect 9137 34017 9171 34051
rect 11529 34017 11563 34051
rect 14381 34017 14415 34051
rect 15025 34017 15059 34051
rect 1869 33949 1903 33983
rect 2789 33949 2823 33983
rect 6837 33949 6871 33983
rect 13553 33949 13587 33983
rect 15669 33949 15703 33983
rect 17325 33949 17359 33983
rect 17969 33949 18003 33983
rect 18613 33949 18647 33983
rect 36093 33949 36127 33983
rect 2145 33881 2179 33915
rect 4261 33881 4295 33915
rect 9413 33881 9447 33915
rect 14473 33881 14507 33915
rect 16221 33881 16255 33915
rect 16313 33881 16347 33915
rect 15485 33813 15519 33847
rect 17417 33813 17451 33847
rect 18705 33813 18739 33847
rect 3801 33609 3835 33643
rect 6009 33609 6043 33643
rect 14013 33609 14047 33643
rect 16037 33609 16071 33643
rect 16865 33609 16899 33643
rect 2329 33541 2363 33575
rect 9873 33541 9907 33575
rect 17877 33541 17911 33575
rect 2053 33473 2087 33507
rect 4261 33473 4295 33507
rect 6561 33473 6595 33507
rect 7205 33473 7239 33507
rect 7297 33473 7331 33507
rect 10333 33473 10367 33507
rect 10977 33473 11011 33507
rect 11713 33473 11747 33507
rect 13921 33473 13955 33507
rect 14565 33473 14599 33507
rect 15209 33473 15243 33507
rect 16221 33473 16255 33507
rect 20177 33473 20211 33507
rect 31493 33473 31527 33507
rect 38025 33473 38059 33507
rect 4537 33405 4571 33439
rect 7849 33405 7883 33439
rect 8125 33405 8159 33439
rect 11989 33405 12023 33439
rect 13461 33405 13495 33439
rect 17785 33405 17819 33439
rect 11069 33337 11103 33371
rect 14657 33337 14691 33371
rect 18337 33337 18371 33371
rect 38209 33337 38243 33371
rect 6653 33269 6687 33303
rect 10425 33269 10459 33303
rect 15301 33269 15335 33303
rect 20269 33269 20303 33303
rect 31585 33269 31619 33303
rect 1777 33065 1811 33099
rect 4077 33065 4111 33099
rect 6824 33065 6858 33099
rect 17601 32997 17635 33031
rect 24869 32997 24903 33031
rect 6561 32929 6595 32963
rect 11253 32929 11287 32963
rect 1593 32861 1627 32895
rect 2329 32861 2363 32895
rect 3157 32861 3191 32895
rect 3985 32861 4019 32895
rect 4629 32861 4663 32895
rect 5273 32861 5307 32895
rect 5917 32861 5951 32895
rect 9137 32861 9171 32895
rect 9781 32861 9815 32895
rect 10425 32861 10459 32895
rect 13645 32861 13679 32895
rect 14565 32861 14599 32895
rect 15025 32861 15059 32895
rect 16221 32861 16255 32895
rect 16865 32861 16899 32895
rect 17509 32861 17543 32895
rect 21557 32861 21591 32895
rect 22201 32861 22235 32895
rect 22661 32861 22695 32895
rect 24777 32861 24811 32895
rect 32321 32861 32355 32895
rect 8585 32793 8619 32827
rect 10517 32793 10551 32827
rect 11529 32793 11563 32827
rect 2421 32725 2455 32759
rect 2973 32725 3007 32759
rect 4721 32725 4755 32759
rect 5365 32725 5399 32759
rect 6009 32725 6043 32759
rect 9229 32725 9263 32759
rect 9873 32725 9907 32759
rect 13001 32725 13035 32759
rect 13461 32725 13495 32759
rect 14381 32725 14415 32759
rect 15117 32725 15151 32759
rect 16313 32725 16347 32759
rect 16957 32725 16991 32759
rect 21373 32725 21407 32759
rect 22017 32725 22051 32759
rect 22753 32725 22787 32759
rect 32413 32725 32447 32759
rect 10977 32521 11011 32555
rect 14013 32521 14047 32555
rect 15945 32521 15979 32555
rect 34345 32521 34379 32555
rect 38117 32521 38151 32555
rect 8033 32453 8067 32487
rect 33701 32453 33735 32487
rect 2053 32385 2087 32419
rect 4997 32385 5031 32419
rect 5641 32385 5675 32419
rect 5733 32385 5767 32419
rect 6561 32385 6595 32419
rect 9781 32385 9815 32419
rect 10425 32385 10459 32419
rect 10885 32385 10919 32419
rect 11713 32385 11747 32419
rect 13921 32385 13955 32419
rect 14565 32385 14599 32419
rect 15209 32385 15243 32419
rect 15853 32385 15887 32419
rect 17049 32385 17083 32419
rect 17509 32385 17543 32419
rect 18889 32385 18923 32419
rect 19533 32385 19567 32419
rect 22569 32385 22603 32419
rect 23949 32385 23983 32419
rect 28457 32385 28491 32419
rect 32321 32385 32355 32419
rect 33609 32385 33643 32419
rect 34253 32385 34287 32419
rect 38301 32385 38335 32419
rect 2697 32317 2731 32351
rect 2973 32317 3007 32351
rect 7757 32317 7791 32351
rect 14657 32317 14691 32351
rect 17601 32317 17635 32351
rect 22385 32317 22419 32351
rect 4445 32249 4479 32283
rect 16865 32249 16899 32283
rect 24041 32249 24075 32283
rect 2145 32181 2179 32215
rect 5089 32181 5123 32215
rect 6653 32181 6687 32215
rect 10241 32181 10275 32215
rect 11976 32181 12010 32215
rect 13461 32181 13495 32215
rect 15301 32181 15335 32215
rect 18705 32181 18739 32215
rect 19625 32181 19659 32215
rect 22845 32181 22879 32215
rect 28549 32181 28583 32215
rect 32413 32181 32447 32215
rect 3341 31977 3375 32011
rect 15025 31977 15059 32011
rect 15669 31977 15703 32011
rect 16313 31977 16347 32011
rect 16957 31977 16991 32011
rect 22385 31977 22419 32011
rect 9597 31909 9631 31943
rect 13645 31909 13679 31943
rect 18705 31909 18739 31943
rect 1593 31841 1627 31875
rect 1869 31841 1903 31875
rect 4905 31841 4939 31875
rect 5181 31841 5215 31875
rect 7481 31841 7515 31875
rect 11345 31841 11379 31875
rect 14381 31841 14415 31875
rect 19625 31841 19659 31875
rect 20545 31841 20579 31875
rect 22201 31841 22235 31875
rect 3985 31773 4019 31807
rect 4077 31773 4111 31807
rect 6929 31773 6963 31807
rect 7389 31773 7423 31807
rect 9781 31773 9815 31807
rect 10241 31773 10275 31807
rect 10333 31773 10367 31807
rect 13553 31773 13587 31807
rect 14289 31773 14323 31807
rect 14933 31773 14967 31807
rect 15577 31773 15611 31807
rect 16221 31773 16255 31807
rect 16865 31773 16899 31807
rect 18889 31773 18923 31807
rect 19533 31773 19567 31807
rect 22017 31773 22051 31807
rect 25145 31773 25179 31807
rect 25789 31773 25823 31807
rect 8401 31705 8435 31739
rect 11621 31705 11655 31739
rect 20269 31705 20303 31739
rect 20361 31705 20395 31739
rect 13093 31637 13127 31671
rect 25237 31637 25271 31671
rect 1961 31433 1995 31467
rect 5733 31433 5767 31467
rect 14197 31433 14231 31467
rect 16957 31433 16991 31467
rect 18889 31365 18923 31399
rect 20085 31365 20119 31399
rect 1869 31297 1903 31331
rect 2697 31297 2731 31331
rect 4997 31297 5031 31331
rect 5641 31297 5675 31331
rect 12357 31297 12391 31331
rect 12817 31297 12851 31331
rect 13461 31297 13495 31331
rect 14105 31297 14139 31331
rect 14749 31297 14783 31331
rect 15393 31297 15427 31331
rect 16037 31297 16071 31331
rect 16865 31297 16899 31331
rect 18245 31297 18279 31331
rect 25053 31297 25087 31331
rect 25697 31297 25731 31331
rect 32321 31297 32355 31331
rect 2973 31229 3007 31263
rect 6561 31229 6595 31263
rect 6837 31229 6871 31263
rect 9137 31229 9171 31263
rect 9413 31229 9447 31263
rect 11161 31229 11195 31263
rect 18797 31229 18831 31263
rect 19993 31229 20027 31263
rect 25513 31229 25547 31263
rect 13553 31161 13587 31195
rect 15485 31161 15519 31195
rect 19349 31161 19383 31195
rect 20545 31161 20579 31195
rect 25881 31161 25915 31195
rect 4445 31093 4479 31127
rect 5089 31093 5123 31127
rect 8309 31093 8343 31127
rect 12173 31093 12207 31127
rect 12909 31093 12943 31127
rect 14841 31093 14875 31127
rect 16129 31093 16163 31127
rect 18061 31093 18095 31127
rect 24869 31093 24903 31127
rect 32413 31093 32447 31127
rect 10609 30889 10643 30923
rect 11989 30889 12023 30923
rect 13277 30889 13311 30923
rect 14381 30889 14415 30923
rect 24685 30889 24719 30923
rect 7849 30821 7883 30855
rect 27353 30821 27387 30855
rect 2145 30753 2179 30787
rect 9413 30753 9447 30787
rect 10149 30753 10183 30787
rect 26157 30753 26191 30787
rect 1869 30685 1903 30719
rect 2789 30685 2823 30719
rect 3985 30685 4019 30719
rect 4629 30685 4663 30719
rect 6009 30685 6043 30719
rect 6653 30685 6687 30719
rect 7113 30685 7147 30719
rect 7757 30685 7791 30719
rect 8585 30685 8619 30719
rect 9321 30685 9355 30719
rect 9965 30685 9999 30719
rect 11253 30685 11287 30719
rect 11897 30685 11931 30719
rect 12541 30685 12575 30719
rect 12633 30685 12667 30719
rect 13185 30685 13219 30719
rect 14289 30685 14323 30719
rect 14933 30685 14967 30719
rect 15761 30685 15795 30719
rect 16497 30685 16531 30719
rect 19625 30685 19659 30719
rect 24593 30685 24627 30719
rect 26617 30685 26651 30719
rect 27261 30685 27295 30719
rect 18245 30617 18279 30651
rect 18337 30617 18371 30651
rect 18889 30617 18923 30651
rect 25513 30617 25547 30651
rect 25605 30617 25639 30651
rect 2881 30549 2915 30583
rect 4077 30549 4111 30583
rect 4721 30549 4755 30583
rect 5825 30549 5859 30583
rect 6469 30549 6503 30583
rect 7205 30549 7239 30583
rect 8401 30549 8435 30583
rect 11069 30549 11103 30583
rect 15025 30549 15059 30583
rect 15577 30549 15611 30583
rect 16313 30549 16347 30583
rect 19441 30549 19475 30583
rect 26709 30549 26743 30583
rect 5825 30345 5859 30379
rect 18705 30345 18739 30379
rect 13461 30277 13495 30311
rect 14381 30277 14415 30311
rect 17693 30277 17727 30311
rect 19809 30277 19843 30311
rect 25513 30277 25547 30311
rect 25605 30277 25639 30311
rect 26157 30277 26191 30311
rect 1869 30209 1903 30243
rect 4537 30209 4571 30243
rect 4997 30209 5031 30243
rect 6009 30209 6043 30243
rect 13001 30209 13035 30243
rect 13921 30209 13955 30243
rect 14933 30209 14967 30243
rect 15669 30209 15703 30243
rect 17601 30209 17635 30243
rect 18613 30209 18647 30243
rect 24869 30209 24903 30243
rect 28089 30209 28123 30243
rect 34437 30209 34471 30243
rect 38301 30209 38335 30243
rect 2145 30141 2179 30175
rect 3893 30141 3927 30175
rect 6653 30141 6687 30175
rect 6929 30141 6963 30175
rect 8861 30141 8895 30175
rect 9137 30141 9171 30175
rect 11713 30141 11747 30175
rect 15485 30141 15519 30175
rect 19717 30141 19751 30175
rect 28181 30141 28215 30175
rect 14013 30073 14047 30107
rect 15853 30073 15887 30107
rect 20269 30073 20303 30107
rect 24685 30073 24719 30107
rect 34253 30073 34287 30107
rect 4353 30005 4387 30039
rect 5089 30005 5123 30039
rect 8401 30005 8435 30039
rect 10609 30005 10643 30039
rect 12817 30005 12851 30039
rect 14749 30005 14783 30039
rect 38117 30005 38151 30039
rect 7297 29801 7331 29835
rect 12081 29801 12115 29835
rect 13553 29733 13587 29767
rect 17509 29733 17543 29767
rect 2145 29665 2179 29699
rect 3065 29665 3099 29699
rect 4629 29665 4663 29699
rect 8125 29665 8159 29699
rect 17325 29665 17359 29699
rect 1869 29597 1903 29631
rect 2789 29597 2823 29631
rect 4169 29597 4203 29631
rect 7481 29597 7515 29631
rect 7941 29597 7975 29631
rect 9137 29597 9171 29631
rect 11437 29597 11471 29631
rect 11621 29597 11655 29631
rect 12633 29597 12667 29631
rect 13737 29597 13771 29631
rect 14657 29597 14691 29631
rect 15301 29597 15335 29631
rect 17141 29597 17175 29631
rect 18889 29597 18923 29631
rect 19625 29607 19659 29641
rect 20269 29597 20303 29631
rect 21557 29597 21591 29631
rect 24777 29597 24811 29631
rect 4905 29529 4939 29563
rect 6653 29529 6687 29563
rect 9413 29529 9447 29563
rect 19717 29529 19751 29563
rect 3985 29461 4019 29495
rect 8585 29461 8619 29495
rect 10885 29461 10919 29495
rect 12725 29461 12759 29495
rect 14473 29461 14507 29495
rect 15117 29461 15151 29495
rect 18705 29461 18739 29495
rect 20361 29461 20395 29495
rect 20913 29461 20947 29495
rect 21649 29461 21683 29495
rect 24593 29461 24627 29495
rect 4721 29257 4755 29291
rect 6009 29257 6043 29291
rect 21097 29257 21131 29291
rect 23489 29257 23523 29291
rect 10609 29189 10643 29223
rect 1961 29121 1995 29155
rect 3985 29121 4019 29155
rect 4905 29121 4939 29155
rect 5549 29121 5583 29155
rect 7113 29121 7147 29155
rect 7297 29121 7331 29155
rect 8217 29121 8251 29155
rect 11713 29121 11747 29155
rect 14197 29121 14231 29155
rect 15025 29121 15059 29155
rect 16037 29121 16071 29155
rect 17049 29121 17083 29155
rect 17785 29121 17819 29155
rect 18889 29121 18923 29155
rect 20177 29121 20211 29155
rect 21281 29121 21315 29155
rect 22201 29121 22235 29155
rect 22753 29121 22787 29155
rect 23397 29121 23431 29155
rect 25237 29121 25271 29155
rect 38301 29121 38335 29155
rect 5365 29053 5399 29087
rect 9965 29053 9999 29087
rect 10517 29053 10551 29087
rect 11161 29053 11195 29087
rect 11989 29053 12023 29087
rect 13737 29053 13771 29087
rect 17969 29053 18003 29087
rect 18429 29053 18463 29087
rect 19993 29053 20027 29087
rect 7481 28985 7515 29019
rect 14289 28985 14323 29019
rect 14841 28985 14875 29019
rect 15853 28985 15887 29019
rect 16865 28985 16899 29019
rect 18981 28985 19015 29019
rect 20637 28985 20671 29019
rect 22017 28985 22051 29019
rect 25329 28985 25363 29019
rect 38117 28985 38151 29019
rect 2224 28917 2258 28951
rect 8480 28917 8514 28951
rect 22845 28917 22879 28951
rect 8401 28713 8435 28747
rect 16681 28713 16715 28747
rect 7665 28645 7699 28679
rect 17969 28645 18003 28679
rect 21741 28645 21775 28679
rect 1869 28577 1903 28611
rect 4997 28577 5031 28611
rect 6193 28577 6227 28611
rect 10057 28577 10091 28611
rect 10333 28577 10367 28611
rect 12081 28577 12115 28611
rect 13185 28577 13219 28611
rect 19533 28577 19567 28611
rect 19993 28577 20027 28611
rect 20637 28577 20671 28611
rect 20821 28577 20855 28611
rect 22753 28577 22787 28611
rect 22937 28577 22971 28611
rect 1593 28509 1627 28543
rect 4169 28509 4203 28543
rect 4813 28509 4847 28543
rect 5917 28509 5951 28543
rect 8585 28509 8619 28543
rect 9413 28509 9447 28543
rect 12541 28509 12575 28543
rect 12725 28509 12759 28543
rect 14749 28509 14783 28543
rect 15761 28509 15795 28543
rect 16865 28509 16899 28543
rect 17325 28509 17359 28543
rect 18153 28509 18187 28543
rect 18797 28509 18831 28543
rect 21925 28509 21959 28543
rect 17417 28441 17451 28475
rect 19625 28441 19659 28475
rect 3341 28373 3375 28407
rect 4261 28373 4295 28407
rect 5457 28373 5491 28407
rect 9505 28373 9539 28407
rect 14841 28373 14875 28407
rect 15853 28373 15887 28407
rect 18613 28373 18647 28407
rect 21281 28373 21315 28407
rect 23397 28373 23431 28407
rect 11069 28169 11103 28203
rect 13461 28169 13495 28203
rect 22661 28169 22695 28203
rect 1869 28101 1903 28135
rect 4353 28101 4387 28135
rect 9045 28101 9079 28135
rect 9965 28101 9999 28135
rect 20821 28101 20855 28135
rect 20913 28101 20947 28135
rect 23213 28101 23247 28135
rect 4077 28033 4111 28067
rect 7021 28033 7055 28067
rect 10977 28033 11011 28067
rect 11713 28033 11747 28067
rect 14381 28033 14415 28067
rect 15209 28033 15243 28067
rect 15853 28033 15887 28067
rect 17417 28033 17451 28067
rect 19625 28033 19659 28067
rect 20085 28033 20119 28067
rect 22017 28033 22051 28067
rect 22201 28033 22235 28067
rect 23121 28033 23155 28067
rect 24961 28033 24995 28067
rect 1593 27965 1627 27999
rect 3617 27965 3651 27999
rect 5825 27965 5859 27999
rect 7304 27965 7338 27999
rect 9873 27965 9907 27999
rect 11989 27965 12023 27999
rect 15669 27965 15703 27999
rect 17233 27965 17267 27999
rect 18521 27965 18555 27999
rect 21465 27965 21499 27999
rect 23765 27965 23799 27999
rect 10425 27897 10459 27931
rect 14473 27829 14507 27863
rect 15025 27829 15059 27863
rect 16313 27829 16347 27863
rect 17601 27829 17635 27863
rect 19441 27829 19475 27863
rect 20177 27829 20211 27863
rect 24777 27829 24811 27863
rect 1856 27625 1890 27659
rect 5444 27625 5478 27659
rect 10885 27625 10919 27659
rect 4721 27557 4755 27591
rect 8585 27557 8619 27591
rect 20729 27557 20763 27591
rect 21649 27557 21683 27591
rect 22753 27557 22787 27591
rect 5181 27489 5215 27523
rect 9137 27489 9171 27523
rect 9413 27489 9447 27523
rect 11529 27489 11563 27523
rect 15025 27489 15059 27523
rect 16313 27489 16347 27523
rect 18429 27489 18463 27523
rect 20177 27489 20211 27523
rect 22569 27489 22603 27523
rect 1593 27421 1627 27455
rect 4077 27421 4111 27455
rect 4261 27421 4295 27455
rect 7205 27421 7239 27455
rect 7941 27421 7975 27455
rect 8125 27421 8159 27455
rect 14473 27421 14507 27455
rect 16129 27421 16163 27455
rect 17785 27421 17819 27455
rect 18245 27421 18279 27455
rect 19625 27421 19659 27455
rect 21281 27421 21315 27455
rect 21465 27421 21499 27455
rect 22385 27421 22419 27455
rect 23673 27421 23707 27455
rect 24593 27421 24627 27455
rect 31677 27421 31711 27455
rect 38025 27421 38059 27455
rect 11621 27353 11655 27387
rect 12173 27353 12207 27387
rect 12909 27353 12943 27387
rect 13001 27353 13035 27387
rect 13553 27353 13587 27387
rect 15117 27353 15151 27387
rect 15669 27353 15703 27387
rect 18889 27353 18923 27387
rect 20269 27353 20303 27387
rect 3341 27285 3375 27319
rect 14289 27285 14323 27319
rect 16773 27285 16807 27319
rect 17601 27285 17635 27319
rect 19441 27285 19475 27319
rect 23489 27285 23523 27319
rect 24685 27285 24719 27319
rect 31769 27285 31803 27319
rect 38209 27285 38243 27319
rect 1777 27081 1811 27115
rect 2789 27081 2823 27115
rect 5825 27081 5859 27115
rect 14841 27081 14875 27115
rect 18705 27081 18739 27115
rect 25145 27081 25179 27115
rect 29193 27081 29227 27115
rect 3617 27013 3651 27047
rect 5365 27013 5399 27047
rect 11805 27013 11839 27047
rect 11897 27013 11931 27047
rect 1593 26945 1627 26979
rect 2605 26945 2639 26979
rect 6009 26945 6043 26979
rect 7021 26945 7055 26979
rect 9229 26945 9263 26979
rect 13093 26945 13127 26979
rect 13553 26945 13587 26979
rect 14381 26945 14415 26979
rect 17417 26945 17451 26979
rect 19809 26945 19843 26979
rect 23121 26945 23155 26979
rect 24685 26945 24719 26979
rect 29101 26945 29135 26979
rect 32505 26945 32539 26979
rect 3341 26877 3375 26911
rect 7297 26877 7331 26911
rect 9505 26877 9539 26911
rect 14197 26877 14231 26911
rect 15669 26877 15703 26911
rect 15853 26877 15887 26911
rect 18061 26877 18095 26911
rect 18245 26877 18279 26911
rect 20269 26877 20303 26911
rect 20913 26877 20947 26911
rect 22017 26877 22051 26911
rect 22201 26877 22235 26911
rect 23305 26877 23339 26911
rect 24501 26877 24535 26911
rect 12357 26809 12391 26843
rect 16037 26809 16071 26843
rect 8769 26741 8803 26775
rect 10977 26741 11011 26775
rect 12909 26741 12943 26775
rect 13645 26741 13679 26775
rect 17509 26741 17543 26775
rect 19625 26741 19659 26775
rect 22385 26741 22419 26775
rect 23765 26741 23799 26775
rect 32597 26741 32631 26775
rect 1856 26537 1890 26571
rect 5733 26537 5767 26571
rect 7100 26537 7134 26571
rect 11621 26537 11655 26571
rect 15117 26537 15151 26571
rect 25881 26537 25915 26571
rect 34897 26537 34931 26571
rect 3341 26469 3375 26503
rect 6285 26469 6319 26503
rect 8585 26469 8619 26503
rect 12909 26469 12943 26503
rect 16773 26469 16807 26503
rect 17509 26469 17543 26503
rect 18153 26469 18187 26503
rect 3985 26401 4019 26435
rect 4261 26401 4295 26435
rect 6837 26401 6871 26435
rect 9505 26401 9539 26435
rect 10149 26401 10183 26435
rect 14657 26401 14691 26435
rect 16482 26401 16516 26435
rect 23397 26401 23431 26435
rect 23581 26401 23615 26435
rect 1593 26333 1627 26367
rect 6193 26333 6227 26367
rect 10977 26333 11011 26367
rect 11805 26333 11839 26367
rect 12265 26333 12299 26367
rect 13093 26333 13127 26367
rect 13737 26333 13771 26367
rect 14473 26333 14507 26367
rect 15669 26333 15703 26367
rect 16313 26333 16347 26367
rect 17693 26333 17727 26367
rect 18337 26333 18371 26367
rect 20821 26333 20855 26367
rect 22109 26333 22143 26367
rect 22569 26333 22603 26367
rect 24777 26333 24811 26367
rect 25421 26333 25455 26367
rect 26065 26333 26099 26367
rect 35081 26333 35115 26367
rect 9597 26265 9631 26299
rect 11069 26265 11103 26299
rect 15761 26265 15795 26299
rect 19533 26265 19567 26299
rect 19625 26265 19659 26299
rect 20177 26265 20211 26299
rect 24041 26265 24075 26299
rect 12357 26197 12391 26231
rect 13553 26197 13587 26231
rect 20637 26197 20671 26231
rect 21281 26197 21315 26231
rect 21925 26197 21959 26231
rect 22661 26197 22695 26231
rect 24593 26197 24627 26231
rect 25237 26197 25271 26231
rect 13185 25993 13219 26027
rect 15853 25993 15887 26027
rect 16957 25993 16991 26027
rect 18981 25993 19015 26027
rect 24409 25993 24443 26027
rect 4353 25925 4387 25959
rect 8493 25925 8527 25959
rect 20821 25925 20855 25959
rect 20913 25925 20947 25959
rect 21465 25925 21499 25959
rect 22753 25925 22787 25959
rect 23305 25925 23339 25959
rect 4077 25857 4111 25891
rect 8217 25857 8251 25891
rect 10977 25857 11011 25891
rect 12081 25857 12115 25891
rect 12725 25857 12759 25891
rect 14105 25857 14139 25891
rect 14565 25857 14599 25891
rect 15393 25857 15427 25891
rect 17141 25857 17175 25891
rect 17785 25857 17819 25891
rect 18429 25857 18463 25891
rect 19165 25857 19199 25891
rect 19625 25857 19659 25891
rect 23765 25857 23799 25891
rect 24593 25857 24627 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 34621 25857 34655 25891
rect 1593 25789 1627 25823
rect 1869 25789 1903 25823
rect 3617 25789 3651 25823
rect 5825 25789 5859 25823
rect 7113 25789 7147 25823
rect 7297 25789 7331 25823
rect 11069 25789 11103 25823
rect 12541 25789 12575 25823
rect 15209 25789 15243 25823
rect 19809 25789 19843 25823
rect 22661 25789 22695 25823
rect 25053 25789 25087 25823
rect 14657 25721 14691 25755
rect 17601 25721 17635 25755
rect 19993 25721 20027 25755
rect 7757 25653 7791 25687
rect 9965 25653 9999 25687
rect 11897 25653 11931 25687
rect 13921 25653 13955 25687
rect 18245 25653 18279 25687
rect 23857 25653 23891 25687
rect 34437 25653 34471 25687
rect 1856 25449 1890 25483
rect 3985 25449 4019 25483
rect 5549 25449 5583 25483
rect 6837 25449 6871 25483
rect 7481 25449 7515 25483
rect 12357 25449 12391 25483
rect 16589 25449 16623 25483
rect 17417 25449 17451 25483
rect 18613 25449 18647 25483
rect 20913 25449 20947 25483
rect 22293 25449 22327 25483
rect 23489 25449 23523 25483
rect 9321 25381 9355 25415
rect 10149 25381 10183 25415
rect 1593 25313 1627 25347
rect 8125 25313 8159 25347
rect 14657 25313 14691 25347
rect 16129 25313 16163 25347
rect 17233 25313 17267 25347
rect 18429 25313 18463 25347
rect 20269 25313 20303 25347
rect 20453 25313 20487 25347
rect 21833 25313 21867 25347
rect 23029 25313 23063 25347
rect 4169 25245 4203 25279
rect 4905 25245 4939 25279
rect 5733 25245 5767 25279
rect 6745 25245 6779 25279
rect 7389 25245 7423 25279
rect 8033 25245 8067 25279
rect 9505 25245 9539 25279
rect 10333 25245 10367 25279
rect 11253 25245 11287 25279
rect 11713 25245 11747 25279
rect 12541 25245 12575 25279
rect 15945 25245 15979 25279
rect 17049 25245 17083 25279
rect 18245 25245 18279 25279
rect 19625 25245 19659 25279
rect 21649 25245 21683 25279
rect 22845 25245 22879 25279
rect 24593 25245 24627 25279
rect 38025 25245 38059 25279
rect 13093 25177 13127 25211
rect 13185 25177 13219 25211
rect 13737 25177 13771 25211
rect 14381 25177 14415 25211
rect 14473 25177 14507 25211
rect 3341 25109 3375 25143
rect 4997 25109 5031 25143
rect 11069 25109 11103 25143
rect 11805 25109 11839 25143
rect 19441 25109 19475 25143
rect 24685 25109 24719 25143
rect 38209 25109 38243 25143
rect 13369 24905 13403 24939
rect 15301 24837 15335 24871
rect 23305 24837 23339 24871
rect 1777 24769 1811 24803
rect 2513 24769 2547 24803
rect 5089 24769 5123 24803
rect 5549 24769 5583 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 7665 24769 7699 24803
rect 8769 24769 8803 24803
rect 9413 24769 9447 24803
rect 9505 24769 9539 24803
rect 10517 24769 10551 24803
rect 11161 24769 11195 24803
rect 12081 24769 12115 24803
rect 12909 24769 12943 24803
rect 17325 24769 17359 24803
rect 18521 24769 18555 24803
rect 18705 24769 18739 24803
rect 19901 24769 19935 24803
rect 21189 24769 21223 24803
rect 22477 24769 22511 24803
rect 24501 24769 24535 24803
rect 24961 24769 24995 24803
rect 25789 24769 25823 24803
rect 27537 24769 27571 24803
rect 27629 24769 27663 24803
rect 2789 24701 2823 24735
rect 4261 24701 4295 24735
rect 5641 24701 5675 24735
rect 14013 24701 14047 24735
rect 14197 24701 14231 24735
rect 15209 24701 15243 24735
rect 15853 24701 15887 24735
rect 17509 24701 17543 24735
rect 20361 24701 20395 24735
rect 23213 24701 23247 24735
rect 4905 24633 4939 24667
rect 10333 24633 10367 24667
rect 10977 24633 11011 24667
rect 12173 24633 12207 24667
rect 12725 24633 12759 24667
rect 17693 24633 17727 24667
rect 18889 24633 18923 24667
rect 23765 24633 23799 24667
rect 1593 24565 1627 24599
rect 7757 24565 7791 24599
rect 8861 24565 8895 24599
rect 14381 24565 14415 24599
rect 19717 24565 19751 24599
rect 21005 24565 21039 24599
rect 22293 24565 22327 24599
rect 24317 24565 24351 24599
rect 25053 24565 25087 24599
rect 25605 24565 25639 24599
rect 2421 24361 2455 24395
rect 3065 24361 3099 24395
rect 4077 24361 4111 24395
rect 5733 24361 5767 24395
rect 6745 24361 6779 24395
rect 9965 24361 9999 24395
rect 11345 24361 11379 24395
rect 13001 24361 13035 24395
rect 14565 24361 14599 24395
rect 23673 24361 23707 24395
rect 24961 24361 24995 24395
rect 26341 24361 26375 24395
rect 16497 24293 16531 24327
rect 9781 24225 9815 24259
rect 11161 24225 11195 24259
rect 23213 24225 23247 24259
rect 24593 24225 24627 24259
rect 24777 24225 24811 24259
rect 1593 24157 1627 24191
rect 2329 24157 2363 24191
rect 2973 24157 3007 24191
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 5917 24157 5951 24191
rect 6929 24157 6963 24191
rect 7573 24157 7607 24191
rect 9597 24157 9631 24191
rect 10977 24157 11011 24191
rect 12265 24157 12299 24191
rect 12909 24157 12943 24191
rect 13737 24157 13771 24191
rect 14749 24157 14783 24191
rect 15209 24157 15243 24191
rect 17877 24157 17911 24191
rect 18061 24157 18095 24191
rect 19717 24157 19751 24191
rect 20545 24157 20579 24191
rect 21189 24157 21223 24191
rect 21833 24157 21867 24191
rect 23029 24157 23063 24191
rect 25881 24157 25915 24191
rect 26525 24157 26559 24191
rect 28825 24157 28859 24191
rect 38301 24157 38335 24191
rect 4721 24089 4755 24123
rect 15945 24089 15979 24123
rect 16037 24089 16071 24123
rect 1777 24021 1811 24055
rect 7665 24021 7699 24055
rect 12357 24021 12391 24055
rect 13553 24021 13587 24055
rect 15301 24021 15335 24055
rect 17233 24021 17267 24055
rect 18521 24021 18555 24055
rect 19809 24021 19843 24055
rect 20361 24021 20395 24055
rect 21005 24021 21039 24055
rect 21925 24021 21959 24055
rect 25697 24021 25731 24055
rect 28917 24021 28951 24055
rect 38117 24021 38151 24055
rect 2329 23817 2363 23851
rect 2973 23817 3007 23851
rect 8585 23817 8619 23851
rect 18429 23817 18463 23851
rect 20821 23817 20855 23851
rect 3617 23749 3651 23783
rect 8033 23749 8067 23783
rect 9413 23749 9447 23783
rect 9965 23749 9999 23783
rect 14841 23749 14875 23783
rect 22293 23749 22327 23783
rect 22845 23749 22879 23783
rect 25053 23749 25087 23783
rect 1593 23681 1627 23715
rect 2237 23681 2271 23715
rect 2881 23681 2915 23715
rect 3525 23681 3559 23715
rect 6745 23681 6779 23715
rect 7941 23681 7975 23715
rect 8769 23681 8803 23715
rect 11161 23681 11195 23715
rect 11713 23681 11747 23715
rect 11897 23681 11931 23715
rect 13553 23681 13587 23715
rect 14197 23681 14231 23715
rect 17325 23681 17359 23715
rect 17785 23681 17819 23715
rect 17969 23681 18003 23715
rect 19073 23681 19107 23715
rect 20361 23681 20395 23715
rect 21465 23681 21499 23715
rect 23305 23681 23339 23715
rect 23949 23681 23983 23715
rect 24593 23681 24627 23715
rect 6837 23613 6871 23647
rect 9321 23613 9355 23647
rect 14749 23613 14783 23647
rect 15301 23613 15335 23647
rect 18889 23613 18923 23647
rect 20177 23613 20211 23647
rect 22201 23613 22235 23647
rect 23489 23613 23523 23647
rect 1685 23545 1719 23579
rect 12173 23545 12207 23579
rect 24409 23545 24443 23579
rect 10977 23477 11011 23511
rect 13369 23477 13403 23511
rect 14013 23477 14047 23511
rect 17141 23477 17175 23511
rect 19257 23477 19291 23511
rect 21281 23477 21315 23511
rect 1593 23273 1627 23307
rect 2973 23273 3007 23307
rect 8401 23273 8435 23307
rect 11529 23273 11563 23307
rect 16313 23273 16347 23307
rect 24593 23273 24627 23307
rect 11989 23205 12023 23239
rect 13277 23205 13311 23239
rect 14749 23205 14783 23239
rect 15669 23205 15703 23239
rect 18889 23205 18923 23239
rect 20269 23205 20303 23239
rect 9413 23137 9447 23171
rect 9597 23137 9631 23171
rect 10885 23137 10919 23171
rect 12817 23137 12851 23171
rect 14565 23137 14599 23171
rect 17601 23137 17635 23171
rect 18245 23137 18279 23171
rect 20085 23137 20119 23171
rect 21005 23137 21039 23171
rect 22845 23137 22879 23171
rect 23397 23137 23431 23171
rect 23857 23137 23891 23171
rect 1777 23069 1811 23103
rect 2237 23069 2271 23103
rect 2881 23069 2915 23103
rect 7113 23069 7147 23103
rect 8585 23069 8619 23103
rect 11069 23069 11103 23103
rect 12173 23069 12207 23103
rect 12633 23069 12667 23103
rect 14381 23069 14415 23103
rect 15577 23069 15611 23103
rect 16221 23069 16255 23103
rect 18429 23069 18463 23103
rect 19901 23069 19935 23103
rect 21189 23069 21223 23103
rect 24777 23069 24811 23103
rect 2329 23001 2363 23035
rect 7205 23001 7239 23035
rect 16957 23001 16991 23035
rect 17049 23001 17083 23035
rect 22201 23001 22235 23035
rect 22293 23001 22327 23035
rect 23489 23001 23523 23035
rect 7757 22933 7791 22967
rect 10057 22933 10091 22967
rect 21649 22933 21683 22967
rect 1593 22729 1627 22763
rect 8493 22729 8527 22763
rect 13093 22729 13127 22763
rect 13737 22729 13771 22763
rect 17693 22729 17727 22763
rect 22109 22729 22143 22763
rect 23949 22729 23983 22763
rect 17141 22661 17175 22695
rect 18521 22661 18555 22695
rect 19625 22661 19659 22695
rect 19717 22661 19751 22695
rect 20913 22661 20947 22695
rect 21465 22661 21499 22695
rect 1777 22593 1811 22627
rect 7389 22593 7423 22627
rect 8401 22593 8435 22627
rect 9689 22593 9723 22627
rect 10517 22593 10551 22627
rect 11161 22593 11195 22627
rect 11897 22593 11931 22627
rect 13277 22593 13311 22627
rect 14565 22593 14599 22627
rect 15485 22593 15519 22627
rect 16313 22593 16347 22627
rect 17049 22593 17083 22627
rect 17877 22593 17911 22627
rect 22017 22593 22051 22627
rect 24593 22593 24627 22627
rect 25053 22593 25087 22627
rect 30297 22593 30331 22627
rect 34989 22593 35023 22627
rect 9045 22525 9079 22559
rect 9781 22525 9815 22559
rect 11711 22525 11745 22559
rect 12357 22525 12391 22559
rect 14381 22525 14415 22559
rect 18429 22525 18463 22559
rect 19901 22525 19935 22559
rect 20821 22525 20855 22559
rect 22661 22525 22695 22559
rect 23305 22525 23339 22559
rect 23489 22525 23523 22559
rect 25145 22525 25179 22559
rect 10333 22457 10367 22491
rect 14749 22457 14783 22491
rect 15577 22457 15611 22491
rect 18981 22457 19015 22491
rect 24409 22457 24443 22491
rect 7205 22389 7239 22423
rect 10977 22389 11011 22423
rect 16129 22389 16163 22423
rect 30389 22389 30423 22423
rect 34805 22389 34839 22423
rect 7389 22117 7423 22151
rect 10701 22117 10735 22151
rect 12357 22117 12391 22151
rect 18521 22117 18555 22151
rect 19809 22117 19843 22151
rect 8125 22049 8159 22083
rect 9137 22049 9171 22083
rect 9321 22049 9355 22083
rect 9781 22049 9815 22083
rect 11989 22049 12023 22083
rect 13093 22049 13127 22083
rect 14933 22049 14967 22083
rect 16773 22049 16807 22083
rect 17417 22049 17451 22083
rect 19441 22049 19475 22083
rect 20821 22049 20855 22083
rect 21557 22049 21591 22083
rect 31309 22049 31343 22083
rect 6653 21981 6687 22015
rect 7297 21981 7331 22015
rect 7941 21981 7975 22015
rect 10885 21981 10919 22015
rect 11345 21981 11379 22015
rect 12173 21981 12207 22015
rect 13277 21981 13311 22015
rect 16221 21981 16255 22015
rect 19625 21981 19659 22015
rect 20729 21981 20763 22015
rect 21373 21981 21407 22015
rect 31217 21981 31251 22015
rect 38301 21981 38335 22015
rect 11437 21913 11471 21947
rect 15025 21913 15059 21947
rect 15577 21913 15611 21947
rect 16865 21913 16899 21947
rect 17969 21913 18003 21947
rect 18061 21913 18095 21947
rect 22017 21913 22051 21947
rect 23029 21913 23063 21947
rect 23121 21913 23155 21947
rect 23673 21913 23707 21947
rect 6745 21845 6779 21879
rect 8585 21845 8619 21879
rect 13737 21845 13771 21879
rect 16037 21845 16071 21879
rect 38117 21845 38151 21879
rect 8401 21641 8435 21675
rect 9689 21641 9723 21675
rect 17141 21641 17175 21675
rect 18429 21641 18463 21675
rect 21465 21641 21499 21675
rect 22661 21641 22695 21675
rect 14565 21573 14599 21607
rect 7757 21505 7791 21539
rect 8585 21505 8619 21539
rect 10517 21505 10551 21539
rect 10977 21505 11011 21539
rect 11713 21505 11747 21539
rect 16313 21505 16347 21539
rect 17325 21505 17359 21539
rect 17785 21505 17819 21539
rect 19073 21505 19107 21539
rect 19533 21505 19567 21539
rect 22017 21505 22051 21539
rect 23305 21505 23339 21539
rect 23949 21505 23983 21539
rect 7113 21437 7147 21471
rect 9045 21437 9079 21471
rect 9229 21437 9263 21471
rect 11897 21437 11931 21471
rect 13001 21437 13035 21471
rect 13185 21437 13219 21471
rect 14473 21437 14507 21471
rect 17969 21437 18003 21471
rect 19717 21437 19751 21471
rect 20821 21437 20855 21471
rect 21005 21437 21039 21471
rect 22201 21437 22235 21471
rect 7849 21369 7883 21403
rect 10333 21369 10367 21403
rect 13369 21369 13403 21403
rect 15025 21369 15059 21403
rect 16129 21369 16163 21403
rect 18889 21369 18923 21403
rect 23121 21369 23155 21403
rect 11069 21301 11103 21335
rect 12357 21301 12391 21335
rect 20177 21301 20211 21335
rect 23765 21301 23799 21335
rect 1593 21097 1627 21131
rect 6561 21097 6595 21131
rect 10793 21097 10827 21131
rect 11713 21097 11747 21131
rect 16589 21097 16623 21131
rect 18061 21097 18095 21131
rect 22937 21097 22971 21131
rect 14289 21029 14323 21063
rect 19901 21029 19935 21063
rect 10149 20961 10183 20995
rect 10333 20961 10367 20995
rect 13461 20961 13495 20995
rect 16221 20961 16255 20995
rect 16405 20961 16439 20995
rect 21189 20961 21223 20995
rect 21833 20961 21867 20995
rect 1777 20893 1811 20927
rect 6469 20893 6503 20927
rect 7297 20893 7331 20927
rect 8585 20893 8619 20927
rect 9689 20893 9723 20927
rect 11897 20893 11931 20927
rect 12541 20893 12575 20927
rect 14473 20893 14507 20927
rect 14933 20893 14967 20927
rect 15761 20893 15795 20927
rect 17693 20893 17727 20927
rect 17877 20893 17911 20927
rect 20085 20893 20119 20927
rect 20545 20893 20579 20927
rect 20729 20893 20763 20927
rect 22477 20893 22511 20927
rect 23121 20893 23155 20927
rect 23765 20893 23799 20927
rect 24777 20893 24811 20927
rect 38025 20893 38059 20927
rect 7757 20825 7791 20859
rect 13093 20825 13127 20859
rect 13185 20825 13219 20859
rect 15025 20825 15059 20859
rect 21925 20825 21959 20859
rect 7113 20757 7147 20791
rect 8401 20757 8435 20791
rect 9505 20757 9539 20791
rect 12357 20757 12391 20791
rect 15577 20757 15611 20791
rect 23581 20757 23615 20791
rect 24593 20757 24627 20791
rect 38209 20757 38243 20791
rect 5273 20553 5307 20587
rect 7757 20553 7791 20587
rect 9045 20553 9079 20587
rect 16865 20553 16899 20587
rect 22017 20553 22051 20587
rect 25053 20553 25087 20587
rect 7205 20485 7239 20519
rect 11805 20485 11839 20519
rect 11897 20485 11931 20519
rect 18981 20485 19015 20519
rect 20361 20485 20395 20519
rect 22845 20485 22879 20519
rect 24041 20485 24075 20519
rect 5181 20417 5215 20451
rect 6009 20417 6043 20451
rect 7113 20417 7147 20451
rect 7941 20417 7975 20451
rect 8585 20417 8619 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 14473 20417 14507 20451
rect 15577 20417 15611 20451
rect 17049 20417 17083 20451
rect 18337 20417 18371 20451
rect 25237 20417 25271 20451
rect 10977 20349 11011 20383
rect 13185 20349 13219 20383
rect 13369 20349 13403 20383
rect 14289 20349 14323 20383
rect 15393 20349 15427 20383
rect 17509 20349 17543 20383
rect 18889 20349 18923 20383
rect 20269 20349 20303 20383
rect 22753 20349 22787 20383
rect 23949 20349 23983 20383
rect 9689 20281 9723 20315
rect 12357 20281 12391 20315
rect 18153 20281 18187 20315
rect 19441 20281 19475 20315
rect 20821 20281 20855 20315
rect 23305 20281 23339 20315
rect 24501 20281 24535 20315
rect 5825 20213 5859 20247
rect 8401 20213 8435 20247
rect 10333 20213 10367 20247
rect 13829 20213 13863 20247
rect 14657 20213 14691 20247
rect 15761 20213 15795 20247
rect 5917 20009 5951 20043
rect 15301 20009 15335 20043
rect 16773 20009 16807 20043
rect 18797 20009 18831 20043
rect 20545 20009 20579 20043
rect 21557 20009 21591 20043
rect 22477 20009 22511 20043
rect 24685 20009 24719 20043
rect 13461 19941 13495 19975
rect 14381 19941 14415 19975
rect 17877 19941 17911 19975
rect 23581 19941 23615 19975
rect 7941 19873 7975 19907
rect 9137 19873 9171 19907
rect 10517 19873 10551 19907
rect 15117 19873 15151 19907
rect 16129 19873 16163 19907
rect 17417 19873 17451 19907
rect 21005 19873 21039 19907
rect 22109 19873 22143 19907
rect 5825 19805 5859 19839
rect 6653 19805 6687 19839
rect 7297 19805 7331 19839
rect 7757 19805 7791 19839
rect 9965 19805 9999 19839
rect 12357 19805 12391 19839
rect 14289 19805 14323 19839
rect 14933 19805 14967 19839
rect 16313 19805 16347 19839
rect 17233 19805 17267 19839
rect 18705 19805 18739 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 21189 19805 21223 19839
rect 22293 19805 22327 19839
rect 23213 19805 23247 19839
rect 23397 19805 23431 19839
rect 24593 19805 24627 19839
rect 10609 19737 10643 19771
rect 11161 19737 11195 19771
rect 12909 19737 12943 19771
rect 13001 19737 13035 19771
rect 6469 19669 6503 19703
rect 7113 19669 7147 19703
rect 8401 19669 8435 19703
rect 9781 19669 9815 19703
rect 12173 19669 12207 19703
rect 1593 19465 1627 19499
rect 7113 19465 7147 19499
rect 7757 19465 7791 19499
rect 9045 19465 9079 19499
rect 9781 19465 9815 19499
rect 16129 19465 16163 19499
rect 18245 19465 18279 19499
rect 18889 19465 18923 19499
rect 19533 19465 19567 19499
rect 20177 19465 20211 19499
rect 20821 19465 20855 19499
rect 22753 19465 22787 19499
rect 23213 19465 23247 19499
rect 23857 19465 23891 19499
rect 12081 19397 12115 19431
rect 14289 19397 14323 19431
rect 14381 19397 14415 19431
rect 1777 19329 1811 19363
rect 7297 19329 7331 19363
rect 7941 19329 7975 19363
rect 8585 19329 8619 19363
rect 9229 19329 9263 19363
rect 9689 19329 9723 19363
rect 10517 19329 10551 19363
rect 10977 19329 11011 19363
rect 13737 19329 13771 19363
rect 16313 19329 16347 19363
rect 17601 19329 17635 19363
rect 18429 19329 18463 19363
rect 19073 19329 19107 19363
rect 19717 19329 19751 19363
rect 21005 19329 21039 19363
rect 22109 19329 22143 19363
rect 23397 19329 23431 19363
rect 28825 19329 28859 19363
rect 28917 19329 28951 19363
rect 11989 19261 12023 19295
rect 12265 19261 12299 19295
rect 15117 19261 15151 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 22293 19261 22327 19295
rect 10333 19193 10367 19227
rect 11069 19193 11103 19227
rect 8401 19125 8435 19159
rect 13553 19125 13587 19159
rect 10517 18921 10551 18955
rect 21557 18921 21591 18955
rect 22937 18921 22971 18955
rect 23489 18921 23523 18955
rect 8401 18853 8435 18887
rect 9873 18853 9907 18887
rect 13461 18853 13495 18887
rect 21005 18853 21039 18887
rect 13277 18785 13311 18819
rect 14381 18785 14415 18819
rect 15393 18785 15427 18819
rect 18245 18785 18279 18819
rect 7113 18717 7147 18751
rect 7941 18717 7975 18751
rect 8585 18717 8619 18751
rect 9413 18717 9447 18751
rect 10057 18717 10091 18751
rect 10701 18717 10735 18751
rect 12449 18717 12483 18751
rect 13093 18717 13127 18751
rect 16221 18717 16255 18751
rect 16405 18717 16439 18751
rect 20913 18717 20947 18751
rect 21741 18717 21775 18751
rect 22201 18717 22235 18751
rect 22845 18717 22879 18751
rect 23673 18717 23707 18751
rect 29745 18717 29779 18751
rect 35081 18717 35115 18751
rect 7205 18649 7239 18683
rect 11253 18649 11287 18683
rect 11345 18649 11379 18683
rect 11897 18649 11931 18683
rect 14473 18649 14507 18683
rect 17417 18649 17451 18683
rect 17509 18649 17543 18683
rect 19533 18649 19567 18683
rect 19625 18649 19659 18683
rect 20177 18649 20211 18683
rect 7757 18581 7791 18615
rect 9229 18581 9263 18615
rect 12541 18581 12575 18615
rect 16865 18581 16899 18615
rect 22293 18581 22327 18615
rect 29837 18581 29871 18615
rect 34897 18581 34931 18615
rect 1593 18377 1627 18411
rect 9229 18377 9263 18411
rect 9873 18377 9907 18411
rect 16313 18377 16347 18411
rect 18613 18377 18647 18411
rect 11805 18309 11839 18343
rect 11897 18309 11931 18343
rect 17049 18309 17083 18343
rect 17601 18309 17635 18343
rect 20545 18309 20579 18343
rect 22201 18309 22235 18343
rect 1777 18241 1811 18275
rect 5917 18241 5951 18275
rect 7481 18241 7515 18275
rect 8125 18241 8159 18275
rect 8769 18241 8803 18275
rect 9413 18241 9447 18275
rect 10057 18241 10091 18275
rect 12909 18241 12943 18275
rect 14565 18241 14599 18275
rect 15853 18241 15887 18275
rect 19257 18241 19291 18275
rect 10517 18173 10551 18207
rect 10701 18173 10735 18207
rect 12081 18173 12115 18207
rect 13093 18173 13127 18207
rect 14749 18173 14783 18207
rect 15669 18173 15703 18207
rect 16957 18173 16991 18207
rect 19441 18173 19475 18207
rect 19901 18173 19935 18207
rect 20453 18173 20487 18207
rect 21465 18173 21499 18207
rect 22109 18173 22143 18207
rect 23121 18173 23155 18207
rect 7941 18105 7975 18139
rect 13277 18105 13311 18139
rect 5733 18037 5767 18071
rect 7297 18037 7331 18071
rect 8585 18037 8619 18071
rect 11161 18037 11195 18071
rect 15209 18037 15243 18071
rect 18061 17833 18095 17867
rect 20269 17833 20303 17867
rect 22661 17833 22695 17867
rect 11069 17765 11103 17799
rect 21557 17765 21591 17799
rect 8493 17697 8527 17731
rect 9505 17697 9539 17731
rect 11713 17697 11747 17731
rect 14749 17697 14783 17731
rect 16497 17697 16531 17731
rect 18797 17697 18831 17731
rect 19993 17697 20027 17731
rect 20913 17697 20947 17731
rect 22017 17697 22051 17731
rect 7941 17629 7975 17663
rect 8401 17629 8435 17663
rect 9321 17629 9355 17663
rect 10425 17629 10459 17663
rect 10609 17629 10643 17663
rect 11529 17629 11563 17663
rect 18245 17629 18279 17663
rect 18705 17629 18739 17663
rect 19809 17629 19843 17663
rect 21097 17629 21131 17663
rect 22845 17629 22879 17663
rect 27813 17629 27847 17663
rect 9965 17561 9999 17595
rect 12725 17561 12759 17595
rect 12817 17561 12851 17595
rect 13369 17561 13403 17595
rect 14841 17561 14875 17595
rect 15393 17561 15427 17595
rect 16589 17561 16623 17595
rect 17141 17561 17175 17595
rect 7757 17493 7791 17527
rect 12173 17493 12207 17527
rect 27905 17493 27939 17527
rect 11069 17289 11103 17323
rect 14013 17289 14047 17323
rect 16129 17289 16163 17323
rect 20545 17289 20579 17323
rect 22017 17289 22051 17323
rect 10425 17221 10459 17255
rect 12909 17221 12943 17255
rect 15393 17221 15427 17255
rect 18337 17221 18371 17255
rect 21189 17221 21223 17255
rect 8493 17153 8527 17187
rect 8953 17153 8987 17187
rect 9873 17153 9907 17187
rect 10333 17153 10367 17187
rect 10977 17153 11011 17187
rect 13553 17153 13587 17187
rect 19349 17153 19383 17187
rect 20453 17153 20487 17187
rect 21097 17153 21131 17187
rect 22201 17153 22235 17187
rect 38025 17153 38059 17187
rect 8309 17085 8343 17119
rect 12265 17085 12299 17119
rect 12449 17085 12483 17119
rect 13369 17085 13403 17119
rect 14749 17085 14783 17119
rect 14933 17085 14967 17119
rect 17049 17085 17083 17119
rect 17233 17085 17267 17119
rect 18245 17085 18279 17119
rect 19533 17085 19567 17119
rect 9689 17017 9723 17051
rect 18797 17017 18831 17051
rect 19993 17017 20027 17051
rect 38209 17017 38243 17051
rect 17417 16949 17451 16983
rect 17877 16745 17911 16779
rect 18613 16745 18647 16779
rect 20085 16745 20119 16779
rect 11253 16609 11287 16643
rect 14473 16609 14507 16643
rect 14657 16609 14691 16643
rect 15853 16609 15887 16643
rect 16497 16609 16531 16643
rect 17509 16609 17543 16643
rect 17693 16609 17727 16643
rect 9505 16541 9539 16575
rect 9965 16541 9999 16575
rect 10609 16541 10643 16575
rect 10701 16541 10735 16575
rect 11437 16541 11471 16575
rect 13093 16541 13127 16575
rect 13553 16541 13587 16575
rect 18797 16541 18831 16575
rect 19625 16541 19659 16575
rect 20269 16541 20303 16575
rect 20913 16541 20947 16575
rect 27169 16541 27203 16575
rect 33609 16541 33643 16575
rect 10057 16473 10091 16507
rect 15945 16473 15979 16507
rect 9321 16405 9355 16439
rect 11897 16405 11931 16439
rect 12909 16405 12943 16439
rect 15117 16405 15151 16439
rect 19441 16405 19475 16439
rect 20729 16405 20763 16439
rect 27261 16405 27295 16439
rect 33701 16405 33735 16439
rect 8953 16201 8987 16235
rect 10425 16201 10459 16235
rect 10977 16201 11011 16235
rect 13553 16201 13587 16235
rect 17693 16201 17727 16235
rect 18337 16201 18371 16235
rect 18981 16201 19015 16235
rect 38117 16201 38151 16235
rect 14105 16133 14139 16167
rect 14197 16133 14231 16167
rect 15577 16133 15611 16167
rect 19625 16133 19659 16167
rect 1593 16065 1627 16099
rect 8861 16065 8895 16099
rect 9505 16065 9539 16099
rect 10333 16065 10367 16099
rect 11161 16065 11195 16099
rect 11989 16065 12023 16099
rect 12449 16065 12483 16099
rect 17049 16065 17083 16099
rect 17877 16065 17911 16099
rect 18521 16065 18555 16099
rect 20453 16065 20487 16099
rect 31585 16065 31619 16099
rect 33609 16065 33643 16099
rect 38301 16065 38335 16099
rect 12909 15997 12943 16031
rect 13093 15997 13127 16031
rect 15485 15997 15519 16031
rect 16129 15997 16163 16031
rect 14657 15929 14691 15963
rect 1777 15861 1811 15895
rect 9597 15861 9631 15895
rect 12265 15861 12299 15895
rect 16865 15861 16899 15895
rect 20269 15861 20303 15895
rect 31677 15861 31711 15895
rect 33425 15861 33459 15895
rect 9781 15657 9815 15691
rect 10425 15657 10459 15691
rect 11713 15657 11747 15691
rect 12265 15657 12299 15691
rect 13645 15657 13679 15691
rect 14565 15657 14599 15691
rect 18429 15657 18463 15691
rect 19441 15589 19475 15623
rect 9321 15521 9355 15555
rect 12909 15521 12943 15555
rect 15117 15521 15151 15555
rect 17325 15521 17359 15555
rect 17509 15521 17543 15555
rect 9137 15453 9171 15487
rect 10609 15453 10643 15487
rect 11621 15453 11655 15487
rect 12449 15453 12483 15487
rect 13553 15453 13587 15487
rect 14473 15453 14507 15487
rect 15301 15453 15335 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 18613 15453 18647 15487
rect 19625 15453 19659 15487
rect 35081 15453 35115 15487
rect 17969 15385 18003 15419
rect 15761 15317 15795 15351
rect 16865 15317 16899 15351
rect 34897 15317 34931 15351
rect 7021 15113 7055 15147
rect 7665 15113 7699 15147
rect 12909 15113 12943 15147
rect 13553 15113 13587 15147
rect 14289 15113 14323 15147
rect 16129 15113 16163 15147
rect 17969 15113 18003 15147
rect 12357 15045 12391 15079
rect 6929 14977 6963 15011
rect 7573 14977 7607 15011
rect 12265 14977 12299 15011
rect 13093 14977 13127 15011
rect 13737 14977 13771 15011
rect 14197 14977 14231 15011
rect 15025 14977 15059 15011
rect 15669 14977 15703 15011
rect 16313 14977 16347 15011
rect 18613 14977 18647 15011
rect 17325 14909 17359 14943
rect 17509 14909 17543 14943
rect 14841 14841 14875 14875
rect 15485 14841 15519 14875
rect 18429 14773 18463 14807
rect 1593 14569 1627 14603
rect 13553 14569 13587 14603
rect 14933 14569 14967 14603
rect 15485 14569 15519 14603
rect 16313 14569 16347 14603
rect 17325 14569 17359 14603
rect 17877 14569 17911 14603
rect 1777 14365 1811 14399
rect 13737 14365 13771 14399
rect 14841 14365 14875 14399
rect 15669 14365 15703 14399
rect 16221 14365 16255 14399
rect 17233 14365 17267 14399
rect 18061 14365 18095 14399
rect 35081 14365 35115 14399
rect 38025 14365 38059 14399
rect 34897 14229 34931 14263
rect 38209 14229 38243 14263
rect 14565 14025 14599 14059
rect 15301 14025 15335 14059
rect 15945 14025 15979 14059
rect 17141 14025 17175 14059
rect 15485 13889 15519 13923
rect 17049 13889 17083 13923
rect 8033 13481 8067 13515
rect 16129 13481 16163 13515
rect 7941 13277 7975 13311
rect 16037 13277 16071 13311
rect 1593 12937 1627 12971
rect 1777 12801 1811 12835
rect 7941 12801 7975 12835
rect 18613 12801 18647 12835
rect 23673 12801 23707 12835
rect 35541 12801 35575 12835
rect 38025 12801 38059 12835
rect 8033 12597 8067 12631
rect 18705 12597 18739 12631
rect 23765 12597 23799 12631
rect 35357 12597 35391 12631
rect 38209 12597 38243 12631
rect 6469 12393 6503 12427
rect 6377 12189 6411 12223
rect 17141 12189 17175 12223
rect 33425 12189 33459 12223
rect 17233 12053 17267 12087
rect 33517 12053 33551 12087
rect 32321 11713 32355 11747
rect 32413 11509 32447 11543
rect 1593 11305 1627 11339
rect 38209 11237 38243 11271
rect 1777 11101 1811 11135
rect 19441 11101 19475 11135
rect 38025 11101 38059 11135
rect 19533 11033 19567 11067
rect 11713 10625 11747 10659
rect 16037 10625 16071 10659
rect 18153 10625 18187 10659
rect 23581 10625 23615 10659
rect 26433 10625 26467 10659
rect 11805 10421 11839 10455
rect 16129 10421 16163 10455
rect 18245 10421 18279 10455
rect 23673 10421 23707 10455
rect 26525 10421 26559 10455
rect 1593 10217 1627 10251
rect 1777 10013 1811 10047
rect 4169 10013 4203 10047
rect 10701 10013 10735 10047
rect 3985 9877 4019 9911
rect 10793 9877 10827 9911
rect 13277 9129 13311 9163
rect 18245 9129 18279 9163
rect 13185 8925 13219 8959
rect 18153 8925 18187 8959
rect 38025 8925 38059 8959
rect 38209 8789 38243 8823
rect 11805 8585 11839 8619
rect 19349 8585 19383 8619
rect 22385 8585 22419 8619
rect 9597 8517 9631 8551
rect 9505 8449 9539 8483
rect 11713 8449 11747 8483
rect 19257 8449 19291 8483
rect 22385 8449 22419 8483
rect 1593 8041 1627 8075
rect 13553 8041 13587 8075
rect 26985 8041 27019 8075
rect 38117 8041 38151 8075
rect 1777 7837 1811 7871
rect 9137 7837 9171 7871
rect 13461 7837 13495 7871
rect 26893 7837 26927 7871
rect 35265 7837 35299 7871
rect 38301 7837 38335 7871
rect 9229 7769 9263 7803
rect 35357 7701 35391 7735
rect 34253 7361 34287 7395
rect 34345 7157 34379 7191
rect 24777 6953 24811 6987
rect 24685 6749 24719 6783
rect 11805 6409 11839 6443
rect 28917 6409 28951 6443
rect 8769 6341 8803 6375
rect 1593 6273 1627 6307
rect 8677 6273 8711 6307
rect 11713 6273 11747 6307
rect 28825 6273 28859 6307
rect 38117 6273 38151 6307
rect 1777 6137 1811 6171
rect 38209 6069 38243 6103
rect 6469 5865 6503 5899
rect 32781 5729 32815 5763
rect 4721 5661 4755 5695
rect 6377 5661 6411 5695
rect 9689 5661 9723 5695
rect 18337 5661 18371 5695
rect 21189 5661 21223 5695
rect 24777 5661 24811 5695
rect 30389 5661 30423 5695
rect 32689 5661 32723 5695
rect 37105 5661 37139 5695
rect 30481 5593 30515 5627
rect 4813 5525 4847 5559
rect 9505 5525 9539 5559
rect 18153 5525 18187 5559
rect 21005 5525 21039 5559
rect 24593 5525 24627 5559
rect 36921 5525 36955 5559
rect 1869 5253 1903 5287
rect 1685 5185 1719 5219
rect 5641 5185 5675 5219
rect 11897 5185 11931 5219
rect 15301 5185 15335 5219
rect 17785 5185 17819 5219
rect 20269 5185 20303 5219
rect 27905 5185 27939 5219
rect 5733 4981 5767 5015
rect 11713 4981 11747 5015
rect 15117 4981 15151 5015
rect 17601 4981 17635 5015
rect 20085 4981 20119 5015
rect 27721 4981 27755 5015
rect 38117 4777 38151 4811
rect 31677 4573 31711 4607
rect 38301 4573 38335 4607
rect 31493 4437 31527 4471
rect 3341 4097 3375 4131
rect 35817 4097 35851 4131
rect 3157 3893 3191 3927
rect 35909 3893 35943 3927
rect 1593 3689 1627 3723
rect 38117 3689 38151 3723
rect 1777 3485 1811 3519
rect 37473 3485 37507 3519
rect 38301 3485 38335 3519
rect 37289 3349 37323 3383
rect 2329 3145 2363 3179
rect 3065 3145 3099 3179
rect 36737 3145 36771 3179
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3249 3009 3283 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 1777 2805 1811 2839
rect 38209 2805 38243 2839
rect 2697 2601 2731 2635
rect 7205 2601 7239 2635
rect 10425 2601 10459 2635
rect 14289 2601 14323 2635
rect 18153 2601 18187 2635
rect 22017 2601 22051 2635
rect 27169 2601 27203 2635
rect 30389 2601 30423 2635
rect 34897 2601 34931 2635
rect 4629 2533 4663 2567
rect 29745 2533 29779 2567
rect 33609 2533 33643 2567
rect 1593 2397 1627 2431
rect 2881 2397 2915 2431
rect 4813 2397 4847 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 11713 2397 11747 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 16865 2397 16899 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 27353 2397 27387 2431
rect 29929 2397 29963 2431
rect 30573 2397 30607 2431
rect 32321 2397 32355 2431
rect 33793 2397 33827 2431
rect 35081 2397 35115 2431
rect 36185 2397 36219 2431
rect 38025 2397 38059 2431
rect 1777 2261 1811 2295
rect 6561 2261 6595 2295
rect 9321 2261 9355 2295
rect 11897 2261 11931 2295
rect 15117 2261 15151 2295
rect 17049 2261 17083 2295
rect 19625 2261 19659 2295
rect 22845 2261 22879 2295
rect 24777 2261 24811 2295
rect 26065 2261 26099 2295
rect 32505 2261 32539 2295
rect 36369 2261 36403 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 5902 37748 5908 37800
rect 5960 37788 5966 37800
rect 11054 37788 11060 37800
rect 5960 37760 11060 37788
rect 5960 37748 5966 37760
rect 11054 37748 11060 37760
rect 11112 37748 11118 37800
rect 4522 37680 4528 37732
rect 4580 37720 4586 37732
rect 6546 37720 6552 37732
rect 4580 37692 6552 37720
rect 4580 37680 4586 37692
rect 6546 37680 6552 37692
rect 6604 37680 6610 37732
rect 7006 37680 7012 37732
rect 7064 37720 7070 37732
rect 13262 37720 13268 37732
rect 7064 37692 13268 37720
rect 7064 37680 7070 37692
rect 13262 37680 13268 37692
rect 13320 37680 13326 37732
rect 4062 37612 4068 37664
rect 4120 37652 4126 37664
rect 19334 37652 19340 37664
rect 4120 37624 19340 37652
rect 4120 37612 4126 37624
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 4236 37451 4294 37457
rect 4236 37417 4248 37451
rect 4282 37448 4294 37451
rect 5902 37448 5908 37460
rect 4282 37420 5908 37448
rect 4282 37417 4294 37420
rect 4236 37411 4294 37417
rect 5902 37408 5908 37420
rect 5960 37408 5966 37460
rect 5994 37408 6000 37460
rect 6052 37448 6058 37460
rect 11054 37448 11060 37460
rect 6052 37420 10824 37448
rect 10967 37420 11060 37448
rect 6052 37408 6058 37420
rect 1857 37315 1915 37321
rect 1857 37281 1869 37315
rect 1903 37312 1915 37315
rect 4706 37312 4712 37324
rect 1903 37284 4712 37312
rect 1903 37281 1915 37284
rect 1857 37275 1915 37281
rect 4706 37272 4712 37284
rect 4764 37272 4770 37324
rect 7006 37312 7012 37324
rect 6967 37284 7012 37312
rect 7006 37272 7012 37284
rect 7064 37272 7070 37324
rect 9585 37315 9643 37321
rect 9585 37281 9597 37315
rect 9631 37312 9643 37315
rect 9950 37312 9956 37324
rect 9631 37284 9956 37312
rect 9631 37281 9643 37284
rect 9585 37275 9643 37281
rect 9950 37272 9956 37284
rect 10008 37272 10014 37324
rect 10796 37312 10824 37420
rect 11054 37408 11060 37420
rect 11112 37448 11118 37460
rect 13906 37448 13912 37460
rect 11112 37420 13912 37448
rect 11112 37408 11118 37420
rect 13906 37408 13912 37420
rect 13964 37408 13970 37460
rect 11977 37315 12035 37321
rect 11977 37312 11989 37315
rect 10796 37284 11989 37312
rect 11977 37281 11989 37284
rect 12023 37281 12035 37315
rect 11977 37275 12035 37281
rect 14200 37284 15884 37312
rect 14 37204 20 37256
rect 72 37244 78 37256
rect 1578 37244 1584 37256
rect 72 37216 1584 37244
rect 72 37204 78 37216
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 3970 37244 3976 37256
rect 3252 37216 3976 37244
rect 3142 37176 3148 37188
rect 3082 37148 3148 37176
rect 3142 37136 3148 37148
rect 3200 37136 3206 37188
rect 1578 37068 1584 37120
rect 1636 37108 1642 37120
rect 3252 37108 3280 37216
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 6730 37244 6736 37256
rect 6691 37216 6736 37244
rect 6730 37204 6736 37216
rect 6788 37204 6794 37256
rect 9122 37204 9128 37256
rect 9180 37244 9186 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 9180 37216 9321 37244
rect 9180 37204 9186 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 11054 37204 11060 37256
rect 11112 37244 11118 37256
rect 11701 37247 11759 37253
rect 11701 37244 11713 37247
rect 11112 37216 11713 37244
rect 11112 37204 11118 37216
rect 11701 37213 11713 37216
rect 11747 37213 11759 37247
rect 14200 37244 14228 37284
rect 13110 37216 14228 37244
rect 14277 37247 14335 37253
rect 11701 37207 11759 37213
rect 14277 37213 14289 37247
rect 14323 37244 14335 37247
rect 15102 37244 15108 37256
rect 14323 37216 15108 37244
rect 14323 37213 14335 37216
rect 14277 37207 14335 37213
rect 15102 37204 15108 37216
rect 15160 37204 15166 37256
rect 15565 37247 15623 37253
rect 15565 37213 15577 37247
rect 15611 37244 15623 37247
rect 15746 37244 15752 37256
rect 15611 37216 15752 37244
rect 15611 37213 15623 37216
rect 15565 37207 15623 37213
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 15856 37244 15884 37284
rect 16666 37244 16672 37256
rect 15856 37216 16672 37244
rect 16666 37204 16672 37216
rect 16724 37204 16730 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19300 37216 19625 37244
rect 19300 37204 19306 37216
rect 19613 37213 19625 37216
rect 19659 37244 19671 37247
rect 19889 37247 19947 37253
rect 19889 37244 19901 37247
rect 19659 37216 19901 37244
rect 19659 37213 19671 37216
rect 19613 37207 19671 37213
rect 19889 37213 19901 37216
rect 19935 37213 19947 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 19889 37207 19947 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21324 37216 22201 37244
rect 21324 37204 21330 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22833 37207 22891 37213
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 26053 37207 26111 37213
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 27985 37247 28043 37253
rect 27985 37244 27997 37247
rect 27764 37216 27997 37244
rect 27764 37204 27770 37216
rect 27985 37213 27997 37216
rect 28031 37213 28043 37247
rect 27985 37207 28043 37213
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29052 37216 29929 37244
rect 29052 37204 29058 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30432 37216 30573 37244
rect 30432 37204 30438 37216
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 30561 37207 30619 37213
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32272 37216 32505 37244
rect 32272 37204 32278 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 36722 37204 36728 37256
rect 36780 37244 36786 37256
rect 36909 37247 36967 37253
rect 36909 37244 36921 37247
rect 36780 37216 36921 37244
rect 36780 37204 36786 37216
rect 36909 37213 36921 37216
rect 36955 37213 36967 37247
rect 36909 37207 36967 37213
rect 37274 37204 37280 37256
rect 37332 37244 37338 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 37332 37216 38025 37244
rect 37332 37204 37338 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 4798 37136 4804 37188
rect 4856 37136 4862 37188
rect 8234 37148 9536 37176
rect 1636 37080 3280 37108
rect 3329 37111 3387 37117
rect 1636 37068 1642 37080
rect 3329 37077 3341 37111
rect 3375 37108 3387 37111
rect 3418 37108 3424 37120
rect 3375 37080 3424 37108
rect 3375 37077 3387 37080
rect 3329 37071 3387 37077
rect 3418 37068 3424 37080
rect 3476 37068 3482 37120
rect 5718 37108 5724 37120
rect 5679 37080 5724 37108
rect 5718 37068 5724 37080
rect 5776 37068 5782 37120
rect 8478 37108 8484 37120
rect 8439 37080 8484 37108
rect 8478 37068 8484 37080
rect 8536 37068 8542 37120
rect 9508 37108 9536 37148
rect 10594 37136 10600 37188
rect 10652 37136 10658 37188
rect 15838 37176 15844 37188
rect 10888 37148 11192 37176
rect 10888 37108 10916 37148
rect 9508 37080 10916 37108
rect 11164 37108 11192 37148
rect 13280 37148 15844 37176
rect 12342 37108 12348 37120
rect 11164 37080 12348 37108
rect 12342 37068 12348 37080
rect 12400 37068 12406 37120
rect 12618 37068 12624 37120
rect 12676 37108 12682 37120
rect 13280 37108 13308 37148
rect 15838 37136 15844 37148
rect 15896 37136 15902 37188
rect 20622 37136 20628 37188
rect 20680 37176 20686 37188
rect 20680 37148 22692 37176
rect 20680 37136 20686 37148
rect 12676 37080 13308 37108
rect 12676 37068 12682 37080
rect 13354 37068 13360 37120
rect 13412 37108 13418 37120
rect 13449 37111 13507 37117
rect 13449 37108 13461 37111
rect 13412 37080 13461 37108
rect 13412 37068 13418 37080
rect 13449 37077 13461 37080
rect 13495 37077 13507 37111
rect 13449 37071 13507 37077
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13596 37080 14473 37108
rect 13596 37068 13602 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 18138 37108 18144 37120
rect 18099 37080 18144 37108
rect 17037 37071 17095 37077
rect 18138 37068 18144 37080
rect 18196 37068 18202 37120
rect 19426 37108 19432 37120
rect 19387 37080 19432 37108
rect 19426 37068 19432 37080
rect 19484 37068 19490 37120
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 20346 37068 20352 37120
rect 20404 37108 20410 37120
rect 22664 37117 22692 37148
rect 23934 37136 23940 37188
rect 23992 37176 23998 37188
rect 23992 37148 25912 37176
rect 23992 37136 23998 37148
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 20404 37080 22017 37108
rect 20404 37068 20410 37080
rect 22005 37077 22017 37080
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 22649 37111 22707 37117
rect 22649 37077 22661 37111
rect 22695 37077 22707 37111
rect 22649 37071 22707 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 25884 37117 25912 37148
rect 31478 37136 31484 37188
rect 31536 37176 31542 37188
rect 31536 37148 35894 37176
rect 31536 37136 31542 37148
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25869 37111 25927 37117
rect 25869 37077 25881 37111
rect 25915 37077 25927 37111
rect 27798 37108 27804 37120
rect 27759 37080 27804 37108
rect 25869 37071 25927 37077
rect 27798 37068 27804 37080
rect 27856 37068 27862 37120
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 30374 37108 30380 37120
rect 30335 37080 30380 37108
rect 30374 37068 30380 37080
rect 30432 37068 30438 37120
rect 30650 37068 30656 37120
rect 30708 37108 30714 37120
rect 32309 37111 32367 37117
rect 32309 37108 32321 37111
rect 30708 37080 32321 37108
rect 30708 37068 30714 37080
rect 32309 37077 32321 37080
rect 32355 37077 32367 37111
rect 32309 37071 32367 37077
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 33597 37111 33655 37117
rect 33597 37108 33609 37111
rect 32456 37080 33609 37108
rect 32456 37068 32462 37080
rect 33597 37077 33609 37080
rect 33643 37077 33655 37111
rect 33597 37071 33655 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 34885 37111 34943 37117
rect 34885 37108 34897 37111
rect 34572 37080 34897 37108
rect 34572 37068 34578 37080
rect 34885 37077 34897 37080
rect 34931 37077 34943 37111
rect 35866 37108 35894 37148
rect 36725 37111 36783 37117
rect 36725 37108 36737 37111
rect 35866 37080 36737 37108
rect 34885 37071 34943 37077
rect 36725 37077 36737 37080
rect 36771 37077 36783 37111
rect 38194 37108 38200 37120
rect 38155 37080 38200 37108
rect 36725 37071 36783 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 5905 36907 5963 36913
rect 5905 36873 5917 36907
rect 5951 36904 5963 36907
rect 7374 36904 7380 36916
rect 5951 36876 7380 36904
rect 5951 36873 5963 36876
rect 5905 36867 5963 36873
rect 7374 36864 7380 36876
rect 7432 36864 7438 36916
rect 12342 36904 12348 36916
rect 7576 36876 12348 36904
rect 4430 36836 4436 36848
rect 3082 36808 4436 36836
rect 4430 36796 4436 36808
rect 4488 36796 4494 36848
rect 7576 36836 7604 36876
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 12526 36864 12532 36916
rect 12584 36904 12590 36916
rect 15933 36907 15991 36913
rect 15933 36904 15945 36907
rect 12584 36876 15945 36904
rect 12584 36864 12590 36876
rect 15933 36873 15945 36876
rect 15979 36873 15991 36907
rect 15933 36867 15991 36873
rect 16206 36864 16212 36916
rect 16264 36904 16270 36916
rect 16853 36907 16911 36913
rect 16853 36904 16865 36907
rect 16264 36876 16865 36904
rect 16264 36864 16270 36876
rect 16853 36873 16865 36876
rect 16899 36873 16911 36907
rect 16853 36867 16911 36873
rect 24670 36864 24676 36916
rect 24728 36904 24734 36916
rect 27798 36904 27804 36916
rect 24728 36876 27804 36904
rect 24728 36864 24734 36876
rect 27798 36864 27804 36876
rect 27856 36864 27862 36916
rect 5920 36808 7604 36836
rect 1578 36768 1584 36780
rect 1539 36740 1584 36768
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 3970 36728 3976 36780
rect 4028 36768 4034 36780
rect 4157 36771 4215 36777
rect 4157 36768 4169 36771
rect 4028 36740 4169 36768
rect 4028 36728 4034 36740
rect 4157 36737 4169 36740
rect 4203 36737 4215 36771
rect 5920 36768 5948 36808
rect 8662 36796 8668 36848
rect 8720 36836 8726 36848
rect 9674 36836 9680 36848
rect 8720 36808 9680 36836
rect 8720 36796 8726 36808
rect 9674 36796 9680 36808
rect 9732 36796 9738 36848
rect 10042 36796 10048 36848
rect 10100 36796 10106 36848
rect 12158 36836 12164 36848
rect 10888 36808 12164 36836
rect 5566 36740 5948 36768
rect 8418 36740 8524 36768
rect 4157 36731 4215 36737
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36700 1915 36703
rect 3234 36700 3240 36712
rect 1903 36672 3240 36700
rect 1903 36669 1915 36672
rect 1857 36663 1915 36669
rect 3234 36660 3240 36672
rect 3292 36660 3298 36712
rect 3602 36700 3608 36712
rect 3563 36672 3608 36700
rect 3602 36660 3608 36672
rect 3660 36660 3666 36712
rect 4433 36703 4491 36709
rect 4433 36669 4445 36703
rect 4479 36700 4491 36703
rect 4479 36672 6684 36700
rect 4479 36669 4491 36672
rect 4433 36663 4491 36669
rect 6656 36632 6684 36672
rect 6730 36660 6736 36712
rect 6788 36700 6794 36712
rect 7009 36703 7067 36709
rect 7009 36700 7021 36703
rect 6788 36672 7021 36700
rect 6788 36660 6794 36672
rect 7009 36669 7021 36672
rect 7055 36669 7067 36703
rect 7282 36700 7288 36712
rect 7243 36672 7288 36700
rect 7009 36663 7067 36669
rect 7282 36660 7288 36672
rect 7340 36660 7346 36712
rect 7374 36660 7380 36712
rect 7432 36700 7438 36712
rect 8018 36700 8024 36712
rect 7432 36672 8024 36700
rect 7432 36660 7438 36672
rect 8018 36660 8024 36672
rect 8076 36660 8082 36712
rect 6914 36632 6920 36644
rect 6656 36604 6920 36632
rect 6914 36592 6920 36604
rect 6972 36592 6978 36644
rect 8496 36564 8524 36740
rect 8754 36700 8760 36712
rect 8715 36672 8760 36700
rect 8754 36660 8760 36672
rect 8812 36660 8818 36712
rect 9122 36660 9128 36712
rect 9180 36700 9186 36712
rect 9309 36703 9367 36709
rect 9309 36700 9321 36703
rect 9180 36672 9321 36700
rect 9180 36660 9186 36672
rect 9309 36669 9321 36672
rect 9355 36669 9367 36703
rect 9582 36700 9588 36712
rect 9309 36663 9367 36669
rect 9416 36672 9588 36700
rect 8570 36592 8576 36644
rect 8628 36632 8634 36644
rect 9416 36632 9444 36672
rect 9582 36660 9588 36672
rect 9640 36660 9646 36712
rect 9674 36660 9680 36712
rect 9732 36700 9738 36712
rect 10888 36700 10916 36808
rect 12158 36796 12164 36808
rect 12216 36796 12222 36848
rect 12618 36796 12624 36848
rect 12676 36796 12682 36848
rect 13722 36796 13728 36848
rect 13780 36836 13786 36848
rect 14461 36839 14519 36845
rect 14461 36836 14473 36839
rect 13780 36808 14473 36836
rect 13780 36796 13786 36808
rect 14461 36805 14473 36808
rect 14507 36805 14519 36839
rect 39298 36836 39304 36848
rect 14461 36799 14519 36805
rect 37660 36808 39304 36836
rect 15562 36728 15568 36780
rect 15620 36728 15626 36780
rect 15838 36728 15844 36780
rect 15896 36768 15902 36780
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 15896 36740 17049 36768
rect 15896 36728 15902 36740
rect 17037 36737 17049 36740
rect 17083 36737 17095 36771
rect 17494 36768 17500 36780
rect 17455 36740 17500 36768
rect 17037 36731 17095 36737
rect 17494 36728 17500 36740
rect 17552 36768 17558 36780
rect 18141 36771 18199 36777
rect 18141 36768 18153 36771
rect 17552 36740 18153 36768
rect 17552 36728 17558 36740
rect 18141 36737 18153 36740
rect 18187 36768 18199 36771
rect 18785 36771 18843 36777
rect 18785 36768 18797 36771
rect 18187 36740 18797 36768
rect 18187 36737 18199 36740
rect 18141 36731 18199 36737
rect 18785 36737 18797 36740
rect 18831 36737 18843 36771
rect 18785 36731 18843 36737
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 37660 36777 37688 36808
rect 39298 36796 39304 36808
rect 39356 36796 39362 36848
rect 19613 36771 19671 36777
rect 19613 36768 19625 36771
rect 19392 36740 19625 36768
rect 19392 36728 19398 36740
rect 19613 36737 19625 36740
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 37645 36771 37703 36777
rect 37645 36737 37657 36771
rect 37691 36737 37703 36771
rect 37645 36731 37703 36737
rect 38010 36728 38016 36780
rect 38068 36768 38074 36780
rect 38289 36771 38347 36777
rect 38289 36768 38301 36771
rect 38068 36740 38301 36768
rect 38068 36728 38074 36740
rect 38289 36737 38301 36740
rect 38335 36737 38347 36771
rect 38289 36731 38347 36737
rect 9732 36672 10916 36700
rect 9732 36660 9738 36672
rect 11054 36660 11060 36712
rect 11112 36700 11118 36712
rect 11885 36703 11943 36709
rect 11885 36700 11897 36703
rect 11112 36672 11897 36700
rect 11112 36660 11118 36672
rect 11885 36669 11897 36672
rect 11931 36669 11943 36703
rect 11885 36663 11943 36669
rect 12161 36703 12219 36709
rect 12161 36669 12173 36703
rect 12207 36700 12219 36703
rect 13354 36700 13360 36712
rect 12207 36672 13360 36700
rect 12207 36669 12219 36672
rect 12161 36663 12219 36669
rect 11790 36632 11796 36644
rect 8628 36604 9444 36632
rect 10980 36604 11796 36632
rect 8628 36592 8634 36604
rect 10980 36564 11008 36604
rect 11790 36592 11796 36604
rect 11848 36592 11854 36644
rect 8496 36536 11008 36564
rect 11057 36567 11115 36573
rect 11057 36533 11069 36567
rect 11103 36564 11115 36567
rect 11146 36564 11152 36576
rect 11103 36536 11152 36564
rect 11103 36533 11115 36536
rect 11057 36527 11115 36533
rect 11146 36524 11152 36536
rect 11204 36524 11210 36576
rect 11900 36564 11928 36663
rect 13354 36660 13360 36672
rect 13412 36660 13418 36712
rect 14182 36700 14188 36712
rect 13556 36672 14188 36700
rect 13556 36564 13584 36672
rect 14182 36660 14188 36672
rect 14240 36660 14246 36712
rect 15654 36660 15660 36712
rect 15712 36700 15718 36712
rect 18233 36703 18291 36709
rect 18233 36700 18245 36703
rect 15712 36672 18245 36700
rect 15712 36660 15718 36672
rect 18233 36669 18245 36672
rect 18279 36669 18291 36703
rect 18233 36663 18291 36669
rect 15470 36592 15476 36644
rect 15528 36632 15534 36644
rect 18877 36635 18935 36641
rect 18877 36632 18889 36635
rect 15528 36604 18889 36632
rect 15528 36592 15534 36604
rect 18877 36601 18889 36604
rect 18923 36601 18935 36635
rect 18877 36595 18935 36601
rect 35894 36592 35900 36644
rect 35952 36632 35958 36644
rect 38105 36635 38163 36641
rect 38105 36632 38117 36635
rect 35952 36604 38117 36632
rect 35952 36592 35958 36604
rect 38105 36601 38117 36604
rect 38151 36601 38163 36635
rect 38105 36595 38163 36601
rect 11900 36536 13584 36564
rect 13630 36524 13636 36576
rect 13688 36564 13694 36576
rect 13688 36536 13733 36564
rect 13688 36524 13694 36536
rect 14274 36524 14280 36576
rect 14332 36564 14338 36576
rect 16758 36564 16764 36576
rect 14332 36536 16764 36564
rect 14332 36524 14338 36536
rect 16758 36524 16764 36536
rect 16816 36524 16822 36576
rect 17586 36564 17592 36576
rect 17547 36536 17592 36564
rect 17586 36524 17592 36536
rect 17644 36524 17650 36576
rect 19334 36524 19340 36576
rect 19392 36564 19398 36576
rect 19429 36567 19487 36573
rect 19429 36564 19441 36567
rect 19392 36536 19441 36564
rect 19392 36524 19398 36536
rect 19429 36533 19441 36536
rect 19475 36533 19487 36567
rect 19429 36527 19487 36533
rect 35986 36524 35992 36576
rect 36044 36564 36050 36576
rect 37461 36567 37519 36573
rect 37461 36564 37473 36567
rect 36044 36536 37473 36564
rect 36044 36524 36050 36536
rect 37461 36533 37473 36536
rect 37507 36533 37519 36567
rect 37461 36527 37519 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 5718 36360 5724 36372
rect 3896 36332 5724 36360
rect 1578 36224 1584 36236
rect 1539 36196 1584 36224
rect 1578 36184 1584 36196
rect 1636 36184 1642 36236
rect 1857 36227 1915 36233
rect 1857 36193 1869 36227
rect 1903 36224 1915 36227
rect 3896 36224 3924 36332
rect 5718 36320 5724 36332
rect 5776 36320 5782 36372
rect 8294 36320 8300 36372
rect 8352 36360 8358 36372
rect 10137 36363 10195 36369
rect 8352 36332 9674 36360
rect 8352 36320 8358 36332
rect 9122 36252 9128 36304
rect 9180 36252 9186 36304
rect 9646 36292 9674 36332
rect 10137 36329 10149 36363
rect 10183 36360 10195 36363
rect 10318 36360 10324 36372
rect 10183 36332 10324 36360
rect 10183 36329 10195 36332
rect 10137 36323 10195 36329
rect 10318 36320 10324 36332
rect 10376 36320 10382 36372
rect 10428 36332 12020 36360
rect 10428 36292 10456 36332
rect 9646 36264 10456 36292
rect 1903 36196 3924 36224
rect 1903 36193 1915 36196
rect 1857 36187 1915 36193
rect 3970 36184 3976 36236
rect 4028 36224 4034 36236
rect 4433 36227 4491 36233
rect 4433 36224 4445 36227
rect 4028 36196 4445 36224
rect 4028 36184 4034 36196
rect 4433 36193 4445 36196
rect 4479 36224 4491 36227
rect 6730 36224 6736 36236
rect 4479 36196 6736 36224
rect 4479 36193 4491 36196
rect 4433 36187 4491 36193
rect 6730 36184 6736 36196
rect 6788 36184 6794 36236
rect 7006 36184 7012 36236
rect 7064 36224 7070 36236
rect 7558 36224 7564 36236
rect 7064 36196 7564 36224
rect 7064 36184 7070 36196
rect 7558 36184 7564 36196
rect 7616 36184 7622 36236
rect 7742 36184 7748 36236
rect 7800 36224 7806 36236
rect 8202 36224 8208 36236
rect 7800 36196 8208 36224
rect 7800 36184 7806 36196
rect 8202 36184 8208 36196
rect 8260 36184 8266 36236
rect 8294 36184 8300 36236
rect 8352 36184 8358 36236
rect 8481 36227 8539 36233
rect 8481 36193 8493 36227
rect 8527 36224 8539 36227
rect 8846 36224 8852 36236
rect 8527 36196 8852 36224
rect 8527 36193 8539 36196
rect 8481 36187 8539 36193
rect 8312 36156 8340 36184
rect 8142 36128 8340 36156
rect 8386 36116 8392 36168
rect 8444 36156 8450 36168
rect 8496 36156 8524 36187
rect 8846 36184 8852 36196
rect 8904 36184 8910 36236
rect 9140 36224 9168 36252
rect 10689 36227 10747 36233
rect 10689 36224 10701 36227
rect 9140 36196 10701 36224
rect 10689 36193 10701 36196
rect 10735 36224 10747 36227
rect 11054 36224 11060 36236
rect 10735 36196 11060 36224
rect 10735 36193 10747 36196
rect 10689 36187 10747 36193
rect 11054 36184 11060 36196
rect 11112 36184 11118 36236
rect 11992 36224 12020 36332
rect 12066 36320 12072 36372
rect 12124 36360 12130 36372
rect 15470 36360 15476 36372
rect 12124 36332 15476 36360
rect 12124 36320 12130 36332
rect 15470 36320 15476 36332
rect 15528 36320 15534 36372
rect 15746 36360 15752 36372
rect 15707 36332 15752 36360
rect 15746 36320 15752 36332
rect 15804 36320 15810 36372
rect 16758 36320 16764 36372
rect 16816 36360 16822 36372
rect 17957 36363 18015 36369
rect 17957 36360 17969 36363
rect 16816 36332 17969 36360
rect 16816 36320 16822 36332
rect 17957 36329 17969 36332
rect 18003 36329 18015 36363
rect 17957 36323 18015 36329
rect 12158 36252 12164 36304
rect 12216 36292 12222 36304
rect 14274 36292 14280 36304
rect 12216 36264 14280 36292
rect 12216 36252 12222 36264
rect 14274 36252 14280 36264
rect 14332 36252 14338 36304
rect 14461 36295 14519 36301
rect 14461 36261 14473 36295
rect 14507 36292 14519 36295
rect 16850 36292 16856 36304
rect 14507 36264 16856 36292
rect 14507 36261 14519 36264
rect 14461 36255 14519 36261
rect 16850 36252 16856 36264
rect 16908 36252 16914 36304
rect 17586 36224 17592 36236
rect 11992 36196 17592 36224
rect 17586 36184 17592 36196
rect 17644 36184 17650 36236
rect 8444 36128 8524 36156
rect 9125 36159 9183 36165
rect 8444 36116 8450 36128
rect 9125 36125 9137 36159
rect 9171 36156 9183 36159
rect 9858 36156 9864 36168
rect 9171 36128 9864 36156
rect 9171 36125 9183 36128
rect 9125 36119 9183 36125
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 9953 36159 10011 36165
rect 9953 36125 9965 36159
rect 9999 36125 10011 36159
rect 9953 36119 10011 36125
rect 3878 36088 3884 36100
rect 3082 36060 3884 36088
rect 3878 36048 3884 36060
rect 3936 36048 3942 36100
rect 4614 36048 4620 36100
rect 4672 36088 4678 36100
rect 4709 36091 4767 36097
rect 4709 36088 4721 36091
rect 4672 36060 4721 36088
rect 4672 36048 4678 36060
rect 4709 36057 4721 36060
rect 4755 36057 4767 36091
rect 4982 36088 4988 36100
rect 4709 36051 4767 36057
rect 4816 36060 4988 36088
rect 3329 36023 3387 36029
rect 3329 35989 3341 36023
rect 3375 36020 3387 36023
rect 4816 36020 4844 36060
rect 4982 36048 4988 36060
rect 5040 36048 5046 36100
rect 5934 36060 6960 36088
rect 3375 35992 4844 36020
rect 3375 35989 3387 35992
rect 3329 35983 3387 35989
rect 4890 35980 4896 36032
rect 4948 36020 4954 36032
rect 6181 36023 6239 36029
rect 6181 36020 6193 36023
rect 4948 35992 6193 36020
rect 4948 35980 4954 35992
rect 6181 35989 6193 35992
rect 6227 35989 6239 36023
rect 6932 36020 6960 36060
rect 7006 36048 7012 36100
rect 7064 36088 7070 36100
rect 7064 36060 7109 36088
rect 7064 36048 7070 36060
rect 8294 36048 8300 36100
rect 8352 36088 8358 36100
rect 8352 36060 9352 36088
rect 8352 36048 8358 36060
rect 9214 36020 9220 36032
rect 6932 35992 9220 36020
rect 6181 35983 6239 35989
rect 9214 35980 9220 35992
rect 9272 35980 9278 36032
rect 9324 36029 9352 36060
rect 9309 36023 9367 36029
rect 9309 35989 9321 36023
rect 9355 35989 9367 36023
rect 9968 36020 9996 36119
rect 12434 36116 12440 36168
rect 12492 36156 12498 36168
rect 13357 36159 13415 36165
rect 12492 36128 13308 36156
rect 12492 36116 12498 36128
rect 10962 36088 10968 36100
rect 10923 36060 10968 36088
rect 10962 36048 10968 36060
rect 11020 36048 11026 36100
rect 11422 36048 11428 36100
rect 11480 36048 11486 36100
rect 12986 36088 12992 36100
rect 12268 36060 12992 36088
rect 12268 36020 12296 36060
rect 12986 36048 12992 36060
rect 13044 36048 13050 36100
rect 9968 35992 12296 36020
rect 9309 35983 9367 35989
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 12492 35992 12537 36020
rect 12492 35980 12498 35992
rect 12618 35980 12624 36032
rect 12676 36020 12682 36032
rect 13173 36023 13231 36029
rect 13173 36020 13185 36023
rect 12676 35992 13185 36020
rect 12676 35980 12682 35992
rect 13173 35989 13185 35992
rect 13219 35989 13231 36023
rect 13280 36020 13308 36128
rect 13357 36125 13369 36159
rect 13403 36156 13415 36159
rect 13630 36156 13636 36168
rect 13403 36128 13636 36156
rect 13403 36125 13415 36128
rect 13357 36119 13415 36125
rect 13630 36116 13636 36128
rect 13688 36116 13694 36168
rect 14642 36156 14648 36168
rect 14603 36128 14648 36156
rect 14642 36116 14648 36128
rect 14700 36116 14706 36168
rect 15105 36159 15163 36165
rect 15105 36125 15117 36159
rect 15151 36156 15163 36159
rect 15838 36156 15844 36168
rect 15151 36128 15844 36156
rect 15151 36125 15163 36128
rect 15105 36119 15163 36125
rect 15838 36116 15844 36128
rect 15896 36116 15902 36168
rect 15933 36159 15991 36165
rect 15933 36125 15945 36159
rect 15979 36125 15991 36159
rect 16574 36156 16580 36168
rect 16535 36128 16580 36156
rect 15933 36119 15991 36125
rect 14734 36048 14740 36100
rect 14792 36088 14798 36100
rect 15948 36088 15976 36119
rect 16574 36116 16580 36128
rect 16632 36116 16638 36168
rect 17037 36159 17095 36165
rect 17037 36125 17049 36159
rect 17083 36156 17095 36159
rect 17494 36156 17500 36168
rect 17083 36128 17500 36156
rect 17083 36125 17095 36128
rect 17037 36119 17095 36125
rect 17494 36116 17500 36128
rect 17552 36116 17558 36168
rect 17972 36156 18000 36323
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 17972 36128 18521 36156
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 37182 36116 37188 36168
rect 37240 36156 37246 36168
rect 38289 36159 38347 36165
rect 38289 36156 38301 36159
rect 37240 36128 38301 36156
rect 37240 36116 37246 36128
rect 38289 36125 38301 36128
rect 38335 36125 38347 36159
rect 38289 36119 38347 36125
rect 17126 36088 17132 36100
rect 14792 36060 15976 36088
rect 17087 36060 17132 36088
rect 14792 36048 14798 36060
rect 17126 36048 17132 36060
rect 17184 36048 17190 36100
rect 13538 36020 13544 36032
rect 13280 35992 13544 36020
rect 13173 35983 13231 35989
rect 13538 35980 13544 35992
rect 13596 35980 13602 36032
rect 15197 36023 15255 36029
rect 15197 35989 15209 36023
rect 15243 36020 15255 36023
rect 15378 36020 15384 36032
rect 15243 35992 15384 36020
rect 15243 35989 15255 35992
rect 15197 35983 15255 35989
rect 15378 35980 15384 35992
rect 15436 35980 15442 36032
rect 16298 35980 16304 36032
rect 16356 36020 16362 36032
rect 16393 36023 16451 36029
rect 16393 36020 16405 36023
rect 16356 35992 16405 36020
rect 16356 35980 16362 35992
rect 16393 35989 16405 35992
rect 16439 35989 16451 36023
rect 17586 36020 17592 36032
rect 17547 35992 17592 36020
rect 16393 35983 16451 35989
rect 17586 35980 17592 35992
rect 17644 35980 17650 36032
rect 18325 36023 18383 36029
rect 18325 35989 18337 36023
rect 18371 36020 18383 36023
rect 18414 36020 18420 36032
rect 18371 35992 18420 36020
rect 18371 35989 18383 35992
rect 18325 35983 18383 35989
rect 18414 35980 18420 35992
rect 18472 35980 18478 36032
rect 36078 35980 36084 36032
rect 36136 36020 36142 36032
rect 38105 36023 38163 36029
rect 38105 36020 38117 36023
rect 36136 35992 38117 36020
rect 36136 35980 36142 35992
rect 38105 35989 38117 35992
rect 38151 35989 38163 36023
rect 38105 35983 38163 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 5810 35776 5816 35828
rect 5868 35816 5874 35828
rect 5905 35819 5963 35825
rect 5905 35816 5917 35819
rect 5868 35788 5917 35816
rect 5868 35776 5874 35788
rect 5905 35785 5917 35788
rect 5951 35785 5963 35819
rect 12250 35816 12256 35828
rect 5905 35779 5963 35785
rect 7484 35788 12256 35816
rect 7484 35748 7512 35788
rect 12250 35776 12256 35788
rect 12308 35776 12314 35828
rect 14645 35819 14703 35825
rect 12360 35788 14596 35816
rect 10686 35748 10692 35760
rect 5736 35720 7512 35748
rect 10626 35720 10692 35748
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 1946 35680 1952 35692
rect 1903 35652 1952 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 1946 35640 1952 35652
rect 2004 35640 2010 35692
rect 5736 35689 5764 35720
rect 10686 35708 10692 35720
rect 10744 35708 10750 35760
rect 12360 35748 12388 35788
rect 10796 35720 12388 35748
rect 14568 35748 14596 35788
rect 14645 35785 14657 35819
rect 14691 35816 14703 35819
rect 14734 35816 14740 35828
rect 14691 35788 14740 35816
rect 14691 35785 14703 35788
rect 14645 35779 14703 35785
rect 14734 35776 14740 35788
rect 14792 35776 14798 35828
rect 15102 35776 15108 35828
rect 15160 35816 15166 35828
rect 15197 35819 15255 35825
rect 15197 35816 15209 35819
rect 15160 35788 15209 35816
rect 15160 35776 15166 35788
rect 15197 35785 15209 35788
rect 15243 35785 15255 35819
rect 15197 35779 15255 35785
rect 15286 35776 15292 35828
rect 15344 35816 15350 35828
rect 17126 35816 17132 35828
rect 15344 35788 17132 35816
rect 15344 35776 15350 35788
rect 17126 35776 17132 35788
rect 17184 35776 17190 35828
rect 17586 35748 17592 35760
rect 14568 35720 17592 35748
rect 5721 35683 5779 35689
rect 2133 35615 2191 35621
rect 2133 35581 2145 35615
rect 2179 35612 2191 35615
rect 2958 35612 2964 35624
rect 2179 35584 2964 35612
rect 2179 35581 2191 35584
rect 2133 35575 2191 35581
rect 2958 35572 2964 35584
rect 3016 35572 3022 35624
rect 3053 35615 3111 35621
rect 3053 35581 3065 35615
rect 3099 35581 3111 35615
rect 3326 35612 3332 35624
rect 3287 35584 3332 35612
rect 3053 35575 3111 35581
rect 1578 35504 1584 35556
rect 1636 35544 1642 35556
rect 3068 35544 3096 35575
rect 3326 35572 3332 35584
rect 3384 35572 3390 35624
rect 4448 35612 4476 35666
rect 5721 35649 5733 35683
rect 5767 35649 5779 35683
rect 5721 35643 5779 35649
rect 6730 35640 6736 35692
rect 6788 35680 6794 35692
rect 6825 35683 6883 35689
rect 6825 35680 6837 35683
rect 6788 35652 6837 35680
rect 6788 35640 6794 35652
rect 6825 35649 6837 35652
rect 6871 35649 6883 35683
rect 6825 35643 6883 35649
rect 5902 35612 5908 35624
rect 4448 35584 5908 35612
rect 5902 35572 5908 35584
rect 5960 35572 5966 35624
rect 6178 35572 6184 35624
rect 6236 35612 6242 35624
rect 7101 35615 7159 35621
rect 7101 35612 7113 35615
rect 6236 35584 7113 35612
rect 6236 35572 6242 35584
rect 7101 35581 7113 35584
rect 7147 35612 7159 35615
rect 7834 35612 7840 35624
rect 7147 35584 7840 35612
rect 7147 35581 7159 35584
rect 7101 35575 7159 35581
rect 7834 35572 7840 35584
rect 7892 35572 7898 35624
rect 8220 35544 8248 35666
rect 8570 35612 8576 35624
rect 8531 35584 8576 35612
rect 8570 35572 8576 35584
rect 8628 35572 8634 35624
rect 9122 35612 9128 35624
rect 9083 35584 9128 35612
rect 9122 35572 9128 35584
rect 9180 35572 9186 35624
rect 9401 35615 9459 35621
rect 9401 35581 9413 35615
rect 9447 35612 9459 35615
rect 10410 35612 10416 35624
rect 9447 35584 10416 35612
rect 9447 35581 9459 35584
rect 9401 35575 9459 35581
rect 10410 35572 10416 35584
rect 10468 35572 10474 35624
rect 1636 35516 3096 35544
rect 4632 35516 6960 35544
rect 8220 35516 9260 35544
rect 1636 35504 1642 35516
rect 3510 35436 3516 35488
rect 3568 35476 3574 35488
rect 4632 35476 4660 35516
rect 3568 35448 4660 35476
rect 3568 35436 3574 35448
rect 4706 35436 4712 35488
rect 4764 35476 4770 35488
rect 4801 35479 4859 35485
rect 4801 35476 4813 35479
rect 4764 35448 4813 35476
rect 4764 35436 4770 35448
rect 4801 35445 4813 35448
rect 4847 35476 4859 35479
rect 5074 35476 5080 35488
rect 4847 35448 5080 35476
rect 4847 35445 4859 35448
rect 4801 35439 4859 35445
rect 5074 35436 5080 35448
rect 5132 35436 5138 35488
rect 6932 35476 6960 35516
rect 8386 35476 8392 35488
rect 6932 35448 8392 35476
rect 8386 35436 8392 35448
rect 8444 35436 8450 35488
rect 9232 35476 9260 35516
rect 10796 35476 10824 35720
rect 17586 35708 17592 35720
rect 17644 35708 17650 35760
rect 14093 35683 14151 35689
rect 13110 35652 14044 35680
rect 11054 35572 11060 35624
rect 11112 35612 11118 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11112 35584 11713 35612
rect 11112 35572 11118 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11977 35615 12035 35621
rect 11977 35612 11989 35615
rect 11701 35575 11759 35581
rect 11795 35584 11989 35612
rect 10962 35504 10968 35556
rect 11020 35544 11026 35556
rect 11795 35544 11823 35584
rect 11977 35581 11989 35584
rect 12023 35581 12035 35615
rect 11977 35575 12035 35581
rect 12066 35572 12072 35624
rect 12124 35612 12130 35624
rect 13449 35615 13507 35621
rect 13449 35612 13461 35615
rect 12124 35584 13461 35612
rect 12124 35572 12130 35584
rect 13449 35581 13461 35584
rect 13495 35581 13507 35615
rect 14016 35612 14044 35652
rect 14093 35649 14105 35683
rect 14139 35680 14151 35683
rect 14458 35680 14464 35692
rect 14139 35652 14464 35680
rect 14139 35649 14151 35652
rect 14093 35643 14151 35649
rect 14458 35640 14464 35652
rect 14516 35640 14522 35692
rect 14553 35683 14611 35689
rect 14553 35649 14565 35683
rect 14599 35680 14611 35683
rect 14918 35680 14924 35692
rect 14599 35652 14924 35680
rect 14599 35649 14611 35652
rect 14553 35643 14611 35649
rect 14918 35640 14924 35652
rect 14976 35640 14982 35692
rect 15378 35680 15384 35692
rect 15339 35652 15384 35680
rect 15378 35640 15384 35652
rect 15436 35640 15442 35692
rect 15470 35640 15476 35692
rect 15528 35680 15534 35692
rect 15841 35683 15899 35689
rect 15841 35680 15853 35683
rect 15528 35652 15853 35680
rect 15528 35640 15534 35652
rect 15841 35649 15853 35652
rect 15887 35680 15899 35683
rect 16482 35680 16488 35692
rect 15887 35652 16488 35680
rect 15887 35649 15899 35652
rect 15841 35643 15899 35649
rect 16482 35640 16488 35652
rect 16540 35680 16546 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16540 35652 16865 35680
rect 16540 35640 16546 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 17494 35680 17500 35692
rect 17455 35652 17500 35680
rect 16853 35643 16911 35649
rect 17494 35640 17500 35652
rect 17552 35640 17558 35692
rect 18230 35612 18236 35624
rect 14016 35584 18236 35612
rect 13449 35575 13507 35581
rect 18230 35572 18236 35584
rect 18288 35572 18294 35624
rect 11020 35516 11823 35544
rect 11020 35504 11026 35516
rect 12986 35504 12992 35556
rect 13044 35544 13050 35556
rect 13909 35547 13967 35553
rect 13909 35544 13921 35547
rect 13044 35516 13921 35544
rect 13044 35504 13050 35516
rect 13909 35513 13921 35516
rect 13955 35513 13967 35547
rect 16574 35544 16580 35556
rect 13909 35507 13967 35513
rect 14476 35516 16580 35544
rect 9232 35448 10824 35476
rect 10870 35436 10876 35488
rect 10928 35476 10934 35488
rect 10928 35448 10973 35476
rect 10928 35436 10934 35448
rect 11146 35436 11152 35488
rect 11204 35476 11210 35488
rect 14476 35476 14504 35516
rect 16574 35504 16580 35516
rect 16632 35504 16638 35556
rect 11204 35448 14504 35476
rect 11204 35436 11210 35448
rect 14550 35436 14556 35488
rect 14608 35476 14614 35488
rect 15102 35476 15108 35488
rect 14608 35448 15108 35476
rect 14608 35436 14614 35448
rect 15102 35436 15108 35448
rect 15160 35436 15166 35488
rect 15930 35476 15936 35488
rect 15891 35448 15936 35476
rect 15930 35436 15936 35448
rect 15988 35436 15994 35488
rect 16942 35476 16948 35488
rect 16903 35448 16948 35476
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 17586 35476 17592 35488
rect 17547 35448 17592 35476
rect 17586 35436 17592 35448
rect 17644 35436 17650 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 4696 35275 4754 35281
rect 4696 35241 4708 35275
rect 4742 35272 4754 35275
rect 6362 35272 6368 35284
rect 4742 35244 6368 35272
rect 4742 35241 4754 35244
rect 4696 35235 4754 35241
rect 6362 35232 6368 35244
rect 6420 35232 6426 35284
rect 6638 35232 6644 35284
rect 6696 35272 6702 35284
rect 6696 35244 10916 35272
rect 6696 35232 6702 35244
rect 6178 35204 6184 35216
rect 6139 35176 6184 35204
rect 6178 35164 6184 35176
rect 6236 35164 6242 35216
rect 1578 35136 1584 35148
rect 1539 35108 1584 35136
rect 1578 35096 1584 35108
rect 1636 35096 1642 35148
rect 1857 35139 1915 35145
rect 1857 35105 1869 35139
rect 1903 35136 1915 35139
rect 3234 35136 3240 35148
rect 1903 35108 3240 35136
rect 1903 35105 1915 35108
rect 1857 35099 1915 35105
rect 3234 35096 3240 35108
rect 3292 35136 3298 35148
rect 3418 35136 3424 35148
rect 3292 35108 3424 35136
rect 3292 35096 3298 35108
rect 3418 35096 3424 35108
rect 3476 35096 3482 35148
rect 3970 35096 3976 35148
rect 4028 35136 4034 35148
rect 4433 35139 4491 35145
rect 4433 35136 4445 35139
rect 4028 35108 4445 35136
rect 4028 35096 4034 35108
rect 4433 35105 4445 35108
rect 4479 35136 4491 35139
rect 6641 35139 6699 35145
rect 6641 35136 6653 35139
rect 4479 35108 6653 35136
rect 4479 35105 4491 35108
rect 4433 35099 4491 35105
rect 6641 35105 6653 35108
rect 6687 35136 6699 35139
rect 9122 35136 9128 35148
rect 6687 35108 9128 35136
rect 6687 35105 6699 35108
rect 6641 35099 6699 35105
rect 9122 35096 9128 35108
rect 9180 35096 9186 35148
rect 9398 35136 9404 35148
rect 9359 35108 9404 35136
rect 9398 35096 9404 35108
rect 9456 35096 9462 35148
rect 10888 35136 10916 35244
rect 11514 35232 11520 35284
rect 11572 35272 11578 35284
rect 15930 35272 15936 35284
rect 11572 35244 15936 35272
rect 11572 35232 11578 35244
rect 15930 35232 15936 35244
rect 15988 35232 15994 35284
rect 22741 35275 22799 35281
rect 22741 35241 22753 35275
rect 22787 35272 22799 35275
rect 24578 35272 24584 35284
rect 22787 35244 24584 35272
rect 22787 35241 22799 35244
rect 22741 35235 22799 35241
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 12802 35164 12808 35216
rect 12860 35204 12866 35216
rect 17405 35207 17463 35213
rect 12860 35176 14412 35204
rect 12860 35164 12866 35176
rect 14090 35136 14096 35148
rect 10888 35108 14096 35136
rect 14090 35096 14096 35108
rect 14148 35096 14154 35148
rect 14182 35096 14188 35148
rect 14240 35136 14246 35148
rect 14277 35139 14335 35145
rect 14277 35136 14289 35139
rect 14240 35108 14289 35136
rect 14240 35096 14246 35108
rect 14277 35105 14289 35108
rect 14323 35105 14335 35139
rect 14384 35136 14412 35176
rect 17405 35173 17417 35207
rect 17451 35204 17463 35207
rect 20070 35204 20076 35216
rect 17451 35176 20076 35204
rect 17451 35173 17463 35176
rect 17405 35167 17463 35173
rect 20070 35164 20076 35176
rect 20128 35164 20134 35216
rect 17862 35136 17868 35148
rect 14384 35108 17868 35136
rect 14277 35099 14335 35105
rect 17862 35096 17868 35108
rect 17920 35096 17926 35148
rect 8018 35028 8024 35080
rect 8076 35028 8082 35080
rect 10502 35028 10508 35080
rect 10560 35028 10566 35080
rect 11054 35028 11060 35080
rect 11112 35068 11118 35080
rect 11517 35071 11575 35077
rect 11517 35068 11529 35071
rect 11112 35040 11529 35068
rect 11112 35028 11118 35040
rect 11517 35037 11529 35040
rect 11563 35037 11575 35071
rect 16114 35068 16120 35080
rect 15686 35040 16120 35068
rect 11517 35031 11575 35037
rect 16114 35028 16120 35040
rect 16172 35028 16178 35080
rect 16390 35028 16396 35080
rect 16448 35068 16454 35080
rect 16485 35071 16543 35077
rect 16485 35068 16497 35071
rect 16448 35040 16497 35068
rect 16448 35028 16454 35040
rect 16485 35037 16497 35040
rect 16531 35037 16543 35071
rect 16485 35031 16543 35037
rect 17589 35071 17647 35077
rect 17589 35037 17601 35071
rect 17635 35068 17647 35071
rect 17678 35068 17684 35080
rect 17635 35040 17684 35068
rect 17635 35037 17647 35040
rect 17589 35031 17647 35037
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 22922 35068 22928 35080
rect 22883 35040 22928 35068
rect 22922 35028 22928 35040
rect 22980 35028 22986 35080
rect 34238 35028 34244 35080
rect 34296 35068 34302 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 34296 35040 38025 35068
rect 34296 35028 34302 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 3082 34972 5028 35000
rect 5934 34972 6868 35000
rect 3326 34932 3332 34944
rect 3287 34904 3332 34932
rect 3326 34892 3332 34904
rect 3384 34892 3390 34944
rect 5000 34932 5028 34972
rect 6086 34932 6092 34944
rect 5000 34904 6092 34932
rect 6086 34892 6092 34904
rect 6144 34892 6150 34944
rect 6840 34932 6868 34972
rect 6914 34960 6920 35012
rect 6972 35000 6978 35012
rect 6972 34972 7017 35000
rect 8220 34972 8524 35000
rect 6972 34960 6978 34972
rect 8220 34932 8248 34972
rect 8386 34932 8392 34944
rect 6840 34904 8248 34932
rect 8347 34904 8392 34932
rect 8386 34892 8392 34904
rect 8444 34892 8450 34944
rect 8496 34932 8524 34972
rect 10704 34972 11008 35000
rect 10704 34932 10732 34972
rect 8496 34904 10732 34932
rect 10778 34892 10784 34944
rect 10836 34932 10842 34944
rect 10873 34935 10931 34941
rect 10873 34932 10885 34935
rect 10836 34904 10885 34932
rect 10836 34892 10842 34904
rect 10873 34901 10885 34904
rect 10919 34901 10931 34935
rect 10980 34932 11008 34972
rect 11146 34960 11152 35012
rect 11204 35000 11210 35012
rect 11793 35003 11851 35009
rect 11793 35000 11805 35003
rect 11204 34972 11805 35000
rect 11204 34960 11210 34972
rect 11793 34969 11805 34972
rect 11839 34969 11851 35003
rect 11793 34963 11851 34969
rect 12526 34960 12532 35012
rect 12584 34960 12590 35012
rect 14550 35000 14556 35012
rect 14511 34972 14556 35000
rect 14550 34960 14556 34972
rect 14608 34960 14614 35012
rect 16577 35003 16635 35009
rect 16577 35000 16589 35003
rect 15856 34972 16589 35000
rect 13170 34932 13176 34944
rect 10980 34904 13176 34932
rect 10873 34895 10931 34901
rect 13170 34892 13176 34904
rect 13228 34892 13234 34944
rect 13262 34892 13268 34944
rect 13320 34932 13326 34944
rect 13320 34904 13365 34932
rect 13320 34892 13326 34904
rect 13446 34892 13452 34944
rect 13504 34932 13510 34944
rect 15856 34932 15884 34972
rect 16577 34969 16589 34972
rect 16623 34969 16635 35003
rect 16577 34963 16635 34969
rect 13504 34904 15884 34932
rect 13504 34892 13510 34904
rect 15930 34892 15936 34944
rect 15988 34932 15994 34944
rect 16025 34935 16083 34941
rect 16025 34932 16037 34935
rect 15988 34904 16037 34932
rect 15988 34892 15994 34904
rect 16025 34901 16037 34904
rect 16071 34901 16083 34935
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 16025 34895 16083 34901
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2682 34688 2688 34740
rect 2740 34728 2746 34740
rect 13998 34728 14004 34740
rect 2740 34700 14004 34728
rect 2740 34688 2746 34700
rect 13998 34688 14004 34700
rect 14056 34688 14062 34740
rect 14090 34688 14096 34740
rect 14148 34728 14154 34740
rect 14829 34731 14887 34737
rect 14829 34728 14841 34731
rect 14148 34700 14841 34728
rect 14148 34688 14154 34700
rect 14829 34697 14841 34700
rect 14875 34697 14887 34731
rect 14829 34691 14887 34697
rect 15010 34688 15016 34740
rect 15068 34728 15074 34740
rect 17494 34728 17500 34740
rect 15068 34700 17500 34728
rect 15068 34688 15074 34700
rect 17494 34688 17500 34700
rect 17552 34688 17558 34740
rect 18230 34728 18236 34740
rect 18191 34700 18236 34728
rect 18230 34688 18236 34700
rect 18288 34688 18294 34740
rect 2133 34663 2191 34669
rect 2133 34629 2145 34663
rect 2179 34660 2191 34663
rect 4706 34660 4712 34672
rect 2179 34632 4712 34660
rect 2179 34629 2191 34632
rect 2133 34623 2191 34629
rect 4706 34620 4712 34632
rect 4764 34620 4770 34672
rect 7650 34660 7656 34672
rect 5920 34632 7656 34660
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 1946 34592 1952 34604
rect 1903 34564 1952 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 1946 34552 1952 34564
rect 2004 34592 2010 34604
rect 2682 34592 2688 34604
rect 2004 34564 2688 34592
rect 2004 34552 2010 34564
rect 2682 34552 2688 34564
rect 2740 34592 2746 34604
rect 2777 34595 2835 34601
rect 2777 34592 2789 34595
rect 2740 34564 2789 34592
rect 2740 34552 2746 34564
rect 2777 34561 2789 34564
rect 2823 34561 2835 34595
rect 2777 34555 2835 34561
rect 3970 34552 3976 34604
rect 4028 34592 4034 34604
rect 4157 34595 4215 34601
rect 4157 34592 4169 34595
rect 4028 34564 4169 34592
rect 4028 34552 4034 34564
rect 4157 34561 4169 34564
rect 4203 34561 4215 34595
rect 4157 34555 4215 34561
rect 5534 34552 5540 34604
rect 5592 34552 5598 34604
rect 3050 34524 3056 34536
rect 3011 34496 3056 34524
rect 3050 34484 3056 34496
rect 3108 34484 3114 34536
rect 5920 34533 5948 34632
rect 7650 34620 7656 34632
rect 7708 34620 7714 34672
rect 12066 34660 12072 34672
rect 9338 34632 12072 34660
rect 12066 34620 12072 34632
rect 12124 34620 12130 34672
rect 16942 34660 16948 34672
rect 13202 34632 16948 34660
rect 16942 34620 16948 34632
rect 17000 34620 17006 34672
rect 6549 34595 6607 34601
rect 6549 34561 6561 34595
rect 6595 34592 6607 34595
rect 7190 34592 7196 34604
rect 6595 34564 7196 34592
rect 6595 34561 6607 34564
rect 6549 34555 6607 34561
rect 7190 34552 7196 34564
rect 7248 34552 7254 34604
rect 10321 34595 10379 34601
rect 10321 34561 10333 34595
rect 10367 34561 10379 34595
rect 10321 34555 10379 34561
rect 5905 34527 5963 34533
rect 5905 34493 5917 34527
rect 5951 34493 5963 34527
rect 5905 34487 5963 34493
rect 6822 34484 6828 34536
rect 6880 34524 6886 34536
rect 7837 34527 7895 34533
rect 7837 34524 7849 34527
rect 6880 34496 7849 34524
rect 6880 34484 6886 34496
rect 7837 34493 7849 34496
rect 7883 34493 7895 34527
rect 8110 34524 8116 34536
rect 7837 34487 7895 34493
rect 7944 34496 8116 34524
rect 6546 34416 6552 34468
rect 6604 34456 6610 34468
rect 6733 34459 6791 34465
rect 6733 34456 6745 34459
rect 6604 34428 6745 34456
rect 6604 34416 6610 34428
rect 6733 34425 6745 34428
rect 6779 34425 6791 34459
rect 6733 34419 6791 34425
rect 4420 34391 4478 34397
rect 4420 34357 4432 34391
rect 4466 34388 4478 34391
rect 4890 34388 4896 34400
rect 4466 34360 4896 34388
rect 4466 34357 4478 34360
rect 4420 34351 4478 34357
rect 4890 34348 4896 34360
rect 4948 34388 4954 34400
rect 5166 34388 5172 34400
rect 4948 34360 5172 34388
rect 4948 34348 4954 34360
rect 5166 34348 5172 34360
rect 5224 34348 5230 34400
rect 6362 34348 6368 34400
rect 6420 34388 6426 34400
rect 7944 34388 7972 34496
rect 8110 34484 8116 34496
rect 8168 34484 8174 34536
rect 9122 34484 9128 34536
rect 9180 34524 9186 34536
rect 10336 34524 10364 34555
rect 10502 34552 10508 34604
rect 10560 34592 10566 34604
rect 10781 34595 10839 34601
rect 10781 34592 10793 34595
rect 10560 34564 10793 34592
rect 10560 34552 10566 34564
rect 10781 34561 10793 34564
rect 10827 34561 10839 34595
rect 10781 34555 10839 34561
rect 11054 34552 11060 34604
rect 11112 34592 11118 34604
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11112 34564 11713 34592
rect 11112 34552 11118 34564
rect 11701 34561 11713 34564
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34561 14243 34595
rect 14185 34555 14243 34561
rect 10870 34524 10876 34536
rect 9180 34496 10364 34524
rect 10831 34496 10876 34524
rect 9180 34484 9186 34496
rect 10870 34484 10876 34496
rect 10928 34484 10934 34536
rect 11330 34484 11336 34536
rect 11388 34524 11394 34536
rect 11974 34524 11980 34536
rect 11388 34496 11980 34524
rect 11388 34484 11394 34496
rect 11974 34484 11980 34496
rect 12032 34484 12038 34536
rect 12066 34484 12072 34536
rect 12124 34524 12130 34536
rect 12434 34524 12440 34536
rect 12124 34496 12440 34524
rect 12124 34484 12130 34496
rect 12434 34484 12440 34496
rect 12492 34484 12498 34536
rect 12526 34484 12532 34536
rect 12584 34524 12590 34536
rect 13449 34527 13507 34533
rect 13449 34524 13461 34527
rect 12584 34496 13461 34524
rect 12584 34484 12590 34496
rect 13449 34493 13461 34496
rect 13495 34493 13507 34527
rect 13449 34487 13507 34493
rect 13722 34484 13728 34536
rect 13780 34524 13786 34536
rect 14200 34524 14228 34555
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 14792 34564 14837 34592
rect 14792 34552 14798 34564
rect 15286 34552 15292 34604
rect 15344 34592 15350 34604
rect 15381 34595 15439 34601
rect 15381 34592 15393 34595
rect 15344 34564 15393 34592
rect 15344 34552 15350 34564
rect 15381 34561 15393 34564
rect 15427 34561 15439 34595
rect 15381 34555 15439 34561
rect 15470 34552 15476 34604
rect 15528 34592 15534 34604
rect 16025 34595 16083 34601
rect 15528 34564 15573 34592
rect 15528 34552 15534 34564
rect 16025 34561 16037 34595
rect 16071 34592 16083 34595
rect 16390 34592 16396 34604
rect 16071 34564 16396 34592
rect 16071 34561 16083 34564
rect 16025 34555 16083 34561
rect 16390 34552 16396 34564
rect 16448 34592 16454 34604
rect 16853 34595 16911 34601
rect 16853 34592 16865 34595
rect 16448 34564 16865 34592
rect 16448 34552 16454 34564
rect 16853 34561 16865 34564
rect 16899 34561 16911 34595
rect 17497 34595 17555 34601
rect 17497 34592 17509 34595
rect 16853 34555 16911 34561
rect 17052 34564 17509 34592
rect 16206 34524 16212 34536
rect 13780 34496 14136 34524
rect 14200 34496 16212 34524
rect 13780 34484 13786 34496
rect 11238 34456 11244 34468
rect 9508 34428 11244 34456
rect 6420 34360 7972 34388
rect 8100 34391 8158 34397
rect 6420 34348 6426 34360
rect 8100 34357 8112 34391
rect 8146 34388 8158 34391
rect 9508 34388 9536 34428
rect 11238 34416 11244 34428
rect 11296 34416 11302 34468
rect 14108 34456 14136 34496
rect 16206 34484 16212 34496
rect 16264 34484 16270 34536
rect 16942 34524 16948 34536
rect 16903 34496 16948 34524
rect 16942 34484 16948 34496
rect 17000 34484 17006 34536
rect 16117 34459 16175 34465
rect 16117 34456 16129 34459
rect 14108 34428 16129 34456
rect 16117 34425 16129 34428
rect 16163 34425 16175 34459
rect 16117 34419 16175 34425
rect 16482 34416 16488 34468
rect 16540 34456 16546 34468
rect 17052 34456 17080 34564
rect 17497 34561 17509 34564
rect 17543 34592 17555 34595
rect 18141 34595 18199 34601
rect 18141 34592 18153 34595
rect 17543 34564 18153 34592
rect 17543 34561 17555 34564
rect 17497 34555 17555 34561
rect 18141 34561 18153 34564
rect 18187 34592 18199 34595
rect 18598 34592 18604 34604
rect 18187 34564 18604 34592
rect 18187 34561 18199 34564
rect 18141 34555 18199 34561
rect 18598 34552 18604 34564
rect 18656 34552 18662 34604
rect 16540 34428 17080 34456
rect 16540 34416 16546 34428
rect 8146 34360 9536 34388
rect 8146 34357 8158 34360
rect 8100 34351 8158 34357
rect 9582 34348 9588 34400
rect 9640 34388 9646 34400
rect 10134 34388 10140 34400
rect 9640 34360 9685 34388
rect 10095 34360 10140 34388
rect 9640 34348 9646 34360
rect 10134 34348 10140 34360
rect 10192 34348 10198 34400
rect 12342 34348 12348 34400
rect 12400 34388 12406 34400
rect 14090 34388 14096 34400
rect 12400 34360 14096 34388
rect 12400 34348 12406 34360
rect 14090 34348 14096 34360
rect 14148 34348 14154 34400
rect 14185 34391 14243 34397
rect 14185 34357 14197 34391
rect 14231 34388 14243 34391
rect 14366 34388 14372 34400
rect 14231 34360 14372 34388
rect 14231 34357 14243 34360
rect 14185 34351 14243 34357
rect 14366 34348 14372 34360
rect 14424 34348 14430 34400
rect 15102 34348 15108 34400
rect 15160 34388 15166 34400
rect 16850 34388 16856 34400
rect 15160 34360 16856 34388
rect 15160 34348 15166 34360
rect 16850 34348 16856 34360
rect 16908 34348 16914 34400
rect 17586 34388 17592 34400
rect 17547 34360 17592 34388
rect 17586 34348 17592 34360
rect 17644 34348 17650 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 2869 34187 2927 34193
rect 2869 34153 2881 34187
rect 2915 34184 2927 34187
rect 6730 34184 6736 34196
rect 2915 34156 6736 34184
rect 2915 34153 2927 34156
rect 2869 34147 2927 34153
rect 6730 34144 6736 34156
rect 6788 34144 6794 34196
rect 7088 34187 7146 34193
rect 7088 34153 7100 34187
rect 7134 34184 7146 34187
rect 10778 34184 10784 34196
rect 7134 34156 10784 34184
rect 7134 34153 7146 34156
rect 7088 34147 7146 34153
rect 10778 34144 10784 34156
rect 10836 34184 10842 34196
rect 11780 34187 11838 34193
rect 10836 34156 11652 34184
rect 10836 34144 10842 34156
rect 8110 34076 8116 34128
rect 8168 34116 8174 34128
rect 8573 34119 8631 34125
rect 8573 34116 8585 34119
rect 8168 34088 8585 34116
rect 8168 34076 8174 34088
rect 8573 34085 8585 34088
rect 8619 34116 8631 34119
rect 10873 34119 10931 34125
rect 8619 34088 9260 34116
rect 8619 34085 8631 34088
rect 8573 34079 8631 34085
rect 3970 34048 3976 34060
rect 3931 34020 3976 34048
rect 3970 34008 3976 34020
rect 4028 34008 4034 34060
rect 4706 34008 4712 34060
rect 4764 34048 4770 34060
rect 5994 34048 6000 34060
rect 4764 34020 5856 34048
rect 5955 34020 6000 34048
rect 4764 34008 4770 34020
rect 1857 33983 1915 33989
rect 1857 33949 1869 33983
rect 1903 33980 1915 33983
rect 1946 33980 1952 33992
rect 1903 33952 1952 33980
rect 1903 33949 1915 33952
rect 1857 33943 1915 33949
rect 1946 33940 1952 33952
rect 2004 33940 2010 33992
rect 2777 33983 2835 33989
rect 2777 33949 2789 33983
rect 2823 33980 2835 33983
rect 3234 33980 3240 33992
rect 2823 33952 3240 33980
rect 2823 33949 2835 33952
rect 2777 33943 2835 33949
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 5828 33980 5856 34020
rect 5994 34008 6000 34020
rect 6052 34048 6058 34060
rect 6362 34048 6368 34060
rect 6052 34020 6368 34048
rect 6052 34008 6058 34020
rect 6362 34008 6368 34020
rect 6420 34008 6426 34060
rect 9125 34051 9183 34057
rect 9125 34048 9137 34051
rect 6840 34020 9137 34048
rect 6840 33992 6868 34020
rect 9125 34017 9137 34020
rect 9171 34017 9183 34051
rect 9232 34048 9260 34088
rect 10873 34085 10885 34119
rect 10919 34116 10931 34119
rect 11146 34116 11152 34128
rect 10919 34088 11152 34116
rect 10919 34085 10931 34088
rect 10873 34079 10931 34085
rect 11146 34076 11152 34088
rect 11204 34076 11210 34128
rect 9766 34048 9772 34060
rect 9232 34020 9772 34048
rect 9125 34011 9183 34017
rect 9766 34008 9772 34020
rect 9824 34008 9830 34060
rect 10042 34008 10048 34060
rect 10100 34048 10106 34060
rect 10962 34048 10968 34060
rect 10100 34020 10968 34048
rect 10100 34008 10106 34020
rect 10962 34008 10968 34020
rect 11020 34008 11026 34060
rect 11054 34008 11060 34060
rect 11112 34048 11118 34060
rect 11517 34051 11575 34057
rect 11517 34048 11529 34051
rect 11112 34020 11529 34048
rect 11112 34008 11118 34020
rect 11517 34017 11529 34020
rect 11563 34017 11575 34051
rect 11624 34048 11652 34156
rect 11780 34153 11792 34187
rect 11826 34184 11838 34187
rect 13262 34184 13268 34196
rect 11826 34156 13268 34184
rect 11826 34153 11838 34156
rect 11780 34147 11838 34153
rect 13262 34144 13268 34156
rect 13320 34144 13326 34196
rect 13538 34144 13544 34196
rect 13596 34184 13602 34196
rect 15102 34184 15108 34196
rect 13596 34156 15108 34184
rect 13596 34144 13602 34156
rect 15102 34144 15108 34156
rect 15160 34144 15166 34196
rect 15304 34156 17816 34184
rect 12342 34048 12348 34060
rect 11624 34020 12348 34048
rect 11517 34011 11575 34017
rect 12342 34008 12348 34020
rect 12400 34008 12406 34060
rect 14366 34048 14372 34060
rect 14327 34020 14372 34048
rect 14366 34008 14372 34020
rect 14424 34008 14430 34060
rect 15013 34051 15071 34057
rect 15013 34017 15025 34051
rect 15059 34048 15071 34051
rect 15304 34048 15332 34156
rect 15838 34076 15844 34128
rect 15896 34116 15902 34128
rect 16482 34116 16488 34128
rect 15896 34088 16488 34116
rect 15896 34076 15902 34088
rect 16482 34076 16488 34088
rect 16540 34116 16546 34128
rect 16761 34119 16819 34125
rect 16761 34116 16773 34119
rect 16540 34088 16773 34116
rect 16540 34076 16546 34088
rect 16761 34085 16773 34088
rect 16807 34085 16819 34119
rect 17788 34116 17816 34156
rect 17862 34144 17868 34196
rect 17920 34184 17926 34196
rect 18049 34187 18107 34193
rect 18049 34184 18061 34187
rect 17920 34156 18061 34184
rect 17920 34144 17926 34156
rect 18049 34153 18061 34156
rect 18095 34153 18107 34187
rect 18049 34147 18107 34153
rect 35897 34187 35955 34193
rect 35897 34153 35909 34187
rect 35943 34184 35955 34187
rect 37274 34184 37280 34196
rect 35943 34156 37280 34184
rect 35943 34153 35955 34156
rect 35897 34147 35955 34153
rect 37274 34144 37280 34156
rect 37332 34144 37338 34196
rect 19150 34116 19156 34128
rect 17788 34088 19156 34116
rect 16761 34079 16819 34085
rect 19150 34076 19156 34088
rect 19208 34076 19214 34128
rect 19242 34048 19248 34060
rect 15059 34020 15332 34048
rect 15396 34020 19248 34048
rect 15059 34017 15071 34020
rect 15013 34011 15071 34017
rect 6546 33980 6552 33992
rect 5828 33952 6552 33980
rect 6546 33940 6552 33952
rect 6604 33940 6610 33992
rect 6822 33980 6828 33992
rect 6783 33952 6828 33980
rect 6822 33940 6828 33952
rect 6880 33940 6886 33992
rect 8202 33940 8208 33992
rect 8260 33940 8266 33992
rect 10778 33980 10784 33992
rect 10534 33952 10784 33980
rect 10778 33940 10784 33952
rect 10836 33940 10842 33992
rect 13170 33940 13176 33992
rect 13228 33980 13234 33992
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 13228 33952 13553 33980
rect 13228 33940 13234 33952
rect 13541 33949 13553 33952
rect 13587 33949 13599 33983
rect 13541 33943 13599 33949
rect 1394 33872 1400 33924
rect 1452 33912 1458 33924
rect 2133 33915 2191 33921
rect 2133 33912 2145 33915
rect 1452 33884 2145 33912
rect 1452 33872 1458 33884
rect 2133 33881 2145 33884
rect 2179 33881 2191 33915
rect 2133 33875 2191 33881
rect 2148 33844 2176 33875
rect 4154 33872 4160 33924
rect 4212 33912 4218 33924
rect 4249 33915 4307 33921
rect 4249 33912 4261 33915
rect 4212 33884 4261 33912
rect 4212 33872 4218 33884
rect 4249 33881 4261 33884
rect 4295 33881 4307 33915
rect 6638 33912 6644 33924
rect 5474 33884 6644 33912
rect 4249 33875 4307 33881
rect 6638 33872 6644 33884
rect 6696 33872 6702 33924
rect 8478 33872 8484 33924
rect 8536 33912 8542 33924
rect 9030 33912 9036 33924
rect 8536 33884 9036 33912
rect 8536 33872 8542 33884
rect 9030 33872 9036 33884
rect 9088 33912 9094 33924
rect 9401 33915 9459 33921
rect 9401 33912 9413 33915
rect 9088 33884 9413 33912
rect 9088 33872 9094 33884
rect 9401 33881 9413 33884
rect 9447 33881 9459 33915
rect 11882 33912 11888 33924
rect 9401 33875 9459 33881
rect 10704 33884 11888 33912
rect 10704 33844 10732 33884
rect 11882 33872 11888 33884
rect 11940 33872 11946 33924
rect 13446 33912 13452 33924
rect 13018 33884 13452 33912
rect 13446 33872 13452 33884
rect 13504 33872 13510 33924
rect 13998 33872 14004 33924
rect 14056 33912 14062 33924
rect 14461 33915 14519 33921
rect 14461 33912 14473 33915
rect 14056 33884 14473 33912
rect 14056 33872 14062 33884
rect 14461 33881 14473 33884
rect 14507 33881 14519 33915
rect 14461 33875 14519 33881
rect 2148 33816 10732 33844
rect 12710 33804 12716 33856
rect 12768 33844 12774 33856
rect 15396 33844 15424 34020
rect 19242 34008 19248 34020
rect 19300 34008 19306 34060
rect 15657 33983 15715 33989
rect 15657 33949 15669 33983
rect 15703 33980 15715 33983
rect 16022 33980 16028 33992
rect 15703 33952 16028 33980
rect 15703 33949 15715 33952
rect 15657 33943 15715 33949
rect 16022 33940 16028 33952
rect 16080 33940 16086 33992
rect 17310 33980 17316 33992
rect 17271 33952 17316 33980
rect 17310 33940 17316 33952
rect 17368 33940 17374 33992
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 18598 33980 18604 33992
rect 18559 33952 18604 33980
rect 17957 33943 18015 33949
rect 16206 33912 16212 33924
rect 16167 33884 16212 33912
rect 16206 33872 16212 33884
rect 16264 33872 16270 33924
rect 16301 33915 16359 33921
rect 16301 33881 16313 33915
rect 16347 33881 16359 33915
rect 16301 33875 16359 33881
rect 12768 33816 15424 33844
rect 15473 33847 15531 33853
rect 12768 33804 12774 33816
rect 15473 33813 15485 33847
rect 15519 33844 15531 33847
rect 16316 33844 16344 33875
rect 16390 33872 16396 33924
rect 16448 33912 16454 33924
rect 17972 33912 18000 33943
rect 18598 33940 18604 33952
rect 18656 33940 18662 33992
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 36081 33983 36139 33989
rect 36081 33980 36093 33983
rect 34572 33952 36093 33980
rect 34572 33940 34578 33952
rect 36081 33949 36093 33952
rect 36127 33949 36139 33983
rect 36081 33943 36139 33949
rect 16448 33884 18000 33912
rect 16448 33872 16454 33884
rect 15519 33816 16344 33844
rect 17405 33847 17463 33853
rect 15519 33813 15531 33816
rect 15473 33807 15531 33813
rect 17405 33813 17417 33847
rect 17451 33844 17463 33847
rect 17862 33844 17868 33856
rect 17451 33816 17868 33844
rect 17451 33813 17463 33816
rect 17405 33807 17463 33813
rect 17862 33804 17868 33816
rect 17920 33804 17926 33856
rect 18690 33844 18696 33856
rect 18651 33816 18696 33844
rect 18690 33804 18696 33816
rect 18748 33804 18754 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 2130 33600 2136 33652
rect 2188 33640 2194 33652
rect 3789 33643 3847 33649
rect 2188 33612 2774 33640
rect 2188 33600 2194 33612
rect 2314 33572 2320 33584
rect 2275 33544 2320 33572
rect 2314 33532 2320 33544
rect 2372 33532 2378 33584
rect 2746 33572 2774 33612
rect 3789 33609 3801 33643
rect 3835 33640 3847 33643
rect 5442 33640 5448 33652
rect 3835 33612 5448 33640
rect 3835 33609 3847 33612
rect 3789 33603 3847 33609
rect 5442 33600 5448 33612
rect 5500 33600 5506 33652
rect 5997 33643 6055 33649
rect 5997 33609 6009 33643
rect 6043 33640 6055 33643
rect 6914 33640 6920 33652
rect 6043 33612 6920 33640
rect 6043 33609 6055 33612
rect 5997 33603 6055 33609
rect 6914 33600 6920 33612
rect 6972 33640 6978 33652
rect 7742 33640 7748 33652
rect 6972 33612 7748 33640
rect 6972 33600 6978 33612
rect 7742 33600 7748 33612
rect 7800 33600 7806 33652
rect 7834 33600 7840 33652
rect 7892 33640 7898 33652
rect 9398 33640 9404 33652
rect 7892 33612 9404 33640
rect 7892 33600 7898 33612
rect 9398 33600 9404 33612
rect 9456 33600 9462 33652
rect 11514 33640 11520 33652
rect 9646 33612 11520 33640
rect 2746 33544 2806 33572
rect 1578 33464 1584 33516
rect 1636 33504 1642 33516
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1636 33476 2053 33504
rect 1636 33464 1642 33476
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 3970 33464 3976 33516
rect 4028 33504 4034 33516
rect 4249 33507 4307 33513
rect 4249 33504 4261 33507
rect 4028 33476 4261 33504
rect 4028 33464 4034 33476
rect 4249 33473 4261 33476
rect 4295 33473 4307 33507
rect 6546 33504 6552 33516
rect 4249 33467 4307 33473
rect 4264 33300 4292 33467
rect 4522 33436 4528 33448
rect 4483 33408 4528 33436
rect 4522 33396 4528 33408
rect 4580 33396 4586 33448
rect 5644 33368 5672 33490
rect 6507 33476 6552 33504
rect 6546 33464 6552 33476
rect 6604 33464 6610 33516
rect 7098 33464 7104 33516
rect 7156 33504 7162 33516
rect 7193 33507 7251 33513
rect 7193 33504 7205 33507
rect 7156 33476 7205 33504
rect 7156 33464 7162 33476
rect 7193 33473 7205 33476
rect 7239 33473 7251 33507
rect 7193 33467 7251 33473
rect 7285 33507 7343 33513
rect 7285 33473 7297 33507
rect 7331 33504 7343 33507
rect 7374 33504 7380 33516
rect 7331 33476 7380 33504
rect 7331 33473 7343 33476
rect 7285 33467 7343 33473
rect 7374 33464 7380 33476
rect 7432 33464 7438 33516
rect 9646 33504 9674 33612
rect 11514 33600 11520 33612
rect 11572 33600 11578 33652
rect 12618 33600 12624 33652
rect 12676 33640 12682 33652
rect 13998 33640 14004 33652
rect 12676 33612 13860 33640
rect 13959 33612 14004 33640
rect 12676 33600 12682 33612
rect 9861 33575 9919 33581
rect 9861 33541 9873 33575
rect 9907 33572 9919 33575
rect 10042 33572 10048 33584
rect 9907 33544 10048 33572
rect 9907 33541 9919 33544
rect 9861 33535 9919 33541
rect 10042 33532 10048 33544
rect 10100 33532 10106 33584
rect 13832 33572 13860 33612
rect 13998 33600 14004 33612
rect 14056 33600 14062 33652
rect 14090 33600 14096 33652
rect 14148 33640 14154 33652
rect 15838 33640 15844 33652
rect 14148 33612 15844 33640
rect 14148 33600 14154 33612
rect 15838 33600 15844 33612
rect 15896 33600 15902 33652
rect 16022 33640 16028 33652
rect 15983 33612 16028 33640
rect 16022 33600 16028 33612
rect 16080 33600 16086 33652
rect 16206 33600 16212 33652
rect 16264 33640 16270 33652
rect 16853 33643 16911 33649
rect 16853 33640 16865 33643
rect 16264 33612 16865 33640
rect 16264 33600 16270 33612
rect 16853 33609 16865 33612
rect 16899 33609 16911 33643
rect 16853 33603 16911 33609
rect 17310 33572 17316 33584
rect 13832 33544 17316 33572
rect 9246 33476 9674 33504
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10410 33504 10416 33516
rect 10367 33476 10416 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10962 33504 10968 33516
rect 10923 33476 10968 33504
rect 10962 33464 10968 33476
rect 11020 33464 11026 33516
rect 11054 33464 11060 33516
rect 11112 33504 11118 33516
rect 11701 33507 11759 33513
rect 11701 33504 11713 33507
rect 11112 33476 11713 33504
rect 11112 33464 11118 33476
rect 11701 33473 11713 33476
rect 11747 33473 11759 33507
rect 13906 33504 13912 33516
rect 13110 33476 13768 33504
rect 13867 33476 13912 33504
rect 11701 33467 11759 33473
rect 6822 33396 6828 33448
rect 6880 33436 6886 33448
rect 7837 33439 7895 33445
rect 7837 33436 7849 33439
rect 6880 33408 7849 33436
rect 6880 33396 6886 33408
rect 7837 33405 7849 33408
rect 7883 33405 7895 33439
rect 7837 33399 7895 33405
rect 8113 33439 8171 33445
rect 8113 33405 8125 33439
rect 8159 33436 8171 33439
rect 9306 33436 9312 33448
rect 8159 33408 9312 33436
rect 8159 33405 8171 33408
rect 8113 33399 8171 33405
rect 9306 33396 9312 33408
rect 9364 33396 9370 33448
rect 9398 33396 9404 33448
rect 9456 33436 9462 33448
rect 11514 33436 11520 33448
rect 9456 33408 11520 33436
rect 9456 33396 9462 33408
rect 11514 33396 11520 33408
rect 11572 33396 11578 33448
rect 11977 33439 12035 33445
rect 11977 33436 11989 33439
rect 11624 33408 11989 33436
rect 11057 33371 11115 33377
rect 11057 33368 11069 33371
rect 5644 33340 7972 33368
rect 5534 33300 5540 33312
rect 4264 33272 5540 33300
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 6730 33300 6736 33312
rect 6687 33272 6736 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 6730 33260 6736 33272
rect 6788 33260 6794 33312
rect 7944 33300 7972 33340
rect 9646 33340 11069 33368
rect 9646 33300 9674 33340
rect 11057 33337 11069 33340
rect 11103 33337 11115 33371
rect 11057 33331 11115 33337
rect 11146 33328 11152 33380
rect 11204 33368 11210 33380
rect 11624 33368 11652 33408
rect 11977 33405 11989 33408
rect 12023 33405 12035 33439
rect 11977 33399 12035 33405
rect 12066 33396 12072 33448
rect 12124 33436 12130 33448
rect 12710 33436 12716 33448
rect 12124 33408 12716 33436
rect 12124 33396 12130 33408
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 12986 33396 12992 33448
rect 13044 33436 13050 33448
rect 13449 33439 13507 33445
rect 13449 33436 13461 33439
rect 13044 33408 13461 33436
rect 13044 33396 13050 33408
rect 13449 33405 13461 33408
rect 13495 33405 13507 33439
rect 13740 33436 13768 33476
rect 13906 33464 13912 33476
rect 13964 33464 13970 33516
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 14553 33507 14611 33513
rect 14553 33504 14565 33507
rect 14056 33476 14565 33504
rect 14056 33464 14062 33476
rect 14553 33473 14565 33476
rect 14599 33504 14611 33507
rect 14734 33504 14740 33516
rect 14599 33476 14740 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 14734 33464 14740 33476
rect 14792 33464 14798 33516
rect 15194 33504 15200 33516
rect 15155 33476 15200 33504
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 16224 33513 16252 33544
rect 17310 33532 17316 33544
rect 17368 33532 17374 33584
rect 17862 33572 17868 33584
rect 17823 33544 17868 33572
rect 17862 33532 17868 33544
rect 17920 33532 17926 33584
rect 16209 33507 16267 33513
rect 16209 33473 16221 33507
rect 16255 33473 16267 33507
rect 16209 33467 16267 33473
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33504 20223 33507
rect 20346 33504 20352 33516
rect 20211 33476 20352 33504
rect 20211 33473 20223 33476
rect 20165 33467 20223 33473
rect 20346 33464 20352 33476
rect 20404 33464 20410 33516
rect 31478 33504 31484 33516
rect 31439 33476 31484 33504
rect 31478 33464 31484 33476
rect 31536 33464 31542 33516
rect 37918 33464 37924 33516
rect 37976 33504 37982 33516
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 37976 33476 38025 33504
rect 37976 33464 37982 33476
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 17586 33436 17592 33448
rect 13740 33408 17592 33436
rect 13449 33399 13507 33405
rect 17586 33396 17592 33408
rect 17644 33396 17650 33448
rect 17773 33439 17831 33445
rect 17773 33405 17785 33439
rect 17819 33436 17831 33439
rect 19978 33436 19984 33448
rect 17819 33408 19984 33436
rect 17819 33405 17831 33408
rect 17773 33399 17831 33405
rect 19978 33396 19984 33408
rect 20036 33396 20042 33448
rect 11204 33340 11652 33368
rect 11204 33328 11210 33340
rect 13538 33328 13544 33380
rect 13596 33368 13602 33380
rect 14645 33371 14703 33377
rect 14645 33368 14657 33371
rect 13596 33340 14657 33368
rect 13596 33328 13602 33340
rect 14645 33337 14657 33340
rect 14691 33337 14703 33371
rect 14645 33331 14703 33337
rect 15194 33328 15200 33380
rect 15252 33368 15258 33380
rect 16206 33368 16212 33380
rect 15252 33340 16212 33368
rect 15252 33328 15258 33340
rect 16206 33328 16212 33340
rect 16264 33328 16270 33380
rect 16482 33328 16488 33380
rect 16540 33368 16546 33380
rect 18325 33371 18383 33377
rect 18325 33368 18337 33371
rect 16540 33340 18337 33368
rect 16540 33328 16546 33340
rect 18325 33337 18337 33340
rect 18371 33337 18383 33371
rect 21266 33368 21272 33380
rect 18325 33331 18383 33337
rect 18432 33340 21272 33368
rect 7944 33272 9674 33300
rect 9766 33260 9772 33312
rect 9824 33300 9830 33312
rect 10413 33303 10471 33309
rect 10413 33300 10425 33303
rect 9824 33272 10425 33300
rect 9824 33260 9830 33272
rect 10413 33269 10425 33272
rect 10459 33269 10471 33303
rect 10413 33263 10471 33269
rect 10594 33260 10600 33312
rect 10652 33300 10658 33312
rect 12066 33300 12072 33312
rect 10652 33272 12072 33300
rect 10652 33260 10658 33272
rect 12066 33260 12072 33272
rect 12124 33260 12130 33312
rect 14090 33260 14096 33312
rect 14148 33300 14154 33312
rect 15289 33303 15347 33309
rect 15289 33300 15301 33303
rect 14148 33272 15301 33300
rect 14148 33260 14154 33272
rect 15289 33269 15301 33272
rect 15335 33269 15347 33303
rect 15289 33263 15347 33269
rect 15838 33260 15844 33312
rect 15896 33300 15902 33312
rect 18432 33300 18460 33340
rect 21266 33328 21272 33340
rect 21324 33328 21330 33380
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 20254 33300 20260 33312
rect 15896 33272 18460 33300
rect 20215 33272 20260 33300
rect 15896 33260 15902 33272
rect 20254 33260 20260 33272
rect 20312 33260 20318 33312
rect 28994 33260 29000 33312
rect 29052 33300 29058 33312
rect 31573 33303 31631 33309
rect 31573 33300 31585 33303
rect 29052 33272 31585 33300
rect 29052 33260 29058 33272
rect 31573 33269 31585 33272
rect 31619 33269 31631 33303
rect 31573 33263 31631 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1762 33096 1768 33108
rect 1723 33068 1768 33096
rect 1762 33056 1768 33068
rect 1820 33056 1826 33108
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 4065 33099 4123 33105
rect 4065 33096 4077 33099
rect 3200 33068 4077 33096
rect 3200 33056 3206 33068
rect 4065 33065 4077 33068
rect 4111 33065 4123 33099
rect 4065 33059 4123 33065
rect 6812 33099 6870 33105
rect 6812 33065 6824 33099
rect 6858 33096 6870 33099
rect 6858 33068 8616 33096
rect 6858 33065 6870 33068
rect 6812 33059 6870 33065
rect 8588 33028 8616 33068
rect 8938 33056 8944 33108
rect 8996 33096 9002 33108
rect 13722 33096 13728 33108
rect 8996 33068 13728 33096
rect 8996 33056 9002 33068
rect 13722 33056 13728 33068
rect 13780 33056 13786 33108
rect 13814 33056 13820 33108
rect 13872 33096 13878 33108
rect 18690 33096 18696 33108
rect 13872 33068 18696 33096
rect 13872 33056 13878 33068
rect 18690 33056 18696 33068
rect 18748 33056 18754 33108
rect 9582 33028 9588 33040
rect 8588 33000 9588 33028
rect 9582 32988 9588 33000
rect 9640 32988 9646 33040
rect 9674 32988 9680 33040
rect 9732 33028 9738 33040
rect 11146 33028 11152 33040
rect 9732 33000 11152 33028
rect 9732 32988 9738 33000
rect 11146 32988 11152 33000
rect 11204 32988 11210 33040
rect 15470 33028 15476 33040
rect 12544 33000 15476 33028
rect 2958 32920 2964 32972
rect 3016 32960 3022 32972
rect 3326 32960 3332 32972
rect 3016 32932 3332 32960
rect 3016 32920 3022 32932
rect 3326 32920 3332 32932
rect 3384 32960 3390 32972
rect 4982 32960 4988 32972
rect 3384 32932 4988 32960
rect 3384 32920 3390 32932
rect 1486 32852 1492 32904
rect 1544 32892 1550 32904
rect 1581 32895 1639 32901
rect 1581 32892 1593 32895
rect 1544 32864 1593 32892
rect 1544 32852 1550 32864
rect 1581 32861 1593 32864
rect 1627 32861 1639 32895
rect 2314 32892 2320 32904
rect 2275 32864 2320 32892
rect 1581 32855 1639 32861
rect 2314 32852 2320 32864
rect 2372 32892 2378 32904
rect 3142 32892 3148 32904
rect 2372 32864 2774 32892
rect 3103 32864 3148 32892
rect 2372 32852 2378 32864
rect 2746 32824 2774 32864
rect 3142 32852 3148 32864
rect 3200 32852 3206 32904
rect 3234 32852 3240 32904
rect 3292 32892 3298 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3292 32864 3985 32892
rect 3292 32852 3298 32864
rect 3973 32861 3985 32864
rect 4019 32892 4031 32895
rect 4246 32892 4252 32904
rect 4019 32864 4252 32892
rect 4019 32861 4031 32864
rect 3973 32855 4031 32861
rect 4246 32852 4252 32864
rect 4304 32852 4310 32904
rect 4632 32901 4660 32932
rect 4982 32920 4988 32932
rect 5040 32960 5046 32972
rect 5040 32932 5396 32960
rect 5040 32920 5046 32932
rect 4617 32895 4675 32901
rect 4617 32861 4629 32895
rect 4663 32861 4675 32895
rect 4617 32855 4675 32861
rect 4706 32852 4712 32904
rect 4764 32892 4770 32904
rect 4890 32892 4896 32904
rect 4764 32864 4896 32892
rect 4764 32852 4770 32864
rect 4890 32852 4896 32864
rect 4948 32892 4954 32904
rect 5261 32895 5319 32901
rect 5261 32892 5273 32895
rect 4948 32864 5273 32892
rect 4948 32852 4954 32864
rect 5261 32861 5273 32864
rect 5307 32861 5319 32895
rect 5368 32892 5396 32932
rect 5534 32920 5540 32972
rect 5592 32960 5598 32972
rect 6546 32960 6552 32972
rect 5592 32932 6552 32960
rect 5592 32920 5598 32932
rect 6546 32920 6552 32932
rect 6604 32960 6610 32972
rect 6822 32960 6828 32972
rect 6604 32932 6828 32960
rect 6604 32920 6610 32932
rect 6822 32920 6828 32932
rect 6880 32920 6886 32972
rect 7374 32920 7380 32972
rect 7432 32960 7438 32972
rect 7432 32932 9168 32960
rect 7432 32920 7438 32932
rect 5905 32895 5963 32901
rect 5905 32892 5917 32895
rect 5368 32864 5917 32892
rect 5261 32855 5319 32861
rect 5905 32861 5917 32864
rect 5951 32892 5963 32895
rect 8938 32892 8944 32904
rect 5951 32864 6592 32892
rect 7958 32864 8944 32892
rect 5951 32861 5963 32864
rect 5905 32855 5963 32861
rect 6454 32824 6460 32836
rect 2746 32796 6460 32824
rect 6454 32784 6460 32796
rect 6512 32784 6518 32836
rect 2406 32756 2412 32768
rect 2367 32728 2412 32756
rect 2406 32716 2412 32728
rect 2464 32716 2470 32768
rect 2961 32759 3019 32765
rect 2961 32725 2973 32759
rect 3007 32756 3019 32759
rect 3786 32756 3792 32768
rect 3007 32728 3792 32756
rect 3007 32725 3019 32728
rect 2961 32719 3019 32725
rect 3786 32716 3792 32728
rect 3844 32716 3850 32768
rect 4706 32756 4712 32768
rect 4667 32728 4712 32756
rect 4706 32716 4712 32728
rect 4764 32716 4770 32768
rect 5353 32759 5411 32765
rect 5353 32725 5365 32759
rect 5399 32756 5411 32759
rect 5718 32756 5724 32768
rect 5399 32728 5724 32756
rect 5399 32725 5411 32728
rect 5353 32719 5411 32725
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 5997 32759 6055 32765
rect 5997 32725 6009 32759
rect 6043 32756 6055 32759
rect 6086 32756 6092 32768
rect 6043 32728 6092 32756
rect 6043 32725 6055 32728
rect 5997 32719 6055 32725
rect 6086 32716 6092 32728
rect 6144 32716 6150 32768
rect 6564 32756 6592 32864
rect 8938 32852 8944 32864
rect 8996 32852 9002 32904
rect 9140 32901 9168 32932
rect 9214 32920 9220 32972
rect 9272 32960 9278 32972
rect 9272 32932 10640 32960
rect 9272 32920 9278 32932
rect 9125 32895 9183 32901
rect 9125 32861 9137 32895
rect 9171 32892 9183 32895
rect 9398 32892 9404 32904
rect 9171 32864 9404 32892
rect 9171 32861 9183 32864
rect 9125 32855 9183 32861
rect 9398 32852 9404 32864
rect 9456 32852 9462 32904
rect 9769 32895 9827 32901
rect 9769 32861 9781 32895
rect 9815 32892 9827 32895
rect 9950 32892 9956 32904
rect 9815 32864 9956 32892
rect 9815 32861 9827 32864
rect 9769 32855 9827 32861
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 10410 32892 10416 32904
rect 10371 32864 10416 32892
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 8478 32784 8484 32836
rect 8536 32824 8542 32836
rect 8573 32827 8631 32833
rect 8573 32824 8585 32827
rect 8536 32796 8585 32824
rect 8536 32784 8542 32796
rect 8573 32793 8585 32796
rect 8619 32793 8631 32827
rect 10505 32827 10563 32833
rect 10505 32824 10517 32827
rect 8573 32787 8631 32793
rect 8956 32796 10517 32824
rect 7466 32756 7472 32768
rect 6564 32728 7472 32756
rect 7466 32716 7472 32728
rect 7524 32716 7530 32768
rect 8110 32716 8116 32768
rect 8168 32756 8174 32768
rect 8956 32756 8984 32796
rect 10505 32793 10517 32796
rect 10551 32793 10563 32827
rect 10612 32824 10640 32932
rect 11054 32920 11060 32972
rect 11112 32960 11118 32972
rect 11241 32963 11299 32969
rect 11241 32960 11253 32963
rect 11112 32932 11253 32960
rect 11112 32920 11118 32932
rect 11241 32929 11253 32932
rect 11287 32929 11299 32963
rect 11241 32923 11299 32929
rect 11514 32920 11520 32972
rect 11572 32960 11578 32972
rect 12544 32960 12572 33000
rect 15470 32988 15476 33000
rect 15528 32988 15534 33040
rect 16666 32988 16672 33040
rect 16724 33028 16730 33040
rect 17589 33031 17647 33037
rect 17589 33028 17601 33031
rect 16724 33000 17601 33028
rect 16724 32988 16730 33000
rect 17589 32997 17601 33000
rect 17635 32997 17647 33031
rect 17589 32991 17647 32997
rect 21082 32988 21088 33040
rect 21140 33028 21146 33040
rect 24857 33031 24915 33037
rect 24857 33028 24869 33031
rect 21140 33000 24869 33028
rect 21140 32988 21146 33000
rect 24857 32997 24869 33000
rect 24903 32997 24915 33031
rect 24857 32991 24915 32997
rect 16942 32960 16948 32972
rect 11572 32932 12572 32960
rect 12636 32932 16948 32960
rect 11572 32920 11578 32932
rect 12636 32878 12664 32932
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 22066 32932 22692 32960
rect 13633 32895 13691 32901
rect 13633 32861 13645 32895
rect 13679 32892 13691 32895
rect 13998 32892 14004 32904
rect 13679 32864 14004 32892
rect 13679 32861 13691 32864
rect 13633 32855 13691 32861
rect 13998 32852 14004 32864
rect 14056 32852 14062 32904
rect 14553 32895 14611 32901
rect 14553 32861 14565 32895
rect 14599 32861 14611 32895
rect 15010 32892 15016 32904
rect 14971 32864 15016 32892
rect 14553 32855 14611 32861
rect 11517 32827 11575 32833
rect 11517 32824 11529 32827
rect 10612 32796 11529 32824
rect 10505 32787 10563 32793
rect 11517 32793 11529 32796
rect 11563 32793 11575 32827
rect 11517 32787 11575 32793
rect 12912 32796 13492 32824
rect 9214 32756 9220 32768
rect 8168 32728 8984 32756
rect 9175 32728 9220 32756
rect 8168 32716 8174 32728
rect 9214 32716 9220 32728
rect 9272 32716 9278 32768
rect 9398 32716 9404 32768
rect 9456 32756 9462 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 9456 32728 9873 32756
rect 9456 32716 9462 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9861 32719 9919 32725
rect 10226 32716 10232 32768
rect 10284 32756 10290 32768
rect 12912 32756 12940 32796
rect 10284 32728 12940 32756
rect 12989 32759 13047 32765
rect 10284 32716 10290 32728
rect 12989 32725 13001 32759
rect 13035 32756 13047 32759
rect 13262 32756 13268 32768
rect 13035 32728 13268 32756
rect 13035 32725 13047 32728
rect 12989 32719 13047 32725
rect 13262 32716 13268 32728
rect 13320 32716 13326 32768
rect 13464 32765 13492 32796
rect 13906 32784 13912 32836
rect 13964 32824 13970 32836
rect 14568 32824 14596 32855
rect 15010 32852 15016 32864
rect 15068 32852 15074 32904
rect 16209 32895 16267 32901
rect 16209 32861 16221 32895
rect 16255 32861 16267 32895
rect 16209 32855 16267 32861
rect 13964 32796 14596 32824
rect 13964 32784 13970 32796
rect 14826 32784 14832 32836
rect 14884 32824 14890 32836
rect 15930 32824 15936 32836
rect 14884 32796 15936 32824
rect 14884 32784 14890 32796
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 16224 32824 16252 32855
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 16853 32895 16911 32901
rect 16853 32892 16865 32895
rect 16540 32864 16865 32892
rect 16540 32852 16546 32864
rect 16853 32861 16865 32864
rect 16899 32861 16911 32895
rect 17494 32892 17500 32904
rect 17455 32864 17500 32892
rect 16853 32855 16911 32861
rect 17494 32852 17500 32864
rect 17552 32852 17558 32904
rect 19242 32852 19248 32904
rect 19300 32892 19306 32904
rect 21545 32895 21603 32901
rect 21545 32892 21557 32895
rect 19300 32864 21557 32892
rect 19300 32852 19306 32864
rect 21545 32861 21557 32864
rect 21591 32892 21603 32895
rect 22066 32892 22094 32932
rect 22664 32901 22692 32932
rect 21591 32864 22094 32892
rect 22189 32895 22247 32901
rect 21591 32861 21603 32864
rect 21545 32855 21603 32861
rect 22189 32861 22201 32895
rect 22235 32861 22247 32895
rect 22189 32855 22247 32861
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32861 22707 32895
rect 22649 32855 22707 32861
rect 24765 32895 24823 32901
rect 24765 32861 24777 32895
rect 24811 32892 24823 32895
rect 29730 32892 29736 32904
rect 24811 32864 29736 32892
rect 24811 32861 24823 32864
rect 24765 32855 24823 32861
rect 18138 32824 18144 32836
rect 16224 32796 18144 32824
rect 18138 32784 18144 32796
rect 18196 32784 18202 32836
rect 22204 32824 22232 32855
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32892 32367 32895
rect 35894 32892 35900 32904
rect 32355 32864 35900 32892
rect 32355 32861 32367 32864
rect 32309 32855 32367 32861
rect 35894 32852 35900 32864
rect 35952 32852 35958 32904
rect 21376 32796 22232 32824
rect 13449 32759 13507 32765
rect 13449 32725 13461 32759
rect 13495 32725 13507 32759
rect 14366 32756 14372 32768
rect 14327 32728 14372 32756
rect 13449 32719 13507 32725
rect 14366 32716 14372 32728
rect 14424 32716 14430 32768
rect 14458 32716 14464 32768
rect 14516 32756 14522 32768
rect 15105 32759 15163 32765
rect 15105 32756 15117 32759
rect 14516 32728 15117 32756
rect 14516 32716 14522 32728
rect 15105 32725 15117 32728
rect 15151 32725 15163 32759
rect 15105 32719 15163 32725
rect 16022 32716 16028 32768
rect 16080 32756 16086 32768
rect 16301 32759 16359 32765
rect 16301 32756 16313 32759
rect 16080 32728 16313 32756
rect 16080 32716 16086 32728
rect 16301 32725 16313 32728
rect 16347 32725 16359 32759
rect 16942 32756 16948 32768
rect 16903 32728 16948 32756
rect 16301 32719 16359 32725
rect 16942 32716 16948 32728
rect 17000 32716 17006 32768
rect 21376 32765 21404 32796
rect 21361 32759 21419 32765
rect 21361 32725 21373 32759
rect 21407 32725 21419 32759
rect 21361 32719 21419 32725
rect 22005 32759 22063 32765
rect 22005 32725 22017 32759
rect 22051 32756 22063 32759
rect 22186 32756 22192 32768
rect 22051 32728 22192 32756
rect 22051 32725 22063 32728
rect 22005 32719 22063 32725
rect 22186 32716 22192 32728
rect 22244 32716 22250 32768
rect 22554 32716 22560 32768
rect 22612 32756 22618 32768
rect 22741 32759 22799 32765
rect 22741 32756 22753 32759
rect 22612 32728 22753 32756
rect 22612 32716 22618 32728
rect 22741 32725 22753 32728
rect 22787 32725 22799 32759
rect 22741 32719 22799 32725
rect 31754 32716 31760 32768
rect 31812 32756 31818 32768
rect 32401 32759 32459 32765
rect 32401 32756 32413 32759
rect 31812 32728 32413 32756
rect 31812 32716 31818 32728
rect 32401 32725 32413 32728
rect 32447 32725 32459 32759
rect 32401 32719 32459 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 4246 32512 4252 32564
rect 4304 32552 4310 32564
rect 5810 32552 5816 32564
rect 4304 32524 5816 32552
rect 4304 32512 4310 32524
rect 2866 32484 2872 32496
rect 2056 32456 2872 32484
rect 2056 32425 2084 32456
rect 2866 32444 2872 32456
rect 2924 32444 2930 32496
rect 4798 32484 4804 32496
rect 4186 32456 4804 32484
rect 4798 32444 4804 32456
rect 4856 32444 4862 32496
rect 2041 32419 2099 32425
rect 2041 32385 2053 32419
rect 2087 32385 2099 32419
rect 4982 32416 4988 32428
rect 4943 32388 4988 32416
rect 2041 32379 2099 32385
rect 4982 32376 4988 32388
rect 5040 32376 5046 32428
rect 5644 32425 5672 32524
rect 5810 32512 5816 32524
rect 5868 32552 5874 32564
rect 5868 32524 6224 32552
rect 5868 32512 5874 32524
rect 6196 32484 6224 32524
rect 6454 32512 6460 32564
rect 6512 32552 6518 32564
rect 10594 32552 10600 32564
rect 6512 32524 10600 32552
rect 6512 32512 6518 32524
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 10686 32512 10692 32564
rect 10744 32552 10750 32564
rect 10965 32555 11023 32561
rect 10965 32552 10977 32555
rect 10744 32524 10977 32552
rect 10744 32512 10750 32524
rect 10965 32521 10977 32524
rect 11011 32521 11023 32555
rect 10965 32515 11023 32521
rect 12158 32512 12164 32564
rect 12216 32552 12222 32564
rect 12216 32524 13952 32552
rect 12216 32512 12222 32524
rect 7098 32484 7104 32496
rect 6196 32456 7104 32484
rect 7098 32444 7104 32456
rect 7156 32444 7162 32496
rect 7650 32444 7656 32496
rect 7708 32484 7714 32496
rect 8021 32487 8079 32493
rect 8021 32484 8033 32487
rect 7708 32456 8033 32484
rect 7708 32444 7714 32456
rect 8021 32453 8033 32456
rect 8067 32453 8079 32487
rect 11514 32484 11520 32496
rect 9246 32456 11520 32484
rect 8021 32447 8079 32453
rect 11514 32444 11520 32456
rect 11572 32444 11578 32496
rect 13814 32484 13820 32496
rect 13202 32456 13820 32484
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 5629 32419 5687 32425
rect 5629 32385 5641 32419
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 5721 32419 5779 32425
rect 5721 32385 5733 32419
rect 5767 32416 5779 32419
rect 5994 32416 6000 32428
rect 5767 32388 6000 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 5994 32376 6000 32388
rect 6052 32376 6058 32428
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32416 6607 32419
rect 6822 32416 6828 32428
rect 6595 32388 6828 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 6822 32376 6828 32388
rect 6880 32376 6886 32428
rect 9674 32376 9680 32428
rect 9732 32416 9738 32428
rect 9769 32419 9827 32425
rect 9769 32416 9781 32419
rect 9732 32388 9781 32416
rect 9732 32376 9738 32388
rect 9769 32385 9781 32388
rect 9815 32385 9827 32419
rect 9769 32379 9827 32385
rect 9950 32376 9956 32428
rect 10008 32416 10014 32428
rect 10413 32419 10471 32425
rect 10413 32416 10425 32419
rect 10008 32388 10425 32416
rect 10008 32376 10014 32388
rect 10413 32385 10425 32388
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 10778 32376 10784 32428
rect 10836 32416 10842 32428
rect 10873 32419 10931 32425
rect 10873 32416 10885 32419
rect 10836 32388 10885 32416
rect 10836 32376 10842 32388
rect 10873 32385 10885 32388
rect 10919 32416 10931 32419
rect 10962 32416 10968 32428
rect 10919 32388 10968 32416
rect 10919 32385 10931 32388
rect 10873 32379 10931 32385
rect 10962 32376 10968 32388
rect 11020 32376 11026 32428
rect 11054 32376 11060 32428
rect 11112 32416 11118 32428
rect 13924 32425 13952 32524
rect 13998 32512 14004 32564
rect 14056 32552 14062 32564
rect 14056 32524 14101 32552
rect 14056 32512 14062 32524
rect 14182 32512 14188 32564
rect 14240 32552 14246 32564
rect 14458 32552 14464 32564
rect 14240 32524 14464 32552
rect 14240 32512 14246 32524
rect 14458 32512 14464 32524
rect 14516 32512 14522 32564
rect 14642 32512 14648 32564
rect 14700 32552 14706 32564
rect 15933 32555 15991 32561
rect 15933 32552 15945 32555
rect 14700 32524 15945 32552
rect 14700 32512 14706 32524
rect 15933 32521 15945 32524
rect 15979 32521 15991 32555
rect 15933 32515 15991 32521
rect 16206 32512 16212 32564
rect 16264 32552 16270 32564
rect 16390 32552 16396 32564
rect 16264 32524 16396 32552
rect 16264 32512 16270 32524
rect 16390 32512 16396 32524
rect 16448 32552 16454 32564
rect 16448 32524 17172 32552
rect 16448 32512 16454 32524
rect 14366 32444 14372 32496
rect 14424 32484 14430 32496
rect 14424 32456 17080 32484
rect 14424 32444 14430 32456
rect 11701 32419 11759 32425
rect 11701 32416 11713 32419
rect 11112 32388 11713 32416
rect 11112 32376 11118 32388
rect 11701 32385 11713 32388
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32385 13967 32419
rect 14553 32419 14611 32425
rect 14553 32416 14565 32419
rect 13909 32379 13967 32385
rect 14292 32388 14565 32416
rect 1578 32308 1584 32360
rect 1636 32348 1642 32360
rect 2682 32348 2688 32360
rect 1636 32320 2688 32348
rect 1636 32308 1642 32320
rect 2682 32308 2688 32320
rect 2740 32308 2746 32360
rect 2961 32351 3019 32357
rect 2961 32317 2973 32351
rect 3007 32348 3019 32351
rect 3007 32320 6592 32348
rect 3007 32317 3019 32320
rect 2961 32311 3019 32317
rect 4433 32283 4491 32289
rect 4433 32249 4445 32283
rect 4479 32280 4491 32283
rect 5166 32280 5172 32292
rect 4479 32252 5172 32280
rect 4479 32249 4491 32252
rect 4433 32243 4491 32249
rect 5166 32240 5172 32252
rect 5224 32240 5230 32292
rect 5626 32240 5632 32292
rect 5684 32280 5690 32292
rect 5902 32280 5908 32292
rect 5684 32252 5908 32280
rect 5684 32240 5690 32252
rect 5902 32240 5908 32252
rect 5960 32240 5966 32292
rect 6564 32280 6592 32320
rect 6638 32308 6644 32360
rect 6696 32348 6702 32360
rect 7745 32351 7803 32357
rect 7745 32348 7757 32351
rect 6696 32320 7757 32348
rect 6696 32308 6702 32320
rect 7745 32317 7757 32320
rect 7791 32317 7803 32351
rect 7745 32311 7803 32317
rect 8386 32308 8392 32360
rect 8444 32348 8450 32360
rect 9692 32348 9720 32376
rect 8444 32320 9720 32348
rect 8444 32308 8450 32320
rect 10594 32308 10600 32360
rect 10652 32348 10658 32360
rect 14292 32348 14320 32388
rect 14553 32385 14565 32388
rect 14599 32416 14611 32419
rect 15010 32416 15016 32428
rect 14599 32388 15016 32416
rect 14599 32385 14611 32388
rect 14553 32379 14611 32385
rect 15010 32376 15016 32388
rect 15068 32376 15074 32428
rect 15197 32419 15255 32425
rect 15197 32385 15209 32419
rect 15243 32416 15255 32419
rect 15378 32416 15384 32428
rect 15243 32388 15384 32416
rect 15243 32385 15255 32388
rect 15197 32379 15255 32385
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 15838 32416 15844 32428
rect 15799 32388 15844 32416
rect 15838 32376 15844 32388
rect 15896 32376 15902 32428
rect 17052 32425 17080 32456
rect 17037 32419 17095 32425
rect 17037 32385 17049 32419
rect 17083 32385 17095 32419
rect 17144 32416 17172 32524
rect 19518 32512 19524 32564
rect 19576 32552 19582 32564
rect 20622 32552 20628 32564
rect 19576 32524 20628 32552
rect 19576 32512 19582 32524
rect 20622 32512 20628 32524
rect 20680 32512 20686 32564
rect 34333 32555 34391 32561
rect 34333 32552 34345 32555
rect 26206 32524 34345 32552
rect 17497 32419 17555 32425
rect 17497 32416 17509 32419
rect 17144 32388 17509 32416
rect 17037 32379 17095 32385
rect 17497 32385 17509 32388
rect 17543 32385 17555 32419
rect 17497 32379 17555 32385
rect 17770 32376 17776 32428
rect 17828 32416 17834 32428
rect 18877 32419 18935 32425
rect 18877 32416 18889 32419
rect 17828 32388 18889 32416
rect 17828 32376 17834 32388
rect 18877 32385 18889 32388
rect 18923 32385 18935 32419
rect 18877 32379 18935 32385
rect 19521 32419 19579 32425
rect 19521 32385 19533 32419
rect 19567 32385 19579 32419
rect 22554 32416 22560 32428
rect 22515 32388 22560 32416
rect 19521 32379 19579 32385
rect 10652 32320 14320 32348
rect 10652 32308 10658 32320
rect 14366 32308 14372 32360
rect 14424 32348 14430 32360
rect 14645 32351 14703 32357
rect 14645 32348 14657 32351
rect 14424 32320 14657 32348
rect 14424 32308 14430 32320
rect 14645 32317 14657 32320
rect 14691 32317 14703 32351
rect 17589 32351 17647 32357
rect 17589 32348 17601 32351
rect 14645 32311 14703 32317
rect 14752 32320 17601 32348
rect 6914 32280 6920 32292
rect 6564 32252 6920 32280
rect 6914 32240 6920 32252
rect 6972 32240 6978 32292
rect 9030 32240 9036 32292
rect 9088 32280 9094 32292
rect 9398 32280 9404 32292
rect 9088 32252 9404 32280
rect 9088 32240 9094 32252
rect 9398 32240 9404 32252
rect 9456 32240 9462 32292
rect 14182 32240 14188 32292
rect 14240 32280 14246 32292
rect 14752 32280 14780 32320
rect 17589 32317 17601 32320
rect 17635 32317 17647 32351
rect 17589 32311 17647 32317
rect 18046 32308 18052 32360
rect 18104 32348 18110 32360
rect 19536 32348 19564 32379
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 23934 32416 23940 32428
rect 23895 32388 23940 32416
rect 23934 32376 23940 32388
rect 23992 32376 23998 32428
rect 18104 32320 19564 32348
rect 22373 32351 22431 32357
rect 18104 32308 18110 32320
rect 22373 32317 22385 32351
rect 22419 32348 22431 32351
rect 26206 32348 26234 32524
rect 34333 32521 34345 32524
rect 34379 32521 34391 32555
rect 38105 32555 38163 32561
rect 38105 32552 38117 32555
rect 34333 32515 34391 32521
rect 35866 32524 38117 32552
rect 33689 32487 33747 32493
rect 22419 32320 26234 32348
rect 28368 32456 33640 32484
rect 22419 32317 22431 32320
rect 22373 32311 22431 32317
rect 14240 32252 14780 32280
rect 15120 32252 15424 32280
rect 14240 32240 14246 32252
rect 2133 32215 2191 32221
rect 2133 32181 2145 32215
rect 2179 32212 2191 32215
rect 2590 32212 2596 32224
rect 2179 32184 2596 32212
rect 2179 32181 2191 32184
rect 2133 32175 2191 32181
rect 2590 32172 2596 32184
rect 2648 32172 2654 32224
rect 3510 32172 3516 32224
rect 3568 32212 3574 32224
rect 5077 32215 5135 32221
rect 5077 32212 5089 32215
rect 3568 32184 5089 32212
rect 3568 32172 3574 32184
rect 5077 32181 5089 32184
rect 5123 32181 5135 32215
rect 5077 32175 5135 32181
rect 6641 32215 6699 32221
rect 6641 32181 6653 32215
rect 6687 32212 6699 32215
rect 9674 32212 9680 32224
rect 6687 32184 9680 32212
rect 6687 32181 6699 32184
rect 6641 32175 6699 32181
rect 9674 32172 9680 32184
rect 9732 32172 9738 32224
rect 10226 32212 10232 32224
rect 10187 32184 10232 32212
rect 10226 32172 10232 32184
rect 10284 32172 10290 32224
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10778 32212 10784 32224
rect 10468 32184 10784 32212
rect 10468 32172 10474 32184
rect 10778 32172 10784 32184
rect 10836 32172 10842 32224
rect 11790 32172 11796 32224
rect 11848 32212 11854 32224
rect 11964 32215 12022 32221
rect 11964 32212 11976 32215
rect 11848 32184 11976 32212
rect 11848 32172 11854 32184
rect 11964 32181 11976 32184
rect 12010 32212 12022 32215
rect 12526 32212 12532 32224
rect 12010 32184 12532 32212
rect 12010 32181 12022 32184
rect 11964 32175 12022 32181
rect 12526 32172 12532 32184
rect 12584 32172 12590 32224
rect 12710 32172 12716 32224
rect 12768 32212 12774 32224
rect 13449 32215 13507 32221
rect 13449 32212 13461 32215
rect 12768 32184 13461 32212
rect 12768 32172 12774 32184
rect 13449 32181 13461 32184
rect 13495 32212 13507 32215
rect 14550 32212 14556 32224
rect 13495 32184 14556 32212
rect 13495 32181 13507 32184
rect 13449 32175 13507 32181
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 14734 32172 14740 32224
rect 14792 32212 14798 32224
rect 15120 32212 15148 32252
rect 14792 32184 15148 32212
rect 14792 32172 14798 32184
rect 15194 32172 15200 32224
rect 15252 32212 15258 32224
rect 15289 32215 15347 32221
rect 15289 32212 15301 32215
rect 15252 32184 15301 32212
rect 15252 32172 15258 32184
rect 15289 32181 15301 32184
rect 15335 32181 15347 32215
rect 15396 32212 15424 32252
rect 15470 32240 15476 32292
rect 15528 32280 15534 32292
rect 16482 32280 16488 32292
rect 15528 32252 16488 32280
rect 15528 32240 15534 32252
rect 16482 32240 16488 32252
rect 16540 32240 16546 32292
rect 16853 32283 16911 32289
rect 16853 32249 16865 32283
rect 16899 32280 16911 32283
rect 18598 32280 18604 32292
rect 16899 32252 18604 32280
rect 16899 32249 16911 32252
rect 16853 32243 16911 32249
rect 18598 32240 18604 32252
rect 18656 32240 18662 32292
rect 22738 32240 22744 32292
rect 22796 32280 22802 32292
rect 24029 32283 24087 32289
rect 24029 32280 24041 32283
rect 22796 32252 24041 32280
rect 22796 32240 22802 32252
rect 24029 32249 24041 32252
rect 24075 32249 24087 32283
rect 24029 32243 24087 32249
rect 26142 32240 26148 32292
rect 26200 32280 26206 32292
rect 28368 32280 28396 32456
rect 28445 32419 28503 32425
rect 28445 32385 28457 32419
rect 28491 32416 28503 32419
rect 32214 32416 32220 32428
rect 28491 32388 32220 32416
rect 28491 32385 28503 32388
rect 28445 32379 28503 32385
rect 32214 32376 32220 32388
rect 32272 32376 32278 32428
rect 33612 32425 33640 32456
rect 33689 32453 33701 32487
rect 33735 32484 33747 32487
rect 34514 32484 34520 32496
rect 33735 32456 34520 32484
rect 33735 32453 33747 32456
rect 33689 32447 33747 32453
rect 34514 32444 34520 32456
rect 34572 32444 34578 32496
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32385 32367 32419
rect 32309 32379 32367 32385
rect 33597 32419 33655 32425
rect 33597 32385 33609 32419
rect 33643 32385 33655 32419
rect 33597 32379 33655 32385
rect 34241 32419 34299 32425
rect 34241 32385 34253 32419
rect 34287 32416 34299 32419
rect 35866 32416 35894 32524
rect 38105 32521 38117 32524
rect 38151 32521 38163 32555
rect 38105 32515 38163 32521
rect 38286 32416 38292 32428
rect 34287 32388 35894 32416
rect 38247 32388 38292 32416
rect 34287 32385 34299 32388
rect 34241 32379 34299 32385
rect 32324 32348 32352 32379
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 35986 32348 35992 32360
rect 32324 32320 35992 32348
rect 35986 32308 35992 32320
rect 36044 32308 36050 32360
rect 26200 32252 28396 32280
rect 26200 32240 26206 32252
rect 17494 32212 17500 32224
rect 15396 32184 17500 32212
rect 15289 32175 15347 32181
rect 17494 32172 17500 32184
rect 17552 32172 17558 32224
rect 18693 32215 18751 32221
rect 18693 32181 18705 32215
rect 18739 32212 18751 32215
rect 18874 32212 18880 32224
rect 18739 32184 18880 32212
rect 18739 32181 18751 32184
rect 18693 32175 18751 32181
rect 18874 32172 18880 32184
rect 18932 32172 18938 32224
rect 19613 32215 19671 32221
rect 19613 32181 19625 32215
rect 19659 32212 19671 32215
rect 20346 32212 20352 32224
rect 19659 32184 20352 32212
rect 19659 32181 19671 32184
rect 19613 32175 19671 32181
rect 20346 32172 20352 32184
rect 20404 32172 20410 32224
rect 22830 32212 22836 32224
rect 22791 32184 22836 32212
rect 22830 32172 22836 32184
rect 22888 32172 22894 32224
rect 26326 32172 26332 32224
rect 26384 32212 26390 32224
rect 28537 32215 28595 32221
rect 28537 32212 28549 32215
rect 26384 32184 28549 32212
rect 26384 32172 26390 32184
rect 28537 32181 28549 32184
rect 28583 32181 28595 32215
rect 32398 32212 32404 32224
rect 32359 32184 32404 32212
rect 28537 32175 28595 32181
rect 32398 32172 32404 32184
rect 32456 32172 32462 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 3329 32011 3387 32017
rect 3329 31977 3341 32011
rect 3375 32008 3387 32011
rect 3970 32008 3976 32020
rect 3375 31980 3976 32008
rect 3375 31977 3387 31980
rect 3329 31971 3387 31977
rect 3970 31968 3976 31980
rect 4028 31968 4034 32020
rect 5534 32008 5540 32020
rect 4908 31980 5540 32008
rect 1578 31872 1584 31884
rect 1539 31844 1584 31872
rect 1578 31832 1584 31844
rect 1636 31832 1642 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 4908 31881 4936 31980
rect 5534 31968 5540 31980
rect 5592 31968 5598 32020
rect 7484 31980 8064 32008
rect 7484 31940 7512 31980
rect 7208 31912 7512 31940
rect 8036 31940 8064 31980
rect 8110 31968 8116 32020
rect 8168 32008 8174 32020
rect 15013 32011 15071 32017
rect 15013 32008 15025 32011
rect 8168 31980 15025 32008
rect 8168 31968 8174 31980
rect 15013 31977 15025 31980
rect 15059 31977 15071 32011
rect 15654 32008 15660 32020
rect 15615 31980 15660 32008
rect 15013 31971 15071 31977
rect 15654 31968 15660 31980
rect 15712 31968 15718 32020
rect 15930 31968 15936 32020
rect 15988 32008 15994 32020
rect 16301 32011 16359 32017
rect 16301 32008 16313 32011
rect 15988 31980 16313 32008
rect 15988 31968 15994 31980
rect 16301 31977 16313 31980
rect 16347 31977 16359 32011
rect 16301 31971 16359 31977
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 16945 32011 17003 32017
rect 16945 32008 16957 32011
rect 16908 31980 16957 32008
rect 16908 31968 16914 31980
rect 16945 31977 16957 31980
rect 16991 31977 17003 32011
rect 16945 31971 17003 31977
rect 19978 31968 19984 32020
rect 20036 32008 20042 32020
rect 22373 32011 22431 32017
rect 22373 32008 22385 32011
rect 20036 31980 22385 32008
rect 20036 31968 20042 31980
rect 22373 31977 22385 31980
rect 22419 32008 22431 32011
rect 22830 32008 22836 32020
rect 22419 31980 22836 32008
rect 22419 31977 22431 31980
rect 22373 31971 22431 31977
rect 22830 31968 22836 31980
rect 22888 31968 22894 32020
rect 8570 31940 8576 31952
rect 8036 31912 8576 31940
rect 4893 31875 4951 31881
rect 4893 31841 4905 31875
rect 4939 31841 4951 31875
rect 4893 31835 4951 31841
rect 5169 31875 5227 31881
rect 5169 31841 5181 31875
rect 5215 31872 5227 31875
rect 7208 31872 7236 31912
rect 8570 31900 8576 31912
rect 8628 31900 8634 31952
rect 9490 31900 9496 31952
rect 9548 31940 9554 31952
rect 9585 31943 9643 31949
rect 9585 31940 9597 31943
rect 9548 31912 9597 31940
rect 9548 31900 9554 31912
rect 9585 31909 9597 31912
rect 9631 31909 9643 31943
rect 13630 31940 13636 31952
rect 13591 31912 13636 31940
rect 9585 31903 9643 31909
rect 13630 31900 13636 31912
rect 13688 31900 13694 31952
rect 18693 31943 18751 31949
rect 18693 31909 18705 31943
rect 18739 31940 18751 31943
rect 20070 31940 20076 31952
rect 18739 31912 20076 31940
rect 18739 31909 18751 31912
rect 18693 31903 18751 31909
rect 20070 31900 20076 31912
rect 20128 31900 20134 31952
rect 21082 31940 21088 31952
rect 20180 31912 21088 31940
rect 5215 31844 7236 31872
rect 5215 31841 5227 31844
rect 5169 31835 5227 31841
rect 7282 31832 7288 31884
rect 7340 31872 7346 31884
rect 7469 31875 7527 31881
rect 7469 31872 7481 31875
rect 7340 31844 7481 31872
rect 7340 31832 7346 31844
rect 7469 31841 7481 31844
rect 7515 31841 7527 31875
rect 7469 31835 7527 31841
rect 7650 31832 7656 31884
rect 7708 31872 7714 31884
rect 10686 31872 10692 31884
rect 7708 31844 10692 31872
rect 7708 31832 7714 31844
rect 10686 31832 10692 31844
rect 10744 31832 10750 31884
rect 11054 31832 11060 31884
rect 11112 31872 11118 31884
rect 11333 31875 11391 31881
rect 11333 31872 11345 31875
rect 11112 31844 11345 31872
rect 11112 31832 11118 31844
rect 11333 31841 11345 31844
rect 11379 31872 11391 31875
rect 11698 31872 11704 31884
rect 11379 31844 11704 31872
rect 11379 31841 11391 31844
rect 11333 31835 11391 31841
rect 11698 31832 11704 31844
rect 11756 31832 11762 31884
rect 14366 31872 14372 31884
rect 14327 31844 14372 31872
rect 14366 31832 14372 31844
rect 14424 31832 14430 31884
rect 19334 31832 19340 31884
rect 19392 31872 19398 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 19392 31844 19625 31872
rect 19392 31832 19398 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 20180 31872 20208 31912
rect 21082 31900 21088 31912
rect 21140 31900 21146 31952
rect 20530 31872 20536 31884
rect 19613 31835 19671 31841
rect 20088 31844 20208 31872
rect 20491 31844 20536 31872
rect 3970 31804 3976 31816
rect 3931 31776 3976 31804
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31804 4123 31807
rect 4798 31804 4804 31816
rect 4111 31776 4804 31804
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 4798 31764 4804 31776
rect 4856 31764 4862 31816
rect 6914 31804 6920 31816
rect 6875 31776 6920 31804
rect 6914 31764 6920 31776
rect 6972 31804 6978 31816
rect 6972 31776 7328 31804
rect 6972 31764 6978 31776
rect 4614 31736 4620 31748
rect 3082 31708 4620 31736
rect 4614 31696 4620 31708
rect 4672 31696 4678 31748
rect 6178 31696 6184 31748
rect 6236 31696 6242 31748
rect 7300 31736 7328 31776
rect 7374 31764 7380 31816
rect 7432 31804 7438 31816
rect 7432 31776 7477 31804
rect 7432 31764 7438 31776
rect 8662 31764 8668 31816
rect 8720 31804 8726 31816
rect 9769 31807 9827 31813
rect 8720 31776 9674 31804
rect 8720 31764 8726 31776
rect 7466 31736 7472 31748
rect 7300 31708 7472 31736
rect 7466 31696 7472 31708
rect 7524 31696 7530 31748
rect 7926 31696 7932 31748
rect 7984 31736 7990 31748
rect 8389 31739 8447 31745
rect 8389 31736 8401 31739
rect 7984 31708 8401 31736
rect 7984 31696 7990 31708
rect 8389 31705 8401 31708
rect 8435 31705 8447 31739
rect 8389 31699 8447 31705
rect 8846 31696 8852 31748
rect 8904 31736 8910 31748
rect 9398 31736 9404 31748
rect 8904 31708 9404 31736
rect 8904 31696 8910 31708
rect 9398 31696 9404 31708
rect 9456 31696 9462 31748
rect 9646 31736 9674 31776
rect 9769 31773 9781 31807
rect 9815 31804 9827 31807
rect 9858 31804 9864 31816
rect 9815 31776 9864 31804
rect 9815 31773 9827 31776
rect 9769 31767 9827 31773
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 10134 31764 10140 31816
rect 10192 31804 10198 31816
rect 10229 31807 10287 31813
rect 10229 31804 10241 31807
rect 10192 31776 10241 31804
rect 10192 31764 10198 31776
rect 10229 31773 10241 31776
rect 10275 31773 10287 31807
rect 10229 31767 10287 31773
rect 10321 31807 10379 31813
rect 10321 31773 10333 31807
rect 10367 31804 10379 31807
rect 10410 31804 10416 31816
rect 10367 31776 10416 31804
rect 10367 31773 10379 31776
rect 10321 31767 10379 31773
rect 10410 31764 10416 31776
rect 10468 31764 10474 31816
rect 13538 31804 13544 31816
rect 13499 31776 13544 31804
rect 13538 31764 13544 31776
rect 13596 31764 13602 31816
rect 13814 31764 13820 31816
rect 13872 31804 13878 31816
rect 13998 31804 14004 31816
rect 13872 31776 14004 31804
rect 13872 31764 13878 31776
rect 13998 31764 14004 31776
rect 14056 31804 14062 31816
rect 14277 31807 14335 31813
rect 14277 31804 14289 31807
rect 14056 31776 14289 31804
rect 14056 31764 14062 31776
rect 14277 31773 14289 31776
rect 14323 31804 14335 31807
rect 14921 31807 14979 31813
rect 14921 31804 14933 31807
rect 14323 31776 14933 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 14921 31773 14933 31776
rect 14967 31773 14979 31807
rect 14921 31767 14979 31773
rect 15010 31764 15016 31816
rect 15068 31804 15074 31816
rect 15565 31807 15623 31813
rect 15565 31804 15577 31807
rect 15068 31776 15577 31804
rect 15068 31764 15074 31776
rect 15565 31773 15577 31776
rect 15611 31804 15623 31807
rect 16209 31807 16267 31813
rect 16209 31804 16221 31807
rect 15611 31776 16221 31804
rect 15611 31773 15623 31776
rect 15565 31767 15623 31773
rect 16209 31773 16221 31776
rect 16255 31804 16267 31807
rect 16853 31807 16911 31813
rect 16853 31804 16865 31807
rect 16255 31776 16865 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 16853 31773 16865 31776
rect 16899 31773 16911 31807
rect 18874 31804 18880 31816
rect 18835 31776 18880 31804
rect 16853 31767 16911 31773
rect 18874 31764 18880 31776
rect 18932 31764 18938 31816
rect 19518 31804 19524 31816
rect 19479 31776 19524 31804
rect 19518 31764 19524 31776
rect 19576 31764 19582 31816
rect 10778 31736 10784 31748
rect 9646 31708 10784 31736
rect 10778 31696 10784 31708
rect 10836 31696 10842 31748
rect 11606 31736 11612 31748
rect 11567 31708 11612 31736
rect 11606 31696 11612 31708
rect 11664 31696 11670 31748
rect 12066 31696 12072 31748
rect 12124 31696 12130 31748
rect 12986 31696 12992 31748
rect 13044 31736 13050 31748
rect 20088 31736 20116 31844
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 22186 31872 22192 31884
rect 22147 31844 22192 31872
rect 22186 31832 22192 31844
rect 22244 31832 22250 31884
rect 32398 31872 32404 31884
rect 23308 31844 32404 31872
rect 21818 31764 21824 31816
rect 21876 31804 21882 31816
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21876 31776 22017 31804
rect 21876 31764 21882 31776
rect 22005 31773 22017 31776
rect 22051 31804 22063 31807
rect 23308 31804 23336 31844
rect 32398 31832 32404 31844
rect 32456 31832 32462 31884
rect 25130 31804 25136 31816
rect 22051 31776 23336 31804
rect 25091 31776 25136 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 25130 31764 25136 31776
rect 25188 31764 25194 31816
rect 25498 31764 25504 31816
rect 25556 31804 25562 31816
rect 25777 31807 25835 31813
rect 25777 31804 25789 31807
rect 25556 31776 25789 31804
rect 25556 31764 25562 31776
rect 25777 31773 25789 31776
rect 25823 31773 25835 31807
rect 25777 31767 25835 31773
rect 20257 31739 20315 31745
rect 20257 31736 20269 31739
rect 13044 31708 13216 31736
rect 20088 31708 20269 31736
rect 13044 31696 13050 31708
rect 7098 31628 7104 31680
rect 7156 31668 7162 31680
rect 10962 31668 10968 31680
rect 7156 31640 10968 31668
rect 7156 31628 7162 31640
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 12618 31628 12624 31680
rect 12676 31668 12682 31680
rect 13081 31671 13139 31677
rect 13081 31668 13093 31671
rect 12676 31640 13093 31668
rect 12676 31628 12682 31640
rect 13081 31637 13093 31640
rect 13127 31637 13139 31671
rect 13188 31668 13216 31708
rect 20257 31705 20269 31708
rect 20303 31705 20315 31739
rect 20257 31699 20315 31705
rect 20346 31696 20352 31748
rect 20404 31736 20410 31748
rect 20404 31708 20449 31736
rect 20404 31696 20410 31708
rect 24854 31668 24860 31680
rect 13188 31640 24860 31668
rect 13081 31631 13139 31637
rect 24854 31628 24860 31640
rect 24912 31628 24918 31680
rect 25222 31668 25228 31680
rect 25183 31640 25228 31668
rect 25222 31628 25228 31640
rect 25280 31628 25286 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1946 31464 1952 31476
rect 1907 31436 1952 31464
rect 1946 31424 1952 31436
rect 2004 31424 2010 31476
rect 3050 31424 3056 31476
rect 3108 31464 3114 31476
rect 3108 31436 4844 31464
rect 3108 31424 3114 31436
rect 4522 31396 4528 31408
rect 4186 31368 4528 31396
rect 4522 31356 4528 31368
rect 4580 31356 4586 31408
rect 1854 31328 1860 31340
rect 1815 31300 1860 31328
rect 1854 31288 1860 31300
rect 1912 31288 1918 31340
rect 2682 31328 2688 31340
rect 2643 31300 2688 31328
rect 2682 31288 2688 31300
rect 2740 31288 2746 31340
rect 4816 31328 4844 31436
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 5721 31467 5779 31473
rect 5721 31464 5733 31467
rect 5684 31436 5733 31464
rect 5684 31424 5690 31436
rect 5721 31433 5733 31436
rect 5767 31433 5779 31467
rect 5721 31427 5779 31433
rect 6822 31424 6828 31476
rect 6880 31464 6886 31476
rect 9122 31464 9128 31476
rect 6880 31436 9128 31464
rect 6880 31424 6886 31436
rect 9122 31424 9128 31436
rect 9180 31424 9186 31476
rect 9214 31424 9220 31476
rect 9272 31464 9278 31476
rect 9398 31464 9404 31476
rect 9272 31436 9404 31464
rect 9272 31424 9278 31436
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 10870 31464 10876 31476
rect 9784 31436 10876 31464
rect 9784 31396 9812 31436
rect 10870 31424 10876 31436
rect 10928 31424 10934 31476
rect 10962 31424 10968 31476
rect 11020 31464 11026 31476
rect 13078 31464 13084 31476
rect 11020 31436 13084 31464
rect 11020 31424 11026 31436
rect 13078 31424 13084 31436
rect 13136 31424 13142 31476
rect 14185 31467 14243 31473
rect 14185 31433 14197 31467
rect 14231 31464 14243 31467
rect 14274 31464 14280 31476
rect 14231 31436 14280 31464
rect 14231 31433 14243 31436
rect 14185 31427 14243 31433
rect 14274 31424 14280 31436
rect 14332 31424 14338 31476
rect 16945 31467 17003 31473
rect 16945 31433 16957 31467
rect 16991 31464 17003 31467
rect 17126 31464 17132 31476
rect 16991 31436 17132 31464
rect 16991 31433 17003 31436
rect 16945 31427 17003 31433
rect 17126 31424 17132 31436
rect 17184 31424 17190 31476
rect 19978 31464 19984 31476
rect 18524 31436 19984 31464
rect 8050 31368 9812 31396
rect 10778 31356 10784 31408
rect 10836 31396 10842 31408
rect 18524 31396 18552 31436
rect 19978 31424 19984 31436
rect 20036 31424 20042 31476
rect 31754 31464 31760 31476
rect 22066 31436 31760 31464
rect 10836 31368 14136 31396
rect 10836 31356 10842 31368
rect 4816 31326 4936 31328
rect 4982 31326 4988 31340
rect 4816 31300 4988 31326
rect 4908 31298 4988 31300
rect 4982 31288 4988 31298
rect 5040 31328 5046 31340
rect 5626 31328 5632 31340
rect 5040 31300 5133 31328
rect 5539 31300 5632 31328
rect 5040 31288 5046 31300
rect 5626 31288 5632 31300
rect 5684 31328 5690 31340
rect 5810 31328 5816 31340
rect 5684 31300 5816 31328
rect 5684 31288 5690 31300
rect 5810 31288 5816 31300
rect 5868 31288 5874 31340
rect 10962 31328 10968 31340
rect 10534 31300 10968 31328
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11974 31288 11980 31340
rect 12032 31328 12038 31340
rect 12345 31331 12403 31337
rect 12345 31328 12357 31331
rect 12032 31300 12357 31328
rect 12032 31288 12038 31300
rect 12345 31297 12357 31300
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 12526 31288 12532 31340
rect 12584 31328 12590 31340
rect 12805 31331 12863 31337
rect 12805 31328 12817 31331
rect 12584 31300 12817 31328
rect 12584 31288 12590 31300
rect 12805 31297 12817 31300
rect 12851 31328 12863 31331
rect 12851 31300 13400 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 2961 31263 3019 31269
rect 2961 31229 2973 31263
rect 3007 31260 3019 31263
rect 5902 31260 5908 31272
rect 3007 31232 5908 31260
rect 3007 31229 3019 31232
rect 2961 31223 3019 31229
rect 5902 31220 5908 31232
rect 5960 31220 5966 31272
rect 6546 31260 6552 31272
rect 6507 31232 6552 31260
rect 6546 31220 6552 31232
rect 6604 31220 6610 31272
rect 6822 31260 6828 31272
rect 6783 31232 6828 31260
rect 6822 31220 6828 31232
rect 6880 31220 6886 31272
rect 7190 31220 7196 31272
rect 7248 31260 7254 31272
rect 7248 31232 8708 31260
rect 7248 31220 7254 31232
rect 4433 31127 4491 31133
rect 4433 31093 4445 31127
rect 4479 31124 4491 31127
rect 4614 31124 4620 31136
rect 4479 31096 4620 31124
rect 4479 31093 4491 31096
rect 4433 31087 4491 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 5077 31127 5135 31133
rect 5077 31093 5089 31127
rect 5123 31124 5135 31127
rect 6914 31124 6920 31136
rect 5123 31096 6920 31124
rect 5123 31093 5135 31096
rect 5077 31087 5135 31093
rect 6914 31084 6920 31096
rect 6972 31084 6978 31136
rect 8297 31127 8355 31133
rect 8297 31093 8309 31127
rect 8343 31124 8355 31127
rect 8478 31124 8484 31136
rect 8343 31096 8484 31124
rect 8343 31093 8355 31096
rect 8297 31087 8355 31093
rect 8478 31084 8484 31096
rect 8536 31084 8542 31136
rect 8680 31124 8708 31232
rect 8754 31220 8760 31272
rect 8812 31260 8818 31272
rect 9125 31263 9183 31269
rect 9125 31260 9137 31263
rect 8812 31232 9137 31260
rect 8812 31220 8818 31232
rect 9125 31229 9137 31232
rect 9171 31229 9183 31263
rect 9398 31260 9404 31272
rect 9311 31232 9404 31260
rect 9125 31223 9183 31229
rect 9398 31220 9404 31232
rect 9456 31260 9462 31272
rect 9456 31232 10456 31260
rect 9456 31220 9462 31232
rect 10428 31192 10456 31232
rect 10594 31220 10600 31272
rect 10652 31260 10658 31272
rect 11149 31263 11207 31269
rect 11149 31260 11161 31263
rect 10652 31232 11161 31260
rect 10652 31220 10658 31232
rect 11149 31229 11161 31232
rect 11195 31229 11207 31263
rect 12894 31260 12900 31272
rect 11149 31223 11207 31229
rect 11256 31232 12900 31260
rect 11256 31192 11284 31232
rect 12894 31220 12900 31232
rect 12952 31220 12958 31272
rect 13372 31260 13400 31300
rect 13446 31288 13452 31340
rect 13504 31328 13510 31340
rect 14108 31337 14136 31368
rect 16868 31368 18552 31396
rect 14093 31331 14151 31337
rect 13504 31300 14044 31328
rect 13504 31288 13510 31300
rect 13814 31260 13820 31272
rect 13372 31232 13820 31260
rect 13814 31220 13820 31232
rect 13872 31220 13878 31272
rect 14016 31260 14044 31300
rect 14093 31297 14105 31331
rect 14139 31328 14151 31331
rect 14274 31328 14280 31340
rect 14139 31300 14280 31328
rect 14139 31297 14151 31300
rect 14093 31291 14151 31297
rect 14274 31288 14280 31300
rect 14332 31288 14338 31340
rect 14734 31328 14740 31340
rect 14695 31300 14740 31328
rect 14734 31288 14740 31300
rect 14792 31288 14798 31340
rect 15378 31328 15384 31340
rect 15291 31300 15384 31328
rect 15378 31288 15384 31300
rect 15436 31288 15442 31340
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16390 31328 16396 31340
rect 16071 31300 16396 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16390 31288 16396 31300
rect 16448 31288 16454 31340
rect 16868 31337 16896 31368
rect 18598 31356 18604 31408
rect 18656 31396 18662 31408
rect 18877 31399 18935 31405
rect 18877 31396 18889 31399
rect 18656 31368 18889 31396
rect 18656 31356 18662 31368
rect 18877 31365 18889 31368
rect 18923 31365 18935 31399
rect 20070 31396 20076 31408
rect 20031 31368 20076 31396
rect 18877 31359 18935 31365
rect 20070 31356 20076 31368
rect 20128 31356 20134 31408
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18233 31331 18291 31337
rect 18233 31328 18245 31331
rect 18012 31300 18245 31328
rect 18012 31288 18018 31300
rect 18233 31297 18245 31300
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 15396 31260 15424 31288
rect 18782 31260 18788 31272
rect 14016 31232 15424 31260
rect 18743 31232 18788 31260
rect 18782 31220 18788 31232
rect 18840 31220 18846 31272
rect 18966 31220 18972 31272
rect 19024 31260 19030 31272
rect 19981 31263 20039 31269
rect 19024 31232 19932 31260
rect 19024 31220 19030 31232
rect 10428 31164 11284 31192
rect 12066 31152 12072 31204
rect 12124 31192 12130 31204
rect 13541 31195 13599 31201
rect 13541 31192 13553 31195
rect 12124 31164 13553 31192
rect 12124 31152 12130 31164
rect 13541 31161 13553 31164
rect 13587 31161 13599 31195
rect 13541 31155 13599 31161
rect 13630 31152 13636 31204
rect 13688 31192 13694 31204
rect 15473 31195 15531 31201
rect 15473 31192 15485 31195
rect 13688 31164 15485 31192
rect 13688 31152 13694 31164
rect 15473 31161 15485 31164
rect 15519 31161 15531 31195
rect 15473 31155 15531 31161
rect 19150 31152 19156 31204
rect 19208 31192 19214 31204
rect 19337 31195 19395 31201
rect 19337 31192 19349 31195
rect 19208 31164 19349 31192
rect 19208 31152 19214 31164
rect 19337 31161 19349 31164
rect 19383 31192 19395 31195
rect 19904 31192 19932 31232
rect 19981 31229 19993 31263
rect 20027 31260 20039 31263
rect 22066 31260 22094 31436
rect 31754 31424 31760 31436
rect 31812 31424 31818 31476
rect 25038 31328 25044 31340
rect 24999 31300 25044 31328
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 25222 31288 25228 31340
rect 25280 31328 25286 31340
rect 25685 31331 25743 31337
rect 25685 31328 25697 31331
rect 25280 31300 25697 31328
rect 25280 31288 25286 31300
rect 25685 31297 25697 31300
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31328 32367 31331
rect 36078 31328 36084 31340
rect 32355 31300 36084 31328
rect 32355 31297 32367 31300
rect 32309 31291 32367 31297
rect 36078 31288 36084 31300
rect 36136 31288 36142 31340
rect 20027 31232 22094 31260
rect 25501 31263 25559 31269
rect 20027 31229 20039 31232
rect 19981 31223 20039 31229
rect 25501 31229 25513 31263
rect 25547 31260 25559 31263
rect 28994 31260 29000 31272
rect 25547 31232 29000 31260
rect 25547 31229 25559 31232
rect 25501 31223 25559 31229
rect 28994 31220 29000 31232
rect 29052 31220 29058 31272
rect 20533 31195 20591 31201
rect 20533 31192 20545 31195
rect 19383 31164 19840 31192
rect 19904 31164 20545 31192
rect 19383 31161 19395 31164
rect 19337 31155 19395 31161
rect 12161 31127 12219 31133
rect 12161 31124 12173 31127
rect 8680 31096 12173 31124
rect 12161 31093 12173 31096
rect 12207 31093 12219 31127
rect 12894 31124 12900 31136
rect 12855 31096 12900 31124
rect 12161 31087 12219 31093
rect 12894 31084 12900 31096
rect 12952 31084 12958 31136
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 14829 31127 14887 31133
rect 14829 31124 14841 31127
rect 13872 31096 14841 31124
rect 13872 31084 13878 31096
rect 14829 31093 14841 31096
rect 14875 31093 14887 31127
rect 14829 31087 14887 31093
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 16117 31127 16175 31133
rect 16117 31124 16129 31127
rect 15344 31096 16129 31124
rect 15344 31084 15350 31096
rect 16117 31093 16129 31096
rect 16163 31093 16175 31127
rect 16117 31087 16175 31093
rect 18049 31127 18107 31133
rect 18049 31093 18061 31127
rect 18095 31124 18107 31127
rect 19610 31124 19616 31136
rect 18095 31096 19616 31124
rect 18095 31093 18107 31096
rect 18049 31087 18107 31093
rect 19610 31084 19616 31096
rect 19668 31084 19674 31136
rect 19812 31124 19840 31164
rect 20533 31161 20545 31164
rect 20579 31161 20591 31195
rect 20533 31155 20591 31161
rect 25314 31152 25320 31204
rect 25372 31192 25378 31204
rect 25869 31195 25927 31201
rect 25869 31192 25881 31195
rect 25372 31164 25881 31192
rect 25372 31152 25378 31164
rect 25869 31161 25881 31164
rect 25915 31161 25927 31195
rect 25869 31155 25927 31161
rect 20714 31124 20720 31136
rect 19812 31096 20720 31124
rect 20714 31084 20720 31096
rect 20772 31084 20778 31136
rect 24857 31127 24915 31133
rect 24857 31093 24869 31127
rect 24903 31124 24915 31127
rect 25590 31124 25596 31136
rect 24903 31096 25596 31124
rect 24903 31093 24915 31096
rect 24857 31087 24915 31093
rect 25590 31084 25596 31096
rect 25648 31084 25654 31136
rect 32398 31124 32404 31136
rect 32359 31096 32404 31124
rect 32398 31084 32404 31096
rect 32456 31084 32462 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 4890 30880 4896 30932
rect 4948 30920 4954 30932
rect 5350 30920 5356 30932
rect 4948 30892 5356 30920
rect 4948 30880 4954 30892
rect 5350 30880 5356 30892
rect 5408 30880 5414 30932
rect 5902 30880 5908 30932
rect 5960 30880 5966 30932
rect 6270 30880 6276 30932
rect 6328 30920 6334 30932
rect 6822 30920 6828 30932
rect 6328 30892 6828 30920
rect 6328 30880 6334 30892
rect 6822 30880 6828 30892
rect 6880 30920 6886 30932
rect 9582 30920 9588 30932
rect 6880 30892 9588 30920
rect 6880 30880 6886 30892
rect 9582 30880 9588 30892
rect 9640 30880 9646 30932
rect 10597 30923 10655 30929
rect 10597 30889 10609 30923
rect 10643 30920 10655 30923
rect 11974 30920 11980 30932
rect 10643 30892 11744 30920
rect 11935 30892 11980 30920
rect 10643 30889 10655 30892
rect 10597 30883 10655 30889
rect 5920 30852 5948 30880
rect 7374 30852 7380 30864
rect 5920 30824 7380 30852
rect 7374 30812 7380 30824
rect 7432 30812 7438 30864
rect 7837 30855 7895 30861
rect 7837 30821 7849 30855
rect 7883 30852 7895 30855
rect 11606 30852 11612 30864
rect 7883 30824 11612 30852
rect 7883 30821 7895 30824
rect 7837 30815 7895 30821
rect 11606 30812 11612 30824
rect 11664 30812 11670 30864
rect 11716 30852 11744 30892
rect 11974 30880 11980 30892
rect 12032 30880 12038 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 13265 30923 13323 30929
rect 13265 30920 13277 30923
rect 12492 30892 13277 30920
rect 12492 30880 12498 30892
rect 13265 30889 13277 30892
rect 13311 30889 13323 30923
rect 13265 30883 13323 30889
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 14369 30923 14427 30929
rect 14369 30920 14381 30923
rect 13780 30892 14381 30920
rect 13780 30880 13786 30892
rect 14369 30889 14381 30892
rect 14415 30889 14427 30923
rect 14369 30883 14427 30889
rect 18782 30880 18788 30932
rect 18840 30920 18846 30932
rect 21174 30920 21180 30932
rect 18840 30892 21180 30920
rect 18840 30880 18846 30892
rect 21174 30880 21180 30892
rect 21232 30920 21238 30932
rect 24673 30923 24731 30929
rect 24673 30920 24685 30923
rect 21232 30892 24685 30920
rect 21232 30880 21238 30892
rect 24673 30889 24685 30892
rect 24719 30889 24731 30923
rect 24673 30883 24731 30889
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 26602 30920 26608 30932
rect 24912 30892 26608 30920
rect 24912 30880 24918 30892
rect 26602 30880 26608 30892
rect 26660 30880 26666 30932
rect 11716 30824 12020 30852
rect 11992 30796 12020 30824
rect 12986 30812 12992 30864
rect 13044 30852 13050 30864
rect 15194 30852 15200 30864
rect 13044 30824 15200 30852
rect 13044 30812 13050 30824
rect 15194 30812 15200 30824
rect 15252 30812 15258 30864
rect 18230 30812 18236 30864
rect 18288 30852 18294 30864
rect 27341 30855 27399 30861
rect 27341 30852 27353 30855
rect 18288 30824 27353 30852
rect 18288 30812 18294 30824
rect 27341 30821 27353 30824
rect 27387 30821 27399 30855
rect 27341 30815 27399 30821
rect 2038 30744 2044 30796
rect 2096 30784 2102 30796
rect 2133 30787 2191 30793
rect 2133 30784 2145 30787
rect 2096 30756 2145 30784
rect 2096 30744 2102 30756
rect 2133 30753 2145 30756
rect 2179 30784 2191 30787
rect 2314 30784 2320 30796
rect 2179 30756 2320 30784
rect 2179 30753 2191 30756
rect 2133 30747 2191 30753
rect 2314 30744 2320 30756
rect 2372 30744 2378 30796
rect 4890 30744 4896 30796
rect 4948 30784 4954 30796
rect 9401 30787 9459 30793
rect 4948 30756 7788 30784
rect 4948 30744 4954 30756
rect 1854 30716 1860 30728
rect 1815 30688 1860 30716
rect 1854 30676 1860 30688
rect 1912 30676 1918 30728
rect 2222 30676 2228 30728
rect 2280 30716 2286 30728
rect 2777 30719 2835 30725
rect 2777 30716 2789 30719
rect 2280 30688 2789 30716
rect 2280 30676 2286 30688
rect 2777 30685 2789 30688
rect 2823 30716 2835 30719
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 2823 30688 3985 30716
rect 2823 30685 2835 30688
rect 2777 30679 2835 30685
rect 3973 30685 3985 30688
rect 4019 30716 4031 30719
rect 4617 30719 4675 30725
rect 4617 30716 4629 30719
rect 4019 30688 4629 30716
rect 4019 30685 4031 30688
rect 3973 30679 4031 30685
rect 4617 30685 4629 30688
rect 4663 30716 4675 30719
rect 5626 30716 5632 30728
rect 4663 30688 5632 30716
rect 4663 30685 4675 30688
rect 4617 30679 4675 30685
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 5994 30716 6000 30728
rect 5955 30688 6000 30716
rect 5994 30676 6000 30688
rect 6052 30676 6058 30728
rect 6638 30716 6644 30728
rect 6599 30688 6644 30716
rect 6638 30676 6644 30688
rect 6696 30676 6702 30728
rect 6822 30676 6828 30728
rect 6880 30716 6886 30728
rect 7760 30725 7788 30756
rect 9401 30753 9413 30787
rect 9447 30784 9459 30787
rect 10137 30787 10195 30793
rect 9447 30756 10088 30784
rect 9447 30753 9459 30756
rect 9401 30747 9459 30753
rect 7101 30719 7159 30725
rect 7101 30716 7113 30719
rect 6880 30688 7113 30716
rect 6880 30676 6886 30688
rect 7101 30685 7113 30688
rect 7147 30685 7159 30719
rect 7101 30679 7159 30685
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30716 7803 30719
rect 8573 30719 8631 30725
rect 7791 30688 8524 30716
rect 7791 30685 7803 30688
rect 7745 30679 7803 30685
rect 6086 30608 6092 30660
rect 6144 30648 6150 30660
rect 6144 30620 8432 30648
rect 6144 30608 6150 30620
rect 2869 30583 2927 30589
rect 2869 30549 2881 30583
rect 2915 30580 2927 30583
rect 2958 30580 2964 30592
rect 2915 30552 2964 30580
rect 2915 30549 2927 30552
rect 2869 30543 2927 30549
rect 2958 30540 2964 30552
rect 3016 30540 3022 30592
rect 3878 30540 3884 30592
rect 3936 30580 3942 30592
rect 4065 30583 4123 30589
rect 4065 30580 4077 30583
rect 3936 30552 4077 30580
rect 3936 30540 3942 30552
rect 4065 30549 4077 30552
rect 4111 30549 4123 30583
rect 4065 30543 4123 30549
rect 4614 30540 4620 30592
rect 4672 30580 4678 30592
rect 4709 30583 4767 30589
rect 4709 30580 4721 30583
rect 4672 30552 4721 30580
rect 4672 30540 4678 30552
rect 4709 30549 4721 30552
rect 4755 30549 4767 30583
rect 4709 30543 4767 30549
rect 4982 30540 4988 30592
rect 5040 30580 5046 30592
rect 5813 30583 5871 30589
rect 5813 30580 5825 30583
rect 5040 30552 5825 30580
rect 5040 30540 5046 30552
rect 5813 30549 5825 30552
rect 5859 30549 5871 30583
rect 5813 30543 5871 30549
rect 6457 30583 6515 30589
rect 6457 30549 6469 30583
rect 6503 30580 6515 30583
rect 7098 30580 7104 30592
rect 6503 30552 7104 30580
rect 6503 30549 6515 30552
rect 6457 30543 6515 30549
rect 7098 30540 7104 30552
rect 7156 30540 7162 30592
rect 7190 30540 7196 30592
rect 7248 30580 7254 30592
rect 8404 30589 8432 30620
rect 8389 30583 8447 30589
rect 7248 30552 7293 30580
rect 7248 30540 7254 30552
rect 8389 30549 8401 30583
rect 8435 30549 8447 30583
rect 8496 30580 8524 30688
rect 8573 30685 8585 30719
rect 8619 30716 8631 30719
rect 9306 30716 9312 30728
rect 8619 30688 9312 30716
rect 8619 30685 8631 30688
rect 8573 30679 8631 30685
rect 9306 30676 9312 30688
rect 9364 30676 9370 30728
rect 9953 30719 10011 30725
rect 9953 30685 9965 30719
rect 9999 30685 10011 30719
rect 10060 30716 10088 30756
rect 10137 30753 10149 30787
rect 10183 30784 10195 30787
rect 10226 30784 10232 30796
rect 10183 30756 10232 30784
rect 10183 30753 10195 30756
rect 10137 30747 10195 30753
rect 10226 30744 10232 30756
rect 10284 30744 10290 30796
rect 11974 30744 11980 30796
rect 12032 30744 12038 30796
rect 19426 30784 19432 30796
rect 12452 30756 19432 30784
rect 11054 30716 11060 30728
rect 10060 30688 11060 30716
rect 9953 30679 10011 30685
rect 9968 30648 9996 30679
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 11241 30719 11299 30725
rect 11241 30716 11253 30719
rect 11204 30688 11253 30716
rect 11204 30676 11210 30688
rect 11241 30685 11253 30688
rect 11287 30685 11299 30719
rect 11882 30716 11888 30728
rect 11843 30688 11888 30716
rect 11241 30679 11299 30685
rect 11882 30676 11888 30688
rect 11940 30676 11946 30728
rect 12452 30716 12480 30756
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 26142 30784 26148 30796
rect 26103 30756 26148 30784
rect 26142 30744 26148 30756
rect 26200 30744 26206 30796
rect 12529 30719 12587 30725
rect 12529 30716 12541 30719
rect 12452 30688 12541 30716
rect 12529 30685 12541 30688
rect 12575 30685 12587 30719
rect 12529 30679 12587 30685
rect 12621 30719 12679 30725
rect 12621 30685 12633 30719
rect 12667 30718 12679 30719
rect 12667 30716 12756 30718
rect 12802 30716 12808 30728
rect 12667 30690 12808 30716
rect 12667 30685 12679 30690
rect 12728 30688 12808 30690
rect 12621 30679 12679 30685
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 13078 30676 13084 30728
rect 13136 30716 13142 30728
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 13136 30688 13185 30716
rect 13136 30676 13142 30688
rect 13173 30685 13185 30688
rect 13219 30685 13231 30719
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 13173 30679 13231 30685
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 14734 30676 14740 30728
rect 14792 30716 14798 30728
rect 14921 30719 14979 30725
rect 14921 30716 14933 30719
rect 14792 30688 14933 30716
rect 14792 30676 14798 30688
rect 14921 30685 14933 30688
rect 14967 30716 14979 30719
rect 15749 30719 15807 30725
rect 15749 30716 15761 30719
rect 14967 30688 15761 30716
rect 14967 30685 14979 30688
rect 14921 30679 14979 30685
rect 15749 30685 15761 30688
rect 15795 30685 15807 30719
rect 15749 30679 15807 30685
rect 16485 30719 16543 30725
rect 16485 30685 16497 30719
rect 16531 30685 16543 30719
rect 19610 30716 19616 30728
rect 19571 30688 19616 30716
rect 16485 30679 16543 30685
rect 10870 30648 10876 30660
rect 9968 30620 10876 30648
rect 10870 30608 10876 30620
rect 10928 30608 10934 30660
rect 16500 30648 16528 30679
rect 19610 30676 19616 30688
rect 19668 30676 19674 30728
rect 24581 30719 24639 30725
rect 24581 30685 24593 30719
rect 24627 30716 24639 30719
rect 24670 30716 24676 30728
rect 24627 30688 24676 30716
rect 24627 30685 24639 30688
rect 24581 30679 24639 30685
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 26602 30716 26608 30728
rect 26563 30688 26608 30716
rect 26602 30676 26608 30688
rect 26660 30676 26666 30728
rect 27249 30719 27307 30725
rect 27249 30685 27261 30719
rect 27295 30716 27307 30719
rect 30650 30716 30656 30728
rect 27295 30688 30656 30716
rect 27295 30685 27307 30688
rect 27249 30679 27307 30685
rect 30650 30676 30656 30688
rect 30708 30676 30714 30728
rect 18230 30648 18236 30660
rect 15580 30620 16528 30648
rect 18191 30620 18236 30648
rect 10410 30580 10416 30592
rect 8496 30552 10416 30580
rect 8389 30543 8447 30549
rect 10410 30540 10416 30552
rect 10468 30540 10474 30592
rect 10686 30540 10692 30592
rect 10744 30580 10750 30592
rect 11057 30583 11115 30589
rect 11057 30580 11069 30583
rect 10744 30552 11069 30580
rect 10744 30540 10750 30552
rect 11057 30549 11069 30552
rect 11103 30549 11115 30583
rect 11057 30543 11115 30549
rect 11514 30540 11520 30592
rect 11572 30580 11578 30592
rect 12066 30580 12072 30592
rect 11572 30552 12072 30580
rect 11572 30540 11578 30552
rect 12066 30540 12072 30552
rect 12124 30540 12130 30592
rect 15013 30583 15071 30589
rect 15013 30549 15025 30583
rect 15059 30580 15071 30583
rect 15378 30580 15384 30592
rect 15059 30552 15384 30580
rect 15059 30549 15071 30552
rect 15013 30543 15071 30549
rect 15378 30540 15384 30552
rect 15436 30540 15442 30592
rect 15580 30589 15608 30620
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 18322 30608 18328 30660
rect 18380 30648 18386 30660
rect 18877 30651 18935 30657
rect 18380 30620 18425 30648
rect 18380 30608 18386 30620
rect 18877 30617 18889 30651
rect 18923 30648 18935 30651
rect 18966 30648 18972 30660
rect 18923 30620 18972 30648
rect 18923 30617 18935 30620
rect 18877 30611 18935 30617
rect 18966 30608 18972 30620
rect 19024 30608 19030 30660
rect 25314 30608 25320 30660
rect 25372 30648 25378 30660
rect 25501 30651 25559 30657
rect 25501 30648 25513 30651
rect 25372 30620 25513 30648
rect 25372 30608 25378 30620
rect 25501 30617 25513 30620
rect 25547 30617 25559 30651
rect 25501 30611 25559 30617
rect 25593 30651 25651 30657
rect 25593 30617 25605 30651
rect 25639 30617 25651 30651
rect 25593 30611 25651 30617
rect 15565 30583 15623 30589
rect 15565 30549 15577 30583
rect 15611 30549 15623 30583
rect 16298 30580 16304 30592
rect 16259 30552 16304 30580
rect 15565 30543 15623 30549
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 19426 30580 19432 30592
rect 19387 30552 19432 30580
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 25608 30580 25636 30611
rect 26697 30583 26755 30589
rect 26697 30580 26709 30583
rect 25608 30552 26709 30580
rect 26697 30549 26709 30552
rect 26743 30549 26755 30583
rect 26697 30543 26755 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 5813 30379 5871 30385
rect 5813 30345 5825 30379
rect 5859 30376 5871 30379
rect 6638 30376 6644 30388
rect 5859 30348 6644 30376
rect 5859 30345 5871 30348
rect 5813 30339 5871 30345
rect 6638 30336 6644 30348
rect 6696 30336 6702 30388
rect 7300 30348 8248 30376
rect 7300 30308 7328 30348
rect 3358 30280 7328 30308
rect 8220 30308 8248 30348
rect 9508 30348 10456 30376
rect 9508 30308 9536 30348
rect 8220 30280 9536 30308
rect 10428 30308 10456 30348
rect 12342 30336 12348 30388
rect 12400 30376 12406 30388
rect 12400 30348 14412 30376
rect 12400 30336 12406 30348
rect 13446 30308 13452 30320
rect 10428 30280 13308 30308
rect 13407 30280 13452 30308
rect 1578 30200 1584 30252
rect 1636 30240 1642 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1636 30212 1869 30240
rect 1636 30200 1642 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 1857 30203 1915 30209
rect 4525 30244 4583 30249
rect 4525 30243 4660 30244
rect 4525 30209 4537 30243
rect 4571 30216 4660 30243
rect 4571 30209 4583 30216
rect 4525 30203 4583 30209
rect 2133 30175 2191 30181
rect 2133 30141 2145 30175
rect 2179 30172 2191 30175
rect 3418 30172 3424 30184
rect 2179 30144 3424 30172
rect 2179 30141 2191 30144
rect 2133 30135 2191 30141
rect 3418 30132 3424 30144
rect 3476 30132 3482 30184
rect 3881 30175 3939 30181
rect 3881 30141 3893 30175
rect 3927 30172 3939 30175
rect 3970 30172 3976 30184
rect 3927 30144 3976 30172
rect 3927 30141 3939 30144
rect 3881 30135 3939 30141
rect 3970 30132 3976 30144
rect 4028 30132 4034 30184
rect 4632 30172 4660 30216
rect 4985 30243 5043 30249
rect 4985 30209 4997 30243
rect 5031 30240 5043 30243
rect 5626 30240 5632 30252
rect 5031 30212 5632 30240
rect 5031 30209 5043 30212
rect 4985 30203 5043 30209
rect 5626 30200 5632 30212
rect 5684 30200 5690 30252
rect 5997 30243 6055 30249
rect 5997 30209 6009 30243
rect 6043 30240 6055 30243
rect 6270 30240 6276 30252
rect 6043 30212 6276 30240
rect 6043 30209 6055 30212
rect 5997 30203 6055 30209
rect 6270 30200 6276 30212
rect 6328 30200 6334 30252
rect 5166 30172 5172 30184
rect 4632 30144 5172 30172
rect 5166 30132 5172 30144
rect 5224 30132 5230 30184
rect 5902 30132 5908 30184
rect 5960 30172 5966 30184
rect 6546 30172 6552 30184
rect 5960 30144 6552 30172
rect 5960 30132 5966 30144
rect 6546 30132 6552 30144
rect 6604 30172 6610 30184
rect 6641 30175 6699 30181
rect 6641 30172 6653 30175
rect 6604 30144 6653 30172
rect 6604 30132 6610 30144
rect 6641 30141 6653 30144
rect 6687 30141 6699 30175
rect 6641 30135 6699 30141
rect 6917 30175 6975 30181
rect 6917 30141 6929 30175
rect 6963 30172 6975 30175
rect 6963 30144 7972 30172
rect 6963 30141 6975 30144
rect 6917 30135 6975 30141
rect 1946 29996 1952 30048
rect 2004 30036 2010 30048
rect 4341 30039 4399 30045
rect 4341 30036 4353 30039
rect 2004 30008 4353 30036
rect 2004 29996 2010 30008
rect 4341 30005 4353 30008
rect 4387 30005 4399 30039
rect 5074 30036 5080 30048
rect 5035 30008 5080 30036
rect 4341 29999 4399 30005
rect 5074 29996 5080 30008
rect 5132 29996 5138 30048
rect 7944 30036 7972 30144
rect 8036 30104 8064 30226
rect 10226 30200 10232 30252
rect 10284 30200 10290 30252
rect 10778 30240 10784 30252
rect 10428 30212 10784 30240
rect 8754 30132 8760 30184
rect 8812 30172 8818 30184
rect 8849 30175 8907 30181
rect 8849 30172 8861 30175
rect 8812 30144 8861 30172
rect 8812 30132 8818 30144
rect 8849 30141 8861 30144
rect 8895 30141 8907 30175
rect 8849 30135 8907 30141
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 10428 30172 10456 30212
rect 10778 30200 10784 30212
rect 10836 30200 10842 30252
rect 10962 30200 10968 30252
rect 11020 30240 11026 30252
rect 11020 30212 12296 30240
rect 11020 30200 11026 30212
rect 9171 30144 10456 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 10502 30132 10508 30184
rect 10560 30172 10566 30184
rect 11701 30175 11759 30181
rect 11701 30172 11713 30175
rect 10560 30144 11713 30172
rect 10560 30132 10566 30144
rect 11701 30141 11713 30144
rect 11747 30141 11759 30175
rect 12268 30172 12296 30212
rect 12526 30200 12532 30252
rect 12584 30240 12590 30252
rect 12989 30243 13047 30249
rect 12989 30240 13001 30243
rect 12584 30212 13001 30240
rect 12584 30200 12590 30212
rect 12989 30209 13001 30212
rect 13035 30209 13047 30243
rect 13280 30240 13308 30280
rect 13446 30268 13452 30280
rect 13504 30268 13510 30320
rect 14384 30317 14412 30348
rect 18322 30336 18328 30388
rect 18380 30376 18386 30388
rect 18693 30379 18751 30385
rect 18693 30376 18705 30379
rect 18380 30348 18705 30376
rect 18380 30336 18386 30348
rect 18693 30345 18705 30348
rect 18739 30345 18751 30379
rect 18693 30339 18751 30345
rect 14369 30311 14427 30317
rect 14369 30277 14381 30311
rect 14415 30277 14427 30311
rect 17678 30308 17684 30320
rect 17639 30280 17684 30308
rect 14369 30271 14427 30277
rect 13814 30240 13820 30252
rect 13280 30212 13820 30240
rect 12989 30203 13047 30209
rect 13814 30200 13820 30212
rect 13872 30200 13878 30252
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30240 13967 30243
rect 13998 30240 14004 30252
rect 13955 30212 14004 30240
rect 13955 30209 13967 30212
rect 13909 30203 13967 30209
rect 13998 30200 14004 30212
rect 14056 30200 14062 30252
rect 14384 30240 14412 30271
rect 17678 30268 17684 30280
rect 17736 30268 17742 30320
rect 19426 30268 19432 30320
rect 19484 30308 19490 30320
rect 19797 30311 19855 30317
rect 19797 30308 19809 30311
rect 19484 30280 19809 30308
rect 19484 30268 19490 30280
rect 19797 30277 19809 30280
rect 19843 30277 19855 30311
rect 25498 30308 25504 30320
rect 25459 30280 25504 30308
rect 19797 30271 19855 30277
rect 25498 30268 25504 30280
rect 25556 30268 25562 30320
rect 25590 30268 25596 30320
rect 25648 30308 25654 30320
rect 26142 30308 26148 30320
rect 25648 30280 25693 30308
rect 26103 30280 26148 30308
rect 25648 30268 25654 30280
rect 26142 30268 26148 30280
rect 26200 30268 26206 30320
rect 34606 30308 34612 30320
rect 31726 30280 34612 30308
rect 14921 30243 14979 30249
rect 14921 30240 14933 30243
rect 14384 30212 14933 30240
rect 14921 30209 14933 30212
rect 14967 30209 14979 30243
rect 14921 30203 14979 30209
rect 15378 30200 15384 30252
rect 15436 30240 15442 30252
rect 15657 30243 15715 30249
rect 15657 30240 15669 30243
rect 15436 30212 15669 30240
rect 15436 30200 15442 30212
rect 15657 30209 15669 30212
rect 15703 30209 15715 30243
rect 15657 30203 15715 30209
rect 17494 30200 17500 30252
rect 17552 30240 17558 30252
rect 17589 30243 17647 30249
rect 17589 30240 17601 30243
rect 17552 30212 17601 30240
rect 17552 30200 17558 30212
rect 17589 30209 17601 30212
rect 17635 30209 17647 30243
rect 17589 30203 17647 30209
rect 17862 30200 17868 30252
rect 17920 30240 17926 30252
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 17920 30212 18613 30240
rect 17920 30200 17926 30212
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 24854 30240 24860 30252
rect 24815 30212 24860 30240
rect 18601 30203 18659 30209
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 28077 30243 28135 30249
rect 28077 30209 28089 30243
rect 28123 30240 28135 30243
rect 31726 30240 31754 30280
rect 34606 30268 34612 30280
rect 34664 30268 34670 30320
rect 34422 30240 34428 30252
rect 28123 30212 31754 30240
rect 34383 30212 34428 30240
rect 28123 30209 28135 30212
rect 28077 30203 28135 30209
rect 34422 30200 34428 30212
rect 34480 30200 34486 30252
rect 38286 30240 38292 30252
rect 38247 30212 38292 30240
rect 38286 30200 38292 30212
rect 38344 30200 38350 30252
rect 15473 30175 15531 30181
rect 12268 30144 14044 30172
rect 11701 30135 11759 30141
rect 8036 30076 8984 30104
rect 8294 30036 8300 30048
rect 7944 30008 8300 30036
rect 8294 29996 8300 30008
rect 8352 29996 8358 30048
rect 8389 30039 8447 30045
rect 8389 30005 8401 30039
rect 8435 30036 8447 30039
rect 8662 30036 8668 30048
rect 8435 30008 8668 30036
rect 8435 30005 8447 30008
rect 8389 29999 8447 30005
rect 8662 29996 8668 30008
rect 8720 29996 8726 30048
rect 8956 30036 8984 30076
rect 10410 30064 10416 30116
rect 10468 30104 10474 30116
rect 12434 30104 12440 30116
rect 10468 30076 12440 30104
rect 10468 30064 10474 30076
rect 12434 30064 12440 30076
rect 12492 30064 12498 30116
rect 14016 30113 14044 30144
rect 15473 30141 15485 30175
rect 15519 30172 15531 30175
rect 17678 30172 17684 30184
rect 15519 30144 17684 30172
rect 15519 30141 15531 30144
rect 15473 30135 15531 30141
rect 17678 30132 17684 30144
rect 17736 30132 17742 30184
rect 19426 30132 19432 30184
rect 19484 30172 19490 30184
rect 19705 30175 19763 30181
rect 19705 30172 19717 30175
rect 19484 30144 19717 30172
rect 19484 30132 19490 30144
rect 19705 30141 19717 30144
rect 19751 30172 19763 30175
rect 28169 30175 28227 30181
rect 28169 30172 28181 30175
rect 19751 30144 28181 30172
rect 19751 30141 19763 30144
rect 19705 30135 19763 30141
rect 28169 30141 28181 30144
rect 28215 30141 28227 30175
rect 28169 30135 28227 30141
rect 14001 30107 14059 30113
rect 14001 30073 14013 30107
rect 14047 30073 14059 30107
rect 15838 30104 15844 30116
rect 15799 30076 15844 30104
rect 14001 30067 14059 30073
rect 15838 30064 15844 30076
rect 15896 30064 15902 30116
rect 20257 30107 20315 30113
rect 20257 30073 20269 30107
rect 20303 30104 20315 30107
rect 20438 30104 20444 30116
rect 20303 30076 20444 30104
rect 20303 30073 20315 30076
rect 20257 30067 20315 30073
rect 20438 30064 20444 30076
rect 20496 30064 20502 30116
rect 24673 30107 24731 30113
rect 24673 30073 24685 30107
rect 24719 30104 24731 30107
rect 25038 30104 25044 30116
rect 24719 30076 25044 30104
rect 24719 30073 24731 30076
rect 24673 30067 24731 30073
rect 25038 30064 25044 30076
rect 25096 30064 25102 30116
rect 34238 30104 34244 30116
rect 34199 30076 34244 30104
rect 34238 30064 34244 30076
rect 34296 30064 34302 30116
rect 10134 30036 10140 30048
rect 8956 30008 10140 30036
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 10318 29996 10324 30048
rect 10376 30036 10382 30048
rect 10597 30039 10655 30045
rect 10597 30036 10609 30039
rect 10376 30008 10609 30036
rect 10376 29996 10382 30008
rect 10597 30005 10609 30008
rect 10643 30036 10655 30039
rect 12710 30036 12716 30048
rect 10643 30008 12716 30036
rect 10643 30005 10655 30008
rect 10597 29999 10655 30005
rect 12710 29996 12716 30008
rect 12768 29996 12774 30048
rect 12805 30039 12863 30045
rect 12805 30005 12817 30039
rect 12851 30036 12863 30039
rect 13722 30036 13728 30048
rect 12851 30008 13728 30036
rect 12851 30005 12863 30008
rect 12805 29999 12863 30005
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 13814 29996 13820 30048
rect 13872 30036 13878 30048
rect 14737 30039 14795 30045
rect 14737 30036 14749 30039
rect 13872 30008 14749 30036
rect 13872 29996 13878 30008
rect 14737 30005 14749 30008
rect 14783 30005 14795 30039
rect 14737 29999 14795 30005
rect 36998 29996 37004 30048
rect 37056 30036 37062 30048
rect 38105 30039 38163 30045
rect 38105 30036 38117 30039
rect 37056 30008 38117 30036
rect 37056 29996 37062 30008
rect 38105 30005 38117 30008
rect 38151 30005 38163 30039
rect 38105 29999 38163 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 5442 29832 5448 29844
rect 4172 29804 5448 29832
rect 2133 29699 2191 29705
rect 2133 29665 2145 29699
rect 2179 29696 2191 29699
rect 2222 29696 2228 29708
rect 2179 29668 2228 29696
rect 2179 29665 2191 29668
rect 2133 29659 2191 29665
rect 2222 29656 2228 29668
rect 2280 29656 2286 29708
rect 3053 29699 3111 29705
rect 3053 29665 3065 29699
rect 3099 29696 3111 29699
rect 3694 29696 3700 29708
rect 3099 29668 3700 29696
rect 3099 29665 3111 29668
rect 3053 29659 3111 29665
rect 3694 29656 3700 29668
rect 3752 29696 3758 29708
rect 4062 29696 4068 29708
rect 3752 29668 4068 29696
rect 3752 29656 3758 29668
rect 4062 29656 4068 29668
rect 4120 29656 4126 29708
rect 1854 29628 1860 29640
rect 1815 29600 1860 29628
rect 1854 29588 1860 29600
rect 1912 29628 1918 29640
rect 4172 29637 4200 29804
rect 5442 29792 5448 29804
rect 5500 29792 5506 29844
rect 7285 29835 7343 29841
rect 7285 29801 7297 29835
rect 7331 29832 7343 29835
rect 9858 29832 9864 29844
rect 7331 29804 9864 29832
rect 7331 29801 7343 29804
rect 7285 29795 7343 29801
rect 9858 29792 9864 29804
rect 9916 29792 9922 29844
rect 10134 29792 10140 29844
rect 10192 29832 10198 29844
rect 10870 29832 10876 29844
rect 10192 29804 10876 29832
rect 10192 29792 10198 29804
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 11146 29792 11152 29844
rect 11204 29832 11210 29844
rect 11330 29832 11336 29844
rect 11204 29804 11336 29832
rect 11204 29792 11210 29804
rect 11330 29792 11336 29804
rect 11388 29792 11394 29844
rect 12069 29835 12127 29841
rect 12069 29801 12081 29835
rect 12115 29832 12127 29835
rect 12158 29832 12164 29844
rect 12115 29804 12164 29832
rect 12115 29801 12127 29804
rect 12069 29795 12127 29801
rect 12158 29792 12164 29804
rect 12216 29792 12222 29844
rect 23566 29832 23572 29844
rect 12406 29804 23572 29832
rect 9122 29764 9128 29776
rect 6012 29736 9128 29764
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 5902 29696 5908 29708
rect 4663 29668 5908 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 5902 29656 5908 29668
rect 5960 29656 5966 29708
rect 2777 29631 2835 29637
rect 2777 29628 2789 29631
rect 1912 29600 2789 29628
rect 1912 29588 1918 29600
rect 2777 29597 2789 29600
rect 2823 29597 2835 29631
rect 2777 29591 2835 29597
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29597 4215 29631
rect 6012 29614 6040 29736
rect 9122 29724 9128 29736
rect 9180 29724 9186 29776
rect 12406 29764 12434 29804
rect 23566 29792 23572 29804
rect 23624 29792 23630 29844
rect 12986 29764 12992 29776
rect 10428 29736 12434 29764
rect 12544 29736 12992 29764
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 8113 29699 8171 29705
rect 8113 29696 8125 29699
rect 7156 29668 8125 29696
rect 7156 29656 7162 29668
rect 8113 29665 8125 29668
rect 8159 29665 8171 29699
rect 10428 29696 10456 29736
rect 12544 29696 12572 29736
rect 12986 29724 12992 29736
rect 13044 29724 13050 29776
rect 13078 29724 13084 29776
rect 13136 29764 13142 29776
rect 13262 29764 13268 29776
rect 13136 29736 13268 29764
rect 13136 29724 13142 29736
rect 13262 29724 13268 29736
rect 13320 29724 13326 29776
rect 13541 29767 13599 29773
rect 13541 29733 13553 29767
rect 13587 29764 13599 29767
rect 15102 29764 15108 29776
rect 13587 29736 15108 29764
rect 13587 29733 13599 29736
rect 13541 29727 13599 29733
rect 15102 29724 15108 29736
rect 15160 29724 15166 29776
rect 15838 29724 15844 29776
rect 15896 29764 15902 29776
rect 17497 29767 17555 29773
rect 17497 29764 17509 29767
rect 15896 29736 17509 29764
rect 15896 29724 15902 29736
rect 17497 29733 17509 29736
rect 17543 29733 17555 29767
rect 17497 29727 17555 29733
rect 19610 29724 19616 29776
rect 19668 29724 19674 29776
rect 8113 29659 8171 29665
rect 8496 29668 10456 29696
rect 10520 29668 12572 29696
rect 7469 29631 7527 29637
rect 4157 29591 4215 29597
rect 7469 29597 7481 29631
rect 7515 29628 7527 29631
rect 7650 29628 7656 29640
rect 7515 29600 7656 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 7650 29588 7656 29600
rect 7708 29588 7714 29640
rect 7926 29628 7932 29640
rect 7887 29600 7932 29628
rect 7926 29588 7932 29600
rect 7984 29588 7990 29640
rect 4522 29520 4528 29572
rect 4580 29560 4586 29572
rect 4893 29563 4951 29569
rect 4893 29560 4905 29563
rect 4580 29532 4905 29560
rect 4580 29520 4586 29532
rect 4893 29529 4905 29532
rect 4939 29529 4951 29563
rect 4893 29523 4951 29529
rect 6641 29563 6699 29569
rect 6641 29529 6653 29563
rect 6687 29560 6699 29563
rect 7006 29560 7012 29572
rect 6687 29532 7012 29560
rect 6687 29529 6699 29532
rect 6641 29523 6699 29529
rect 7006 29520 7012 29532
rect 7064 29520 7070 29572
rect 7098 29520 7104 29572
rect 7156 29560 7162 29572
rect 8202 29560 8208 29572
rect 7156 29532 8208 29560
rect 7156 29520 7162 29532
rect 8202 29520 8208 29532
rect 8260 29520 8266 29572
rect 3326 29452 3332 29504
rect 3384 29492 3390 29504
rect 3973 29495 4031 29501
rect 3973 29492 3985 29495
rect 3384 29464 3985 29492
rect 3384 29452 3390 29464
rect 3973 29461 3985 29464
rect 4019 29461 4031 29495
rect 3973 29455 4031 29461
rect 4062 29452 4068 29504
rect 4120 29492 4126 29504
rect 8496 29492 8524 29668
rect 8754 29588 8760 29640
rect 8812 29628 8818 29640
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 8812 29600 9137 29628
rect 8812 29588 8818 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 10520 29614 10548 29668
rect 12710 29656 12716 29708
rect 12768 29696 12774 29708
rect 14182 29696 14188 29708
rect 12768 29668 14188 29696
rect 12768 29656 12774 29668
rect 14182 29656 14188 29668
rect 14240 29696 14246 29708
rect 14240 29668 14688 29696
rect 14240 29656 14246 29668
rect 9125 29591 9183 29597
rect 10870 29588 10876 29640
rect 10928 29628 10934 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 10928 29600 11437 29628
rect 10928 29588 10934 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11606 29628 11612 29640
rect 11567 29600 11612 29628
rect 11425 29591 11483 29597
rect 11606 29588 11612 29600
rect 11664 29588 11670 29640
rect 12621 29631 12679 29637
rect 12621 29597 12633 29631
rect 12667 29597 12679 29631
rect 13722 29628 13728 29640
rect 13683 29600 13728 29628
rect 12621 29591 12679 29597
rect 8662 29520 8668 29572
rect 8720 29560 8726 29572
rect 8938 29560 8944 29572
rect 8720 29532 8944 29560
rect 8720 29520 8726 29532
rect 8938 29520 8944 29532
rect 8996 29560 9002 29572
rect 9401 29563 9459 29569
rect 9401 29560 9413 29563
rect 8996 29532 9413 29560
rect 8996 29520 9002 29532
rect 9401 29529 9413 29532
rect 9447 29529 9459 29563
rect 11882 29560 11888 29572
rect 9401 29523 9459 29529
rect 10704 29532 11888 29560
rect 4120 29464 8524 29492
rect 4120 29452 4126 29464
rect 8570 29452 8576 29504
rect 8628 29492 8634 29504
rect 10704 29492 10732 29532
rect 11882 29520 11888 29532
rect 11940 29520 11946 29572
rect 11974 29520 11980 29572
rect 12032 29560 12038 29572
rect 12526 29560 12532 29572
rect 12032 29532 12532 29560
rect 12032 29520 12038 29532
rect 12526 29520 12532 29532
rect 12584 29560 12590 29572
rect 12636 29560 12664 29591
rect 13722 29588 13728 29600
rect 13780 29588 13786 29640
rect 14660 29637 14688 29668
rect 16298 29656 16304 29708
rect 16356 29696 16362 29708
rect 17313 29699 17371 29705
rect 17313 29696 17325 29699
rect 16356 29668 17325 29696
rect 16356 29656 16362 29668
rect 17313 29665 17325 29668
rect 17359 29665 17371 29699
rect 19518 29696 19524 29708
rect 17313 29659 17371 29665
rect 18708 29668 19524 29696
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29597 14703 29631
rect 14645 29591 14703 29597
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 15068 29600 15301 29628
rect 15068 29588 15074 29600
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 17129 29631 17187 29637
rect 17129 29597 17141 29631
rect 17175 29628 17187 29631
rect 18708 29628 18736 29668
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 19628 29647 19656 29724
rect 19613 29641 19671 29647
rect 18874 29628 18880 29640
rect 17175 29600 18736 29628
rect 18835 29600 18880 29628
rect 17175 29597 17187 29600
rect 17129 29591 17187 29597
rect 18874 29588 18880 29600
rect 18932 29588 18938 29640
rect 19150 29588 19156 29640
rect 19208 29628 19214 29640
rect 19208 29600 19564 29628
rect 19613 29607 19625 29641
rect 19659 29607 19671 29641
rect 19613 29601 19671 29607
rect 19208 29588 19214 29600
rect 12584 29532 12664 29560
rect 12584 29520 12590 29532
rect 10870 29492 10876 29504
rect 8628 29464 10732 29492
rect 10831 29464 10876 29492
rect 8628 29452 8634 29464
rect 10870 29452 10876 29464
rect 10928 29452 10934 29504
rect 12713 29495 12771 29501
rect 12713 29461 12725 29495
rect 12759 29492 12771 29495
rect 12986 29492 12992 29504
rect 12759 29464 12992 29492
rect 12759 29461 12771 29464
rect 12713 29455 12771 29461
rect 12986 29452 12992 29464
rect 13044 29452 13050 29504
rect 14458 29492 14464 29504
rect 14419 29464 14464 29492
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 15105 29495 15163 29501
rect 15105 29461 15117 29495
rect 15151 29492 15163 29495
rect 17034 29492 17040 29504
rect 15151 29464 17040 29492
rect 15151 29461 15163 29464
rect 15105 29455 15163 29461
rect 17034 29452 17040 29464
rect 17092 29452 17098 29504
rect 18693 29495 18751 29501
rect 18693 29461 18705 29495
rect 18739 29492 18751 29495
rect 19242 29492 19248 29504
rect 18739 29464 19248 29492
rect 18739 29461 18751 29464
rect 18693 29455 18751 29461
rect 19242 29452 19248 29464
rect 19300 29452 19306 29504
rect 19536 29492 19564 29600
rect 19794 29588 19800 29640
rect 19852 29628 19858 29640
rect 20257 29631 20315 29637
rect 20257 29628 20269 29631
rect 19852 29600 20269 29628
rect 19852 29588 19858 29600
rect 20257 29597 20269 29600
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 20346 29588 20352 29640
rect 20404 29628 20410 29640
rect 21545 29631 21603 29637
rect 21545 29628 21557 29631
rect 20404 29600 21557 29628
rect 20404 29588 20410 29600
rect 21545 29597 21557 29600
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 24765 29631 24823 29637
rect 24765 29597 24777 29631
rect 24811 29628 24823 29631
rect 25130 29628 25136 29640
rect 24811 29600 25136 29628
rect 24811 29597 24823 29600
rect 24765 29591 24823 29597
rect 25130 29588 25136 29600
rect 25188 29588 25194 29640
rect 19705 29563 19763 29569
rect 19705 29529 19717 29563
rect 19751 29560 19763 29563
rect 20806 29560 20812 29572
rect 19751 29532 20812 29560
rect 19751 29529 19763 29532
rect 19705 29523 19763 29529
rect 20806 29520 20812 29532
rect 20864 29520 20870 29572
rect 19794 29492 19800 29504
rect 19536 29464 19800 29492
rect 19794 29452 19800 29464
rect 19852 29452 19858 29504
rect 20162 29452 20168 29504
rect 20220 29492 20226 29504
rect 20349 29495 20407 29501
rect 20349 29492 20361 29495
rect 20220 29464 20361 29492
rect 20220 29452 20226 29464
rect 20349 29461 20361 29464
rect 20395 29461 20407 29495
rect 20349 29455 20407 29461
rect 20901 29495 20959 29501
rect 20901 29461 20913 29495
rect 20947 29492 20959 29495
rect 21266 29492 21272 29504
rect 20947 29464 21272 29492
rect 20947 29461 20959 29464
rect 20901 29455 20959 29461
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 21637 29495 21695 29501
rect 21637 29461 21649 29495
rect 21683 29492 21695 29495
rect 22186 29492 22192 29504
rect 21683 29464 22192 29492
rect 21683 29461 21695 29464
rect 21637 29455 21695 29461
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 24581 29495 24639 29501
rect 24581 29461 24593 29495
rect 24627 29492 24639 29495
rect 24946 29492 24952 29504
rect 24627 29464 24952 29492
rect 24627 29461 24639 29464
rect 24581 29455 24639 29461
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1854 29248 1860 29300
rect 1912 29288 1918 29300
rect 4062 29288 4068 29300
rect 1912 29260 4068 29288
rect 1912 29248 1918 29260
rect 4062 29248 4068 29260
rect 4120 29248 4126 29300
rect 4709 29291 4767 29297
rect 4709 29257 4721 29291
rect 4755 29288 4767 29291
rect 5997 29291 6055 29297
rect 4755 29260 5488 29288
rect 4755 29257 4767 29260
rect 4709 29251 4767 29257
rect 5258 29220 5264 29232
rect 3450 29192 5264 29220
rect 5258 29180 5264 29192
rect 5316 29180 5322 29232
rect 1578 29112 1584 29164
rect 1636 29152 1642 29164
rect 1949 29155 2007 29161
rect 1949 29152 1961 29155
rect 1636 29124 1961 29152
rect 1636 29112 1642 29124
rect 1949 29121 1961 29124
rect 1995 29121 2007 29155
rect 1949 29115 2007 29121
rect 3973 29155 4031 29161
rect 3973 29121 3985 29155
rect 4019 29152 4031 29155
rect 4062 29152 4068 29164
rect 4019 29124 4068 29152
rect 4019 29121 4031 29124
rect 3973 29115 4031 29121
rect 4062 29112 4068 29124
rect 4120 29112 4126 29164
rect 4890 29152 4896 29164
rect 4851 29124 4896 29152
rect 4890 29112 4896 29124
rect 4948 29112 4954 29164
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29053 5411 29087
rect 5460 29084 5488 29260
rect 5997 29257 6009 29291
rect 6043 29288 6055 29291
rect 8570 29288 8576 29300
rect 6043 29260 8576 29288
rect 6043 29257 6055 29260
rect 5997 29251 6055 29257
rect 8570 29248 8576 29260
rect 8628 29248 8634 29300
rect 8662 29248 8668 29300
rect 8720 29288 8726 29300
rect 10134 29288 10140 29300
rect 8720 29260 10140 29288
rect 8720 29248 8726 29260
rect 10134 29248 10140 29260
rect 10192 29248 10198 29300
rect 14274 29288 14280 29300
rect 10520 29260 14280 29288
rect 7190 29220 7196 29232
rect 5552 29192 7196 29220
rect 5552 29161 5580 29192
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 8754 29220 8760 29232
rect 8220 29192 8760 29220
rect 5537 29155 5595 29161
rect 5537 29121 5549 29155
rect 5583 29121 5595 29155
rect 7098 29152 7104 29164
rect 7059 29124 7104 29152
rect 5537 29115 5595 29121
rect 7098 29112 7104 29124
rect 7156 29112 7162 29164
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7374 29152 7380 29164
rect 7331 29124 7380 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 7926 29112 7932 29164
rect 7984 29152 7990 29164
rect 8220 29161 8248 29192
rect 8754 29180 8760 29192
rect 8812 29180 8818 29232
rect 10520 29220 10548 29260
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 19150 29288 19156 29300
rect 16408 29260 19156 29288
rect 9706 29192 10548 29220
rect 10594 29180 10600 29232
rect 10652 29220 10658 29232
rect 10652 29192 10697 29220
rect 10652 29180 10658 29192
rect 10778 29180 10784 29232
rect 10836 29220 10842 29232
rect 12250 29220 12256 29232
rect 10836 29192 12256 29220
rect 10836 29180 10842 29192
rect 12250 29180 12256 29192
rect 12308 29180 12314 29232
rect 14090 29220 14096 29232
rect 13202 29192 14096 29220
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 14458 29180 14464 29232
rect 14516 29220 14522 29232
rect 14516 29192 16068 29220
rect 14516 29180 14522 29192
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 7984 29124 8217 29152
rect 7984 29112 7990 29124
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 11698 29152 11704 29164
rect 11659 29124 11704 29152
rect 8205 29115 8263 29121
rect 11698 29112 11704 29124
rect 11756 29112 11762 29164
rect 13906 29152 13912 29164
rect 13188 29124 13912 29152
rect 9766 29084 9772 29096
rect 5460 29056 9772 29084
rect 5353 29047 5411 29053
rect 4890 28976 4896 29028
rect 4948 29016 4954 29028
rect 5368 29016 5396 29047
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 9950 29084 9956 29096
rect 9911 29056 9956 29084
rect 9950 29044 9956 29056
rect 10008 29084 10014 29096
rect 10318 29084 10324 29096
rect 10008 29056 10324 29084
rect 10008 29044 10014 29056
rect 10318 29044 10324 29056
rect 10376 29044 10382 29096
rect 10502 29084 10508 29096
rect 10463 29056 10508 29084
rect 10502 29044 10508 29056
rect 10560 29044 10566 29096
rect 11149 29087 11207 29093
rect 11149 29053 11161 29087
rect 11195 29084 11207 29087
rect 11330 29084 11336 29096
rect 11195 29056 11336 29084
rect 11195 29053 11207 29056
rect 11149 29047 11207 29053
rect 11330 29044 11336 29056
rect 11388 29044 11394 29096
rect 11977 29087 12035 29093
rect 11977 29053 11989 29087
rect 12023 29084 12035 29087
rect 12434 29084 12440 29096
rect 12023 29056 12440 29084
rect 12023 29053 12035 29056
rect 11977 29047 12035 29053
rect 12434 29044 12440 29056
rect 12492 29044 12498 29096
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 13188 29084 13216 29124
rect 13906 29112 13912 29124
rect 13964 29112 13970 29164
rect 14182 29152 14188 29164
rect 14143 29124 14188 29152
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 15010 29152 15016 29164
rect 14971 29124 15016 29152
rect 15010 29112 15016 29124
rect 15068 29112 15074 29164
rect 16040 29161 16068 29192
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29121 16083 29155
rect 16025 29115 16083 29121
rect 12584 29056 13216 29084
rect 13725 29087 13783 29093
rect 12584 29044 12590 29056
rect 13725 29053 13737 29087
rect 13771 29084 13783 29087
rect 16408 29084 16436 29260
rect 19150 29248 19156 29260
rect 19208 29248 19214 29300
rect 21085 29291 21143 29297
rect 21085 29257 21097 29291
rect 21131 29288 21143 29291
rect 21131 29260 22094 29288
rect 21131 29257 21143 29260
rect 21085 29251 21143 29257
rect 19334 29220 19340 29232
rect 17788 29192 19340 29220
rect 17034 29152 17040 29164
rect 16995 29124 17040 29152
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 17788 29161 17816 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 17773 29155 17831 29161
rect 17773 29121 17785 29155
rect 17819 29121 17831 29155
rect 17773 29115 17831 29121
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 18877 29155 18935 29161
rect 18877 29152 18889 29155
rect 18104 29124 18889 29152
rect 18104 29112 18110 29124
rect 18877 29121 18889 29124
rect 18923 29121 18935 29155
rect 20162 29152 20168 29164
rect 20123 29124 20168 29152
rect 18877 29115 18935 29121
rect 20162 29112 20168 29124
rect 20220 29112 20226 29164
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21358 29152 21364 29164
rect 21315 29124 21364 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21358 29112 21364 29124
rect 21416 29112 21422 29164
rect 22066 29152 22094 29260
rect 22922 29248 22928 29300
rect 22980 29288 22986 29300
rect 23477 29291 23535 29297
rect 23477 29288 23489 29291
rect 22980 29260 23489 29288
rect 22980 29248 22986 29260
rect 23477 29257 23489 29260
rect 23523 29257 23535 29291
rect 23477 29251 23535 29257
rect 23566 29220 23572 29232
rect 22756 29192 23572 29220
rect 22756 29161 22784 29192
rect 23566 29180 23572 29192
rect 23624 29180 23630 29232
rect 32398 29220 32404 29232
rect 31726 29192 32404 29220
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22066 29124 22201 29152
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22741 29155 22799 29161
rect 22741 29121 22753 29155
rect 22787 29121 22799 29155
rect 23382 29152 23388 29164
rect 23343 29124 23388 29152
rect 22741 29115 22799 29121
rect 23382 29112 23388 29124
rect 23440 29112 23446 29164
rect 25225 29155 25283 29161
rect 25225 29121 25237 29155
rect 25271 29152 25283 29155
rect 30374 29152 30380 29164
rect 25271 29124 30380 29152
rect 25271 29121 25283 29124
rect 25225 29115 25283 29121
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 13771 29056 16436 29084
rect 17957 29087 18015 29093
rect 13771 29053 13783 29056
rect 13725 29047 13783 29053
rect 17957 29053 17969 29087
rect 18003 29053 18015 29087
rect 18414 29084 18420 29096
rect 18375 29056 18420 29084
rect 17957 29047 18015 29053
rect 7469 29019 7527 29025
rect 7469 29016 7481 29019
rect 4948 28988 7481 29016
rect 4948 28976 4954 28988
rect 7469 28985 7481 28988
rect 7515 28985 7527 29019
rect 7469 28979 7527 28985
rect 9582 28976 9588 29028
rect 9640 29016 9646 29028
rect 10594 29016 10600 29028
rect 9640 28988 10600 29016
rect 9640 28976 9646 28988
rect 10594 28976 10600 28988
rect 10652 28976 10658 29028
rect 13170 28976 13176 29028
rect 13228 29016 13234 29028
rect 13740 29016 13768 29047
rect 14274 29016 14280 29028
rect 13228 28988 13768 29016
rect 14235 28988 14280 29016
rect 13228 28976 13234 28988
rect 14274 28976 14280 28988
rect 14332 28976 14338 29028
rect 14829 29019 14887 29025
rect 14829 28985 14841 29019
rect 14875 29016 14887 29019
rect 15194 29016 15200 29028
rect 14875 28988 15200 29016
rect 14875 28985 14887 28988
rect 14829 28979 14887 28985
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 15841 29019 15899 29025
rect 15841 28985 15853 29019
rect 15887 29016 15899 29019
rect 16758 29016 16764 29028
rect 15887 28988 16764 29016
rect 15887 28985 15899 28988
rect 15841 28979 15899 28985
rect 16758 28976 16764 28988
rect 16816 28976 16822 29028
rect 16853 29019 16911 29025
rect 16853 28985 16865 29019
rect 16899 29016 16911 29019
rect 17972 29016 18000 29047
rect 18414 29044 18420 29056
rect 18472 29044 18478 29096
rect 19981 29087 20039 29093
rect 19981 29053 19993 29087
rect 20027 29084 20039 29087
rect 31726 29084 31754 29192
rect 32398 29180 32404 29192
rect 32456 29180 32462 29232
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 20027 29056 31754 29084
rect 20027 29053 20039 29056
rect 19981 29047 20039 29053
rect 16899 28988 18000 29016
rect 16899 28985 16911 28988
rect 16853 28979 16911 28985
rect 18230 28976 18236 29028
rect 18288 29016 18294 29028
rect 18969 29019 19027 29025
rect 18969 29016 18981 29019
rect 18288 28988 18981 29016
rect 18288 28976 18294 28988
rect 18969 28985 18981 28988
rect 19015 28985 19027 29019
rect 18969 28979 19027 28985
rect 20625 29019 20683 29025
rect 20625 28985 20637 29019
rect 20671 29016 20683 29019
rect 20990 29016 20996 29028
rect 20671 28988 20996 29016
rect 20671 28985 20683 28988
rect 20625 28979 20683 28985
rect 20990 28976 20996 28988
rect 21048 28976 21054 29028
rect 22002 29016 22008 29028
rect 21963 28988 22008 29016
rect 22002 28976 22008 28988
rect 22060 28976 22066 29028
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 25317 29019 25375 29025
rect 25317 29016 25329 29019
rect 23348 28988 25329 29016
rect 23348 28976 23354 28988
rect 25317 28985 25329 28988
rect 25363 28985 25375 29019
rect 25317 28979 25375 28985
rect 35434 28976 35440 29028
rect 35492 29016 35498 29028
rect 38105 29019 38163 29025
rect 38105 29016 38117 29019
rect 35492 28988 38117 29016
rect 35492 28976 35498 28988
rect 38105 28985 38117 28988
rect 38151 28985 38163 29019
rect 38105 28979 38163 28985
rect 2212 28951 2270 28957
rect 2212 28917 2224 28951
rect 2258 28948 2270 28951
rect 2314 28948 2320 28960
rect 2258 28920 2320 28948
rect 2258 28917 2270 28920
rect 2212 28911 2270 28917
rect 2314 28908 2320 28920
rect 2372 28908 2378 28960
rect 5810 28908 5816 28960
rect 5868 28948 5874 28960
rect 8202 28948 8208 28960
rect 5868 28920 8208 28948
rect 5868 28908 5874 28920
rect 8202 28908 8208 28920
rect 8260 28908 8266 28960
rect 8468 28951 8526 28957
rect 8468 28917 8480 28951
rect 8514 28948 8526 28951
rect 9858 28948 9864 28960
rect 8514 28920 9864 28948
rect 8514 28917 8526 28920
rect 8468 28911 8526 28917
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 9950 28908 9956 28960
rect 10008 28948 10014 28960
rect 11238 28948 11244 28960
rect 10008 28920 11244 28948
rect 10008 28908 10014 28920
rect 11238 28908 11244 28920
rect 11296 28908 11302 28960
rect 11606 28908 11612 28960
rect 11664 28948 11670 28960
rect 11974 28948 11980 28960
rect 11664 28920 11980 28948
rect 11664 28908 11670 28920
rect 11974 28908 11980 28920
rect 12032 28908 12038 28960
rect 22830 28948 22836 28960
rect 22791 28920 22836 28948
rect 22830 28908 22836 28920
rect 22888 28908 22894 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 2590 28704 2596 28756
rect 2648 28744 2654 28756
rect 4522 28744 4528 28756
rect 2648 28716 4528 28744
rect 2648 28704 2654 28716
rect 4522 28704 4528 28716
rect 4580 28704 4586 28756
rect 7742 28744 7748 28756
rect 5736 28716 7748 28744
rect 5736 28676 5764 28716
rect 7742 28704 7748 28716
rect 7800 28704 7806 28756
rect 8389 28747 8447 28753
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 9582 28744 9588 28756
rect 8435 28716 9588 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 9582 28704 9588 28716
rect 9640 28704 9646 28756
rect 10686 28744 10692 28756
rect 9876 28716 10692 28744
rect 2976 28648 5764 28676
rect 1854 28608 1860 28620
rect 1815 28580 1860 28608
rect 1854 28568 1860 28580
rect 1912 28568 1918 28620
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 2976 28526 3004 28648
rect 7558 28636 7564 28688
rect 7616 28676 7622 28688
rect 7653 28679 7711 28685
rect 7653 28676 7665 28679
rect 7616 28648 7665 28676
rect 7616 28636 7622 28648
rect 7653 28645 7665 28648
rect 7699 28645 7711 28679
rect 7653 28639 7711 28645
rect 4982 28608 4988 28620
rect 4943 28580 4988 28608
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 5810 28568 5816 28620
rect 5868 28608 5874 28620
rect 6181 28611 6239 28617
rect 6181 28608 6193 28611
rect 5868 28580 6193 28608
rect 5868 28568 5874 28580
rect 6181 28577 6193 28580
rect 6227 28608 6239 28611
rect 9876 28608 9904 28716
rect 10686 28704 10692 28716
rect 10744 28704 10750 28756
rect 10778 28704 10784 28756
rect 10836 28744 10842 28756
rect 16669 28747 16727 28753
rect 10836 28716 16620 28744
rect 10836 28704 10842 28716
rect 11422 28636 11428 28688
rect 11480 28676 11486 28688
rect 14090 28676 14096 28688
rect 11480 28648 14096 28676
rect 11480 28636 11486 28648
rect 14090 28636 14096 28648
rect 14148 28676 14154 28688
rect 14642 28676 14648 28688
rect 14148 28648 14648 28676
rect 14148 28636 14154 28648
rect 14642 28636 14648 28648
rect 14700 28636 14706 28688
rect 16592 28676 16620 28716
rect 16669 28713 16681 28747
rect 16715 28744 16727 28747
rect 18874 28744 18880 28756
rect 16715 28716 18880 28744
rect 16715 28713 16727 28716
rect 16669 28707 16727 28713
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 24026 28744 24032 28756
rect 19536 28716 24032 28744
rect 17862 28676 17868 28688
rect 16592 28648 17868 28676
rect 17862 28636 17868 28648
rect 17920 28636 17926 28688
rect 17957 28679 18015 28685
rect 17957 28645 17969 28679
rect 18003 28645 18015 28679
rect 17957 28639 18015 28645
rect 10042 28608 10048 28620
rect 6227 28580 8156 28608
rect 6227 28577 6239 28580
rect 6181 28571 6239 28577
rect 4157 28543 4215 28549
rect 4157 28509 4169 28543
rect 4203 28540 4215 28543
rect 4430 28540 4436 28552
rect 4203 28512 4436 28540
rect 4203 28509 4215 28512
rect 4157 28503 4215 28509
rect 4430 28500 4436 28512
rect 4488 28500 4494 28552
rect 4801 28543 4859 28549
rect 4801 28509 4813 28543
rect 4847 28540 4859 28543
rect 5442 28540 5448 28552
rect 4847 28512 5448 28540
rect 4847 28509 4859 28512
rect 4801 28503 4859 28509
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 5902 28540 5908 28552
rect 5863 28512 5908 28540
rect 5902 28500 5908 28512
rect 5960 28500 5966 28552
rect 3418 28472 3424 28484
rect 3331 28444 3424 28472
rect 3344 28413 3372 28444
rect 3418 28432 3424 28444
rect 3476 28472 3482 28484
rect 4982 28472 4988 28484
rect 3476 28444 4988 28472
rect 3476 28432 3482 28444
rect 4982 28432 4988 28444
rect 5040 28432 5046 28484
rect 8128 28472 8156 28580
rect 8588 28580 9904 28608
rect 10003 28580 10048 28608
rect 8588 28549 8616 28580
rect 10042 28568 10048 28580
rect 10100 28568 10106 28620
rect 10321 28611 10379 28617
rect 10321 28577 10333 28611
rect 10367 28608 10379 28611
rect 10410 28608 10416 28620
rect 10367 28580 10416 28608
rect 10367 28577 10379 28580
rect 10321 28571 10379 28577
rect 10410 28568 10416 28580
rect 10468 28568 10474 28620
rect 10870 28568 10876 28620
rect 10928 28608 10934 28620
rect 12069 28611 12127 28617
rect 10928 28580 11652 28608
rect 10928 28568 10934 28580
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28509 8631 28543
rect 8573 28503 8631 28509
rect 9401 28543 9459 28549
rect 9401 28509 9413 28543
rect 9447 28540 9459 28543
rect 9950 28540 9956 28552
rect 9447 28512 9956 28540
rect 9447 28509 9459 28512
rect 9401 28503 9459 28509
rect 9950 28500 9956 28512
rect 10008 28500 10014 28552
rect 10594 28472 10600 28484
rect 5092 28444 6670 28472
rect 8128 28444 10600 28472
rect 3329 28407 3387 28413
rect 3329 28373 3341 28407
rect 3375 28373 3387 28407
rect 4246 28404 4252 28416
rect 4207 28376 4252 28404
rect 3329 28367 3387 28373
rect 4246 28364 4252 28376
rect 4304 28364 4310 28416
rect 4522 28364 4528 28416
rect 4580 28404 4586 28416
rect 5092 28404 5120 28444
rect 10594 28432 10600 28444
rect 10652 28432 10658 28484
rect 10778 28432 10784 28484
rect 10836 28432 10842 28484
rect 11624 28472 11652 28580
rect 12069 28577 12081 28611
rect 12115 28608 12127 28611
rect 13173 28611 13231 28617
rect 12115 28580 13124 28608
rect 12115 28577 12127 28580
rect 12069 28571 12127 28577
rect 11974 28500 11980 28552
rect 12032 28540 12038 28552
rect 12529 28543 12587 28549
rect 12529 28540 12541 28543
rect 12032 28512 12541 28540
rect 12032 28500 12038 28512
rect 12529 28509 12541 28512
rect 12575 28509 12587 28543
rect 12710 28540 12716 28552
rect 12671 28512 12716 28540
rect 12529 28503 12587 28509
rect 12710 28500 12716 28512
rect 12768 28500 12774 28552
rect 12342 28472 12348 28484
rect 11624 28444 12348 28472
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 13096 28472 13124 28580
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 17678 28608 17684 28620
rect 13219 28580 17684 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 17678 28568 17684 28580
rect 17736 28568 17742 28620
rect 17972 28608 18000 28639
rect 19536 28617 19564 28716
rect 24026 28704 24032 28716
rect 24084 28704 24090 28756
rect 21729 28679 21787 28685
rect 21729 28645 21741 28679
rect 21775 28676 21787 28679
rect 24578 28676 24584 28688
rect 21775 28648 24584 28676
rect 21775 28645 21787 28648
rect 21729 28639 21787 28645
rect 24578 28636 24584 28648
rect 24636 28636 24642 28688
rect 19521 28611 19579 28617
rect 17972 28580 18828 28608
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14424 28512 14749 28540
rect 14424 28500 14430 28512
rect 14737 28509 14749 28512
rect 14783 28540 14795 28543
rect 15010 28540 15016 28552
rect 14783 28512 15016 28540
rect 14783 28509 14795 28512
rect 14737 28503 14795 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 15749 28543 15807 28549
rect 15749 28540 15761 28543
rect 15528 28512 15761 28540
rect 15528 28500 15534 28512
rect 15749 28509 15761 28512
rect 15795 28509 15807 28543
rect 16850 28540 16856 28552
rect 16811 28512 16856 28540
rect 15749 28503 15807 28509
rect 16850 28500 16856 28512
rect 16908 28540 16914 28552
rect 17313 28543 17371 28549
rect 17313 28540 17325 28543
rect 16908 28512 17325 28540
rect 16908 28500 16914 28512
rect 17313 28509 17325 28512
rect 17359 28509 17371 28543
rect 17313 28503 17371 28509
rect 18046 28500 18052 28552
rect 18104 28540 18110 28552
rect 18800 28549 18828 28580
rect 19521 28577 19533 28611
rect 19567 28577 19579 28611
rect 19978 28608 19984 28620
rect 19939 28580 19984 28608
rect 19521 28571 19579 28577
rect 19978 28568 19984 28580
rect 20036 28568 20042 28620
rect 20254 28568 20260 28620
rect 20312 28608 20318 28620
rect 20625 28611 20683 28617
rect 20625 28608 20637 28611
rect 20312 28580 20637 28608
rect 20312 28568 20318 28580
rect 20625 28577 20637 28580
rect 20671 28577 20683 28611
rect 20806 28608 20812 28620
rect 20767 28580 20812 28608
rect 20625 28571 20683 28577
rect 20806 28568 20812 28580
rect 20864 28568 20870 28620
rect 22738 28608 22744 28620
rect 22699 28580 22744 28608
rect 22738 28568 22744 28580
rect 22796 28568 22802 28620
rect 22830 28568 22836 28620
rect 22888 28608 22894 28620
rect 22925 28611 22983 28617
rect 22925 28608 22937 28611
rect 22888 28580 22937 28608
rect 22888 28568 22894 28580
rect 22925 28577 22937 28580
rect 22971 28577 22983 28611
rect 22925 28571 22983 28577
rect 18141 28543 18199 28549
rect 18141 28540 18153 28543
rect 18104 28512 18153 28540
rect 18104 28500 18110 28512
rect 18141 28509 18153 28512
rect 18187 28509 18199 28543
rect 18141 28503 18199 28509
rect 18785 28543 18843 28549
rect 18785 28509 18797 28543
rect 18831 28509 18843 28543
rect 21910 28540 21916 28552
rect 21871 28512 21916 28540
rect 18785 28503 18843 28509
rect 21910 28500 21916 28512
rect 21968 28500 21974 28552
rect 17126 28472 17132 28484
rect 13096 28444 17132 28472
rect 17126 28432 17132 28444
rect 17184 28432 17190 28484
rect 17405 28475 17463 28481
rect 17405 28441 17417 28475
rect 17451 28472 17463 28475
rect 19613 28475 19671 28481
rect 17451 28444 19472 28472
rect 17451 28441 17463 28444
rect 17405 28435 17463 28441
rect 5442 28404 5448 28416
rect 4580 28376 5120 28404
rect 5403 28376 5448 28404
rect 4580 28364 4586 28376
rect 5442 28364 5448 28376
rect 5500 28364 5506 28416
rect 6822 28364 6828 28416
rect 6880 28404 6886 28416
rect 7926 28404 7932 28416
rect 6880 28376 7932 28404
rect 6880 28364 6886 28376
rect 7926 28364 7932 28376
rect 7984 28364 7990 28416
rect 9493 28407 9551 28413
rect 9493 28373 9505 28407
rect 9539 28404 9551 28407
rect 11882 28404 11888 28416
rect 9539 28376 11888 28404
rect 9539 28373 9551 28376
rect 9493 28367 9551 28373
rect 11882 28364 11888 28376
rect 11940 28364 11946 28416
rect 11974 28364 11980 28416
rect 12032 28404 12038 28416
rect 12894 28404 12900 28416
rect 12032 28376 12900 28404
rect 12032 28364 12038 28376
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 14829 28407 14887 28413
rect 14829 28373 14841 28407
rect 14875 28404 14887 28407
rect 15654 28404 15660 28416
rect 14875 28376 15660 28404
rect 14875 28373 14887 28376
rect 14829 28367 14887 28373
rect 15654 28364 15660 28376
rect 15712 28364 15718 28416
rect 15838 28404 15844 28416
rect 15799 28376 15844 28404
rect 15838 28364 15844 28376
rect 15896 28364 15902 28416
rect 18598 28404 18604 28416
rect 18559 28376 18604 28404
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 19444 28404 19472 28444
rect 19613 28441 19625 28475
rect 19659 28441 19671 28475
rect 19613 28435 19671 28441
rect 19628 28404 19656 28435
rect 19444 28376 19656 28404
rect 21082 28364 21088 28416
rect 21140 28404 21146 28416
rect 21269 28407 21327 28413
rect 21269 28404 21281 28407
rect 21140 28376 21281 28404
rect 21140 28364 21146 28376
rect 21269 28373 21281 28376
rect 21315 28373 21327 28407
rect 21269 28367 21327 28373
rect 23385 28407 23443 28413
rect 23385 28373 23397 28407
rect 23431 28404 23443 28407
rect 23658 28404 23664 28416
rect 23431 28376 23664 28404
rect 23431 28373 23443 28376
rect 23385 28367 23443 28373
rect 23658 28364 23664 28376
rect 23716 28364 23722 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 4246 28160 4252 28212
rect 4304 28200 4310 28212
rect 8110 28200 8116 28212
rect 4304 28172 8116 28200
rect 4304 28160 4310 28172
rect 8110 28160 8116 28172
rect 8168 28160 8174 28212
rect 8202 28160 8208 28212
rect 8260 28200 8266 28212
rect 10778 28200 10784 28212
rect 8260 28172 10784 28200
rect 8260 28160 8266 28172
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 11057 28203 11115 28209
rect 11057 28169 11069 28203
rect 11103 28200 11115 28203
rect 12710 28200 12716 28212
rect 11103 28172 12716 28200
rect 11103 28169 11115 28172
rect 11057 28163 11115 28169
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 12894 28160 12900 28212
rect 12952 28200 12958 28212
rect 13449 28203 13507 28209
rect 13449 28200 13461 28203
rect 12952 28172 13461 28200
rect 12952 28160 12958 28172
rect 13449 28169 13461 28172
rect 13495 28169 13507 28203
rect 13449 28163 13507 28169
rect 15010 28160 15016 28212
rect 15068 28200 15074 28212
rect 18506 28200 18512 28212
rect 15068 28172 18512 28200
rect 15068 28160 15074 28172
rect 18506 28160 18512 28172
rect 18564 28160 18570 28212
rect 20714 28160 20720 28212
rect 20772 28200 20778 28212
rect 20772 28172 20852 28200
rect 20772 28160 20778 28172
rect 1854 28132 1860 28144
rect 1815 28104 1860 28132
rect 1854 28092 1860 28104
rect 1912 28092 1918 28144
rect 4338 28132 4344 28144
rect 4299 28104 4344 28132
rect 4338 28092 4344 28104
rect 4396 28092 4402 28144
rect 4798 28092 4804 28144
rect 4856 28092 4862 28144
rect 6914 28092 6920 28144
rect 6972 28132 6978 28144
rect 9030 28132 9036 28144
rect 6972 28104 7774 28132
rect 8991 28104 9036 28132
rect 6972 28092 6978 28104
rect 9030 28092 9036 28104
rect 9088 28092 9094 28144
rect 9674 28092 9680 28144
rect 9732 28132 9738 28144
rect 9953 28135 10011 28141
rect 9953 28132 9965 28135
rect 9732 28104 9965 28132
rect 9732 28092 9738 28104
rect 9953 28101 9965 28104
rect 9999 28101 10011 28135
rect 9953 28095 10011 28101
rect 10042 28092 10048 28144
rect 10100 28132 10106 28144
rect 11974 28132 11980 28144
rect 10100 28104 11980 28132
rect 10100 28092 10106 28104
rect 11974 28092 11980 28104
rect 12032 28092 12038 28144
rect 13630 28132 13636 28144
rect 13202 28104 13636 28132
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 14700 28104 17540 28132
rect 14700 28092 14706 28104
rect 2958 28024 2964 28076
rect 3016 28024 3022 28076
rect 4062 28064 4068 28076
rect 3528 28036 4068 28064
rect 1578 27996 1584 28008
rect 1539 27968 1584 27996
rect 1578 27956 1584 27968
rect 1636 27996 1642 28008
rect 3528 27996 3556 28036
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 5902 28024 5908 28076
rect 5960 28064 5966 28076
rect 6822 28064 6828 28076
rect 5960 28036 6828 28064
rect 5960 28024 5966 28036
rect 6822 28024 6828 28036
rect 6880 28064 6886 28076
rect 7009 28067 7067 28073
rect 7009 28064 7021 28067
rect 6880 28036 7021 28064
rect 6880 28024 6886 28036
rect 7009 28033 7021 28036
rect 7055 28033 7067 28067
rect 7009 28027 7067 28033
rect 10686 28024 10692 28076
rect 10744 28064 10750 28076
rect 10965 28067 11023 28073
rect 10965 28064 10977 28067
rect 10744 28036 10977 28064
rect 10744 28024 10750 28036
rect 10965 28033 10977 28036
rect 11011 28033 11023 28067
rect 11698 28064 11704 28076
rect 11659 28036 11704 28064
rect 10965 28027 11023 28033
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 14369 28067 14427 28073
rect 14369 28033 14381 28067
rect 14415 28064 14427 28067
rect 14918 28064 14924 28076
rect 14415 28036 14924 28064
rect 14415 28033 14427 28036
rect 14369 28027 14427 28033
rect 14918 28024 14924 28036
rect 14976 28024 14982 28076
rect 15194 28064 15200 28076
rect 15155 28036 15200 28064
rect 15194 28024 15200 28036
rect 15252 28024 15258 28076
rect 15838 28064 15844 28076
rect 15799 28036 15844 28064
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 17405 28067 17463 28073
rect 17405 28064 17417 28067
rect 16816 28036 17417 28064
rect 16816 28024 16822 28036
rect 17405 28033 17417 28036
rect 17451 28033 17463 28067
rect 17512 28064 17540 28104
rect 18046 28092 18052 28144
rect 18104 28132 18110 28144
rect 20824 28141 20852 28172
rect 21634 28160 21640 28212
rect 21692 28200 21698 28212
rect 22649 28203 22707 28209
rect 22649 28200 22661 28203
rect 21692 28172 22661 28200
rect 21692 28160 21698 28172
rect 22649 28169 22661 28172
rect 22695 28169 22707 28203
rect 22649 28163 22707 28169
rect 20809 28135 20867 28141
rect 18104 28104 20116 28132
rect 18104 28092 18110 28104
rect 20088 28073 20116 28104
rect 20809 28101 20821 28135
rect 20855 28101 20867 28135
rect 20809 28095 20867 28101
rect 20901 28135 20959 28141
rect 20901 28101 20913 28135
rect 20947 28132 20959 28135
rect 23201 28135 23259 28141
rect 23201 28132 23213 28135
rect 20947 28104 23213 28132
rect 20947 28101 20959 28104
rect 20901 28095 20959 28101
rect 23201 28101 23213 28104
rect 23247 28101 23259 28135
rect 23201 28095 23259 28101
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 17512 28036 19625 28064
rect 17405 28027 17463 28033
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 20073 28067 20131 28073
rect 20073 28033 20085 28067
rect 20119 28033 20131 28067
rect 20073 28027 20131 28033
rect 1636 27968 3556 27996
rect 3605 27999 3663 28005
rect 1636 27956 1642 27968
rect 3605 27965 3617 27999
rect 3651 27996 3663 27999
rect 3786 27996 3792 28008
rect 3651 27968 3792 27996
rect 3651 27965 3663 27968
rect 3605 27959 3663 27965
rect 3786 27956 3792 27968
rect 3844 27956 3850 28008
rect 4430 27956 4436 28008
rect 4488 27996 4494 28008
rect 4798 27996 4804 28008
rect 4488 27968 4804 27996
rect 4488 27956 4494 27968
rect 4798 27956 4804 27968
rect 4856 27956 4862 28008
rect 5810 27996 5816 28008
rect 5771 27968 5816 27996
rect 5810 27956 5816 27968
rect 5868 27956 5874 28008
rect 7292 27999 7350 28005
rect 7292 27965 7304 27999
rect 7338 27996 7350 27999
rect 7650 27996 7656 28008
rect 7338 27968 7656 27996
rect 7338 27965 7350 27968
rect 7292 27959 7350 27965
rect 7650 27956 7656 27968
rect 7708 27956 7714 28008
rect 9861 27999 9919 28005
rect 9861 27965 9873 27999
rect 9907 27996 9919 27999
rect 10502 27996 10508 28008
rect 9907 27968 10508 27996
rect 9907 27965 9919 27968
rect 9861 27959 9919 27965
rect 10502 27956 10508 27968
rect 10560 27956 10566 28008
rect 11977 27999 12035 28005
rect 11977 27965 11989 27999
rect 12023 27996 12035 27999
rect 12342 27996 12348 28008
rect 12023 27968 12348 27996
rect 12023 27965 12035 27968
rect 11977 27959 12035 27965
rect 12342 27956 12348 27968
rect 12400 27996 12406 28008
rect 14458 27996 14464 28008
rect 12400 27968 14464 27996
rect 12400 27956 12406 27968
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 15657 27999 15715 28005
rect 15657 27965 15669 27999
rect 15703 27996 15715 27999
rect 16022 27996 16028 28008
rect 15703 27968 16028 27996
rect 15703 27965 15715 27968
rect 15657 27959 15715 27965
rect 16022 27956 16028 27968
rect 16080 27956 16086 28008
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27965 17279 27999
rect 18506 27996 18512 28008
rect 18467 27968 18512 27996
rect 17221 27959 17279 27965
rect 8570 27888 8576 27940
rect 8628 27928 8634 27940
rect 9306 27928 9312 27940
rect 8628 27900 9312 27928
rect 8628 27888 8634 27900
rect 9306 27888 9312 27900
rect 9364 27928 9370 27940
rect 10042 27928 10048 27940
rect 9364 27900 10048 27928
rect 9364 27888 9370 27900
rect 10042 27888 10048 27900
rect 10100 27888 10106 27940
rect 10413 27931 10471 27937
rect 10413 27897 10425 27931
rect 10459 27928 10471 27931
rect 11698 27928 11704 27940
rect 10459 27900 11704 27928
rect 10459 27897 10471 27900
rect 10413 27891 10471 27897
rect 11698 27888 11704 27900
rect 11756 27888 11762 27940
rect 13722 27888 13728 27940
rect 13780 27928 13786 27940
rect 15470 27928 15476 27940
rect 13780 27900 15476 27928
rect 13780 27888 13786 27900
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 17236 27928 17264 27959
rect 18506 27956 18512 27968
rect 18564 27956 18570 28008
rect 19628 27996 19656 28027
rect 21818 28024 21824 28076
rect 21876 28064 21882 28076
rect 22005 28067 22063 28073
rect 22005 28064 22017 28067
rect 21876 28036 22017 28064
rect 21876 28024 21882 28036
rect 22005 28033 22017 28036
rect 22051 28033 22063 28067
rect 22186 28064 22192 28076
rect 22147 28036 22192 28064
rect 22005 28027 22063 28033
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 23109 28067 23167 28073
rect 23109 28033 23121 28067
rect 23155 28033 23167 28067
rect 24946 28064 24952 28076
rect 24907 28036 24952 28064
rect 23109 28027 23167 28033
rect 20346 27996 20352 28008
rect 19628 27968 20352 27996
rect 20346 27956 20352 27968
rect 20404 27956 20410 28008
rect 21453 27999 21511 28005
rect 21453 27965 21465 27999
rect 21499 27996 21511 27999
rect 21726 27996 21732 28008
rect 21499 27968 21732 27996
rect 21499 27965 21511 27968
rect 21453 27959 21511 27965
rect 21726 27956 21732 27968
rect 21784 27956 21790 28008
rect 20990 27928 20996 27940
rect 17236 27900 20996 27928
rect 20990 27888 20996 27900
rect 21048 27888 21054 27940
rect 21910 27888 21916 27940
rect 21968 27928 21974 27940
rect 23124 27928 23152 28027
rect 24946 28024 24952 28036
rect 25004 28024 25010 28076
rect 23474 27956 23480 28008
rect 23532 27996 23538 28008
rect 23753 27999 23811 28005
rect 23753 27996 23765 27999
rect 23532 27968 23765 27996
rect 23532 27956 23538 27968
rect 23753 27965 23765 27968
rect 23799 27965 23811 27999
rect 23753 27959 23811 27965
rect 21968 27900 23152 27928
rect 21968 27888 21974 27900
rect 5442 27820 5448 27872
rect 5500 27860 5506 27872
rect 8662 27860 8668 27872
rect 5500 27832 8668 27860
rect 5500 27820 5506 27832
rect 8662 27820 8668 27832
rect 8720 27820 8726 27872
rect 9398 27820 9404 27872
rect 9456 27860 9462 27872
rect 14366 27860 14372 27872
rect 9456 27832 14372 27860
rect 9456 27820 9462 27832
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 14461 27863 14519 27869
rect 14461 27829 14473 27863
rect 14507 27860 14519 27863
rect 14642 27860 14648 27872
rect 14507 27832 14648 27860
rect 14507 27829 14519 27832
rect 14461 27823 14519 27829
rect 14642 27820 14648 27832
rect 14700 27820 14706 27872
rect 15013 27863 15071 27869
rect 15013 27829 15025 27863
rect 15059 27860 15071 27863
rect 15746 27860 15752 27872
rect 15059 27832 15752 27860
rect 15059 27829 15071 27832
rect 15013 27823 15071 27829
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 16301 27863 16359 27869
rect 16301 27829 16313 27863
rect 16347 27860 16359 27863
rect 16574 27860 16580 27872
rect 16347 27832 16580 27860
rect 16347 27829 16359 27832
rect 16301 27823 16359 27829
rect 16574 27820 16580 27832
rect 16632 27820 16638 27872
rect 17494 27820 17500 27872
rect 17552 27860 17558 27872
rect 17589 27863 17647 27869
rect 17589 27860 17601 27863
rect 17552 27832 17601 27860
rect 17552 27820 17558 27832
rect 17589 27829 17601 27832
rect 17635 27829 17647 27863
rect 17589 27823 17647 27829
rect 19429 27863 19487 27869
rect 19429 27829 19441 27863
rect 19475 27860 19487 27863
rect 19610 27860 19616 27872
rect 19475 27832 19616 27860
rect 19475 27829 19487 27832
rect 19429 27823 19487 27829
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 20165 27863 20223 27869
rect 20165 27829 20177 27863
rect 20211 27860 20223 27863
rect 22186 27860 22192 27872
rect 20211 27832 22192 27860
rect 20211 27829 20223 27832
rect 20165 27823 20223 27829
rect 22186 27820 22192 27832
rect 22244 27820 22250 27872
rect 24762 27860 24768 27872
rect 24723 27832 24768 27860
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1854 27665 1860 27668
rect 1844 27659 1860 27665
rect 1844 27625 1856 27659
rect 1844 27619 1860 27625
rect 1854 27616 1860 27619
rect 1912 27616 1918 27668
rect 5432 27659 5490 27665
rect 5432 27625 5444 27659
rect 5478 27656 5490 27659
rect 8754 27656 8760 27668
rect 5478 27628 8760 27656
rect 5478 27625 5490 27628
rect 5432 27619 5490 27625
rect 8754 27616 8760 27628
rect 8812 27616 8818 27668
rect 10873 27659 10931 27665
rect 10873 27625 10885 27659
rect 10919 27656 10931 27659
rect 10962 27656 10968 27668
rect 10919 27628 10968 27656
rect 10919 27625 10931 27628
rect 10873 27619 10931 27625
rect 10962 27616 10968 27628
rect 11020 27656 11026 27668
rect 11238 27656 11244 27668
rect 11020 27628 11244 27656
rect 11020 27616 11026 27628
rect 11238 27616 11244 27628
rect 11296 27616 11302 27668
rect 11698 27616 11704 27668
rect 11756 27656 11762 27668
rect 13538 27656 13544 27668
rect 11756 27628 13544 27656
rect 11756 27616 11762 27628
rect 13538 27616 13544 27628
rect 13596 27616 13602 27668
rect 15286 27656 15292 27668
rect 14844 27628 15292 27656
rect 4062 27548 4068 27600
rect 4120 27548 4126 27600
rect 4709 27591 4767 27597
rect 4709 27557 4721 27591
rect 4755 27588 4767 27591
rect 4890 27588 4896 27600
rect 4755 27560 4896 27588
rect 4755 27557 4767 27560
rect 4709 27551 4767 27557
rect 4890 27548 4896 27560
rect 4948 27548 4954 27600
rect 8573 27591 8631 27597
rect 8573 27557 8585 27591
rect 8619 27588 8631 27591
rect 8662 27588 8668 27600
rect 8619 27560 8668 27588
rect 8619 27557 8631 27560
rect 8573 27551 8631 27557
rect 8662 27548 8668 27560
rect 8720 27548 8726 27600
rect 14844 27588 14872 27628
rect 15286 27616 15292 27628
rect 15344 27616 15350 27668
rect 18138 27588 18144 27600
rect 10520 27560 14872 27588
rect 15580 27560 18144 27588
rect 4080 27520 4108 27548
rect 5169 27523 5227 27529
rect 5169 27520 5181 27523
rect 4080 27492 5181 27520
rect 5169 27489 5181 27492
rect 5215 27520 5227 27523
rect 5902 27520 5908 27532
rect 5215 27492 5908 27520
rect 5215 27489 5227 27492
rect 5169 27483 5227 27489
rect 5902 27480 5908 27492
rect 5960 27480 5966 27532
rect 6822 27480 6828 27532
rect 6880 27520 6886 27532
rect 9122 27520 9128 27532
rect 6880 27492 9128 27520
rect 6880 27480 6886 27492
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 9398 27520 9404 27532
rect 9359 27492 9404 27520
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 3142 27412 3148 27464
rect 3200 27452 3206 27464
rect 4065 27455 4123 27461
rect 4065 27452 4077 27455
rect 3200 27424 4077 27452
rect 3200 27412 3206 27424
rect 4065 27421 4077 27424
rect 4111 27421 4123 27455
rect 4065 27415 4123 27421
rect 4249 27455 4307 27461
rect 4249 27421 4261 27455
rect 4295 27452 4307 27455
rect 4890 27452 4896 27464
rect 4295 27424 4896 27452
rect 4295 27421 4307 27424
rect 4249 27415 4307 27421
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 7193 27455 7251 27461
rect 7193 27421 7205 27455
rect 7239 27452 7251 27455
rect 7466 27452 7472 27464
rect 7239 27424 7472 27452
rect 7239 27421 7251 27424
rect 7193 27415 7251 27421
rect 7466 27412 7472 27424
rect 7524 27452 7530 27464
rect 7650 27452 7656 27464
rect 7524 27424 7656 27452
rect 7524 27412 7530 27424
rect 7650 27412 7656 27424
rect 7708 27412 7714 27464
rect 7926 27452 7932 27464
rect 7887 27424 7932 27452
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 8110 27452 8116 27464
rect 8071 27424 8116 27452
rect 8110 27412 8116 27424
rect 8168 27412 8174 27464
rect 8846 27412 8852 27464
rect 8904 27452 8910 27464
rect 8904 27424 9168 27452
rect 10520 27438 10548 27560
rect 11517 27523 11575 27529
rect 11517 27489 11529 27523
rect 11563 27520 11575 27523
rect 13906 27520 13912 27532
rect 11563 27492 13912 27520
rect 11563 27489 11575 27492
rect 11517 27483 11575 27489
rect 13906 27480 13912 27492
rect 13964 27480 13970 27532
rect 15013 27523 15071 27529
rect 15013 27489 15025 27523
rect 15059 27520 15071 27523
rect 15580 27520 15608 27560
rect 18138 27548 18144 27560
rect 18196 27548 18202 27600
rect 19978 27548 19984 27600
rect 20036 27588 20042 27600
rect 20717 27591 20775 27597
rect 20717 27588 20729 27591
rect 20036 27560 20729 27588
rect 20036 27548 20042 27560
rect 20717 27557 20729 27560
rect 20763 27557 20775 27591
rect 21634 27588 21640 27600
rect 21595 27560 21640 27588
rect 20717 27551 20775 27557
rect 21634 27548 21640 27560
rect 21692 27548 21698 27600
rect 22738 27588 22744 27600
rect 22699 27560 22744 27588
rect 22738 27548 22744 27560
rect 22796 27588 22802 27600
rect 23382 27588 23388 27600
rect 22796 27560 23388 27588
rect 22796 27548 22802 27560
rect 23382 27548 23388 27560
rect 23440 27548 23446 27600
rect 15059 27492 15608 27520
rect 15059 27489 15071 27492
rect 15013 27483 15071 27489
rect 15654 27480 15660 27532
rect 15712 27520 15718 27532
rect 16301 27523 16359 27529
rect 16301 27520 16313 27523
rect 15712 27492 16313 27520
rect 15712 27480 15718 27492
rect 16301 27489 16313 27492
rect 16347 27489 16359 27523
rect 16301 27483 16359 27489
rect 18417 27523 18475 27529
rect 18417 27489 18429 27523
rect 18463 27520 18475 27523
rect 18598 27520 18604 27532
rect 18463 27492 18604 27520
rect 18463 27489 18475 27492
rect 18417 27483 18475 27489
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 20165 27523 20223 27529
rect 20165 27489 20177 27523
rect 20211 27520 20223 27523
rect 20211 27492 21588 27520
rect 20211 27489 20223 27492
rect 20165 27483 20223 27489
rect 14458 27452 14464 27464
rect 14419 27424 14464 27452
rect 8904 27412 8910 27424
rect 4614 27384 4620 27396
rect 3082 27356 4620 27384
rect 4614 27344 4620 27356
rect 4672 27344 4678 27396
rect 6730 27384 6736 27396
rect 6670 27356 6736 27384
rect 6730 27344 6736 27356
rect 6788 27344 6794 27396
rect 7558 27344 7564 27396
rect 7616 27384 7622 27396
rect 8938 27384 8944 27396
rect 7616 27356 8944 27384
rect 7616 27344 7622 27356
rect 8938 27344 8944 27356
rect 8996 27344 9002 27396
rect 9140 27384 9168 27424
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27421 16175 27455
rect 16117 27415 16175 27421
rect 9306 27384 9312 27396
rect 9140 27356 9312 27384
rect 9306 27344 9312 27356
rect 9364 27344 9370 27396
rect 11054 27344 11060 27396
rect 11112 27384 11118 27396
rect 11609 27387 11667 27393
rect 11609 27384 11621 27387
rect 11112 27356 11621 27384
rect 11112 27344 11118 27356
rect 11609 27353 11621 27356
rect 11655 27353 11667 27387
rect 11609 27347 11667 27353
rect 11698 27344 11704 27396
rect 11756 27384 11762 27396
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 11756 27356 12173 27384
rect 11756 27344 11762 27356
rect 12161 27353 12173 27356
rect 12207 27353 12219 27387
rect 12161 27347 12219 27353
rect 12710 27344 12716 27396
rect 12768 27384 12774 27396
rect 12897 27387 12955 27393
rect 12897 27384 12909 27387
rect 12768 27356 12909 27384
rect 12768 27344 12774 27356
rect 12897 27353 12909 27356
rect 12943 27353 12955 27387
rect 12897 27347 12955 27353
rect 12986 27344 12992 27396
rect 13044 27384 13050 27396
rect 13541 27387 13599 27393
rect 13044 27356 13089 27384
rect 13044 27344 13050 27356
rect 13541 27353 13553 27387
rect 13587 27384 13599 27387
rect 13587 27356 14872 27384
rect 13587 27353 13599 27356
rect 13541 27347 13599 27353
rect 14844 27328 14872 27356
rect 15102 27344 15108 27396
rect 15160 27384 15166 27396
rect 15657 27387 15715 27393
rect 15160 27356 15205 27384
rect 15160 27344 15166 27356
rect 15657 27353 15669 27387
rect 15703 27353 15715 27387
rect 16132 27384 16160 27415
rect 16206 27412 16212 27464
rect 16264 27452 16270 27464
rect 17773 27455 17831 27461
rect 17773 27452 17785 27455
rect 16264 27424 17785 27452
rect 16264 27412 16270 27424
rect 17773 27421 17785 27424
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 17862 27412 17868 27464
rect 17920 27452 17926 27464
rect 18233 27455 18291 27461
rect 18233 27452 18245 27455
rect 17920 27424 18245 27452
rect 17920 27412 17926 27424
rect 18233 27421 18245 27424
rect 18279 27452 18291 27455
rect 18782 27452 18788 27464
rect 18279 27424 18788 27452
rect 18279 27421 18291 27424
rect 18233 27415 18291 27421
rect 18782 27412 18788 27424
rect 18840 27412 18846 27464
rect 19610 27452 19616 27464
rect 19571 27424 19616 27452
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 21266 27452 21272 27464
rect 21227 27424 21272 27452
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21453 27455 21511 27461
rect 21453 27421 21465 27455
rect 21499 27421 21511 27455
rect 21560 27452 21588 27492
rect 22002 27480 22008 27532
rect 22060 27520 22066 27532
rect 22557 27523 22615 27529
rect 22557 27520 22569 27523
rect 22060 27492 22569 27520
rect 22060 27480 22066 27492
rect 22557 27489 22569 27492
rect 22603 27489 22615 27523
rect 22557 27483 22615 27489
rect 22373 27455 22431 27461
rect 21560 27424 22094 27452
rect 21453 27415 21511 27421
rect 18690 27384 18696 27396
rect 16132 27356 18696 27384
rect 15657 27347 15715 27353
rect 3329 27319 3387 27325
rect 3329 27285 3341 27319
rect 3375 27316 3387 27319
rect 3418 27316 3424 27328
rect 3375 27288 3424 27316
rect 3375 27285 3387 27288
rect 3329 27279 3387 27285
rect 3418 27276 3424 27288
rect 3476 27276 3482 27328
rect 5350 27276 5356 27328
rect 5408 27316 5414 27328
rect 10318 27316 10324 27328
rect 5408 27288 10324 27316
rect 5408 27276 5414 27288
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 13170 27276 13176 27328
rect 13228 27316 13234 27328
rect 14277 27319 14335 27325
rect 14277 27316 14289 27319
rect 13228 27288 14289 27316
rect 13228 27276 13234 27288
rect 14277 27285 14289 27288
rect 14323 27285 14335 27319
rect 14277 27279 14335 27285
rect 14826 27276 14832 27328
rect 14884 27316 14890 27328
rect 15672 27316 15700 27347
rect 18690 27344 18696 27356
rect 18748 27384 18754 27396
rect 18877 27387 18935 27393
rect 18877 27384 18889 27387
rect 18748 27356 18889 27384
rect 18748 27344 18754 27356
rect 18877 27353 18889 27356
rect 18923 27353 18935 27387
rect 18877 27347 18935 27353
rect 19242 27344 19248 27396
rect 19300 27384 19306 27396
rect 20257 27387 20315 27393
rect 20257 27384 20269 27387
rect 19300 27356 20269 27384
rect 19300 27344 19306 27356
rect 20257 27353 20269 27356
rect 20303 27353 20315 27387
rect 20257 27347 20315 27353
rect 16758 27316 16764 27328
rect 14884 27288 15700 27316
rect 16719 27288 16764 27316
rect 14884 27276 14890 27288
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 17589 27319 17647 27325
rect 17589 27285 17601 27319
rect 17635 27316 17647 27319
rect 19058 27316 19064 27328
rect 17635 27288 19064 27316
rect 17635 27285 17647 27288
rect 17589 27279 17647 27285
rect 19058 27276 19064 27288
rect 19116 27276 19122 27328
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 21468 27316 21496 27415
rect 22066 27384 22094 27424
rect 22373 27421 22385 27455
rect 22419 27452 22431 27455
rect 23474 27452 23480 27464
rect 22419 27424 23480 27452
rect 22419 27421 22431 27424
rect 22373 27415 22431 27421
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 23661 27455 23719 27461
rect 23661 27452 23673 27455
rect 23624 27424 23673 27452
rect 23624 27412 23630 27424
rect 23661 27421 23673 27424
rect 23707 27452 23719 27455
rect 24210 27452 24216 27464
rect 23707 27424 24216 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24210 27412 24216 27424
rect 24268 27412 24274 27464
rect 24302 27412 24308 27464
rect 24360 27452 24366 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24360 27424 24593 27452
rect 24360 27412 24366 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 31665 27455 31723 27461
rect 31665 27421 31677 27455
rect 31711 27452 31723 27455
rect 35434 27452 35440 27464
rect 31711 27424 35440 27452
rect 31711 27421 31723 27424
rect 31665 27415 31723 27421
rect 35434 27412 35440 27424
rect 35492 27412 35498 27464
rect 38010 27452 38016 27464
rect 37971 27424 38016 27452
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 23934 27384 23940 27396
rect 22066 27356 23940 27384
rect 23934 27344 23940 27356
rect 23992 27344 23998 27396
rect 19475 27288 21496 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 21542 27276 21548 27328
rect 21600 27316 21606 27328
rect 23290 27316 23296 27328
rect 21600 27288 23296 27316
rect 21600 27276 21606 27288
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 23474 27316 23480 27328
rect 23435 27288 23480 27316
rect 23474 27276 23480 27288
rect 23532 27276 23538 27328
rect 23566 27276 23572 27328
rect 23624 27316 23630 27328
rect 24673 27319 24731 27325
rect 24673 27316 24685 27319
rect 23624 27288 24685 27316
rect 23624 27276 23630 27288
rect 24673 27285 24685 27288
rect 24719 27285 24731 27319
rect 31754 27316 31760 27328
rect 31715 27288 31760 27316
rect 24673 27279 24731 27285
rect 31754 27276 31760 27288
rect 31812 27276 31818 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1762 27112 1768 27124
rect 1723 27084 1768 27112
rect 1762 27072 1768 27084
rect 1820 27072 1826 27124
rect 2777 27115 2835 27121
rect 2777 27081 2789 27115
rect 2823 27112 2835 27115
rect 3142 27112 3148 27124
rect 2823 27084 3148 27112
rect 2823 27081 2835 27084
rect 2777 27075 2835 27081
rect 3142 27072 3148 27084
rect 3200 27072 3206 27124
rect 5813 27115 5871 27121
rect 5813 27081 5825 27115
rect 5859 27112 5871 27115
rect 9674 27112 9680 27124
rect 5859 27084 9680 27112
rect 5859 27081 5871 27084
rect 5813 27075 5871 27081
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 11698 27112 11704 27124
rect 9876 27084 11704 27112
rect 3602 27044 3608 27056
rect 3563 27016 3608 27044
rect 3602 27004 3608 27016
rect 3660 27004 3666 27056
rect 5350 27044 5356 27056
rect 5311 27016 5356 27044
rect 5350 27004 5356 27016
rect 5408 27004 5414 27056
rect 5718 27004 5724 27056
rect 5776 27044 5782 27056
rect 5776 27016 7774 27044
rect 5776 27004 5782 27016
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 9876 27044 9904 27084
rect 11698 27072 11704 27084
rect 11756 27072 11762 27124
rect 14829 27115 14887 27121
rect 11808 27084 14780 27112
rect 11514 27044 11520 27056
rect 8996 27016 9904 27044
rect 10718 27016 11520 27044
rect 8996 27004 9002 27016
rect 11514 27004 11520 27016
rect 11572 27004 11578 27056
rect 11808 27053 11836 27084
rect 11793 27047 11851 27053
rect 11793 27013 11805 27047
rect 11839 27013 11851 27047
rect 11793 27007 11851 27013
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 11940 27016 11985 27044
rect 12912 27016 13584 27044
rect 11940 27004 11946 27016
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26976 1639 26979
rect 1946 26976 1952 26988
rect 1627 26948 1952 26976
rect 1627 26945 1639 26948
rect 1581 26939 1639 26945
rect 1946 26936 1952 26948
rect 2004 26936 2010 26988
rect 2590 26976 2596 26988
rect 2551 26948 2596 26976
rect 2590 26936 2596 26948
rect 2648 26936 2654 26988
rect 4706 26936 4712 26988
rect 4764 26936 4770 26988
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26976 6055 26979
rect 6086 26976 6092 26988
rect 6043 26948 6092 26976
rect 6043 26945 6055 26948
rect 5997 26939 6055 26945
rect 6086 26936 6092 26948
rect 6144 26936 6150 26988
rect 6822 26936 6828 26988
rect 6880 26976 6886 26988
rect 7009 26979 7067 26985
rect 7009 26976 7021 26979
rect 6880 26948 7021 26976
rect 6880 26936 6886 26948
rect 7009 26945 7021 26948
rect 7055 26945 7067 26979
rect 7009 26939 7067 26945
rect 9122 26936 9128 26988
rect 9180 26976 9186 26988
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 9180 26948 9229 26976
rect 9180 26936 9186 26948
rect 9217 26945 9229 26948
rect 9263 26945 9275 26979
rect 12912 26976 12940 27016
rect 13556 26985 13584 27016
rect 14550 27004 14556 27056
rect 14608 27044 14614 27056
rect 14752 27044 14780 27084
rect 14829 27081 14841 27115
rect 14875 27112 14887 27115
rect 17494 27112 17500 27124
rect 14875 27084 17500 27112
rect 14875 27081 14887 27084
rect 14829 27075 14887 27081
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 18690 27112 18696 27124
rect 18651 27084 18696 27112
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 18782 27072 18788 27124
rect 18840 27112 18846 27124
rect 21542 27112 21548 27124
rect 18840 27084 21548 27112
rect 18840 27072 18846 27084
rect 21542 27072 21548 27084
rect 21600 27072 21606 27124
rect 25133 27115 25191 27121
rect 25133 27081 25145 27115
rect 25179 27112 25191 27115
rect 25314 27112 25320 27124
rect 25179 27084 25320 27112
rect 25179 27081 25191 27084
rect 25133 27075 25191 27081
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 29181 27115 29239 27121
rect 29181 27081 29193 27115
rect 29227 27112 29239 27115
rect 34422 27112 34428 27124
rect 29227 27084 34428 27112
rect 29227 27081 29239 27084
rect 29181 27075 29239 27081
rect 34422 27072 34428 27084
rect 34480 27072 34486 27124
rect 15654 27044 15660 27056
rect 14608 27016 14688 27044
rect 14752 27016 15660 27044
rect 14608 27004 14614 27016
rect 9217 26939 9275 26945
rect 12452 26948 12940 26976
rect 13081 26979 13139 26985
rect 13081 26966 13093 26979
rect 1670 26868 1676 26920
rect 1728 26908 1734 26920
rect 3329 26911 3387 26917
rect 3329 26908 3341 26911
rect 1728 26880 3341 26908
rect 1728 26868 1734 26880
rect 3329 26877 3341 26880
rect 3375 26877 3387 26911
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 3329 26871 3387 26877
rect 7024 26880 7297 26908
rect 7024 26852 7052 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 9493 26911 9551 26917
rect 9493 26908 9505 26911
rect 8628 26880 9505 26908
rect 8628 26868 8634 26880
rect 9493 26877 9505 26880
rect 9539 26877 9551 26911
rect 9493 26871 9551 26877
rect 11238 26868 11244 26920
rect 11296 26908 11302 26920
rect 12452 26908 12480 26948
rect 13004 26945 13093 26966
rect 13127 26945 13139 26979
rect 13004 26939 13139 26945
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26976 13599 26979
rect 13722 26976 13728 26988
rect 13587 26948 13728 26976
rect 13587 26945 13599 26948
rect 13541 26939 13599 26945
rect 13004 26938 13124 26939
rect 11296 26880 12480 26908
rect 11296 26868 11302 26880
rect 12526 26868 12532 26920
rect 12584 26908 12590 26920
rect 13004 26908 13032 26938
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 14274 26936 14280 26988
rect 14332 26976 14338 26988
rect 14369 26979 14427 26985
rect 14369 26976 14381 26979
rect 14332 26948 14381 26976
rect 14332 26936 14338 26948
rect 14369 26945 14381 26948
rect 14415 26945 14427 26979
rect 14369 26939 14427 26945
rect 12584 26880 13032 26908
rect 14185 26911 14243 26917
rect 12584 26868 12590 26880
rect 14185 26877 14197 26911
rect 14231 26908 14243 26911
rect 14550 26908 14556 26920
rect 14231 26880 14556 26908
rect 14231 26877 14243 26880
rect 14185 26871 14243 26877
rect 14550 26868 14556 26880
rect 14608 26868 14614 26920
rect 14660 26908 14688 27016
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 15746 27004 15752 27056
rect 15804 27004 15810 27056
rect 16666 27004 16672 27056
rect 16724 27044 16730 27056
rect 16724 27016 18092 27044
rect 16724 27004 16730 27016
rect 14826 26908 14832 26920
rect 14660 26880 14832 26908
rect 14826 26868 14832 26880
rect 14884 26868 14890 26920
rect 15470 26868 15476 26920
rect 15528 26908 15534 26920
rect 15657 26911 15715 26917
rect 15657 26908 15669 26911
rect 15528 26880 15669 26908
rect 15528 26868 15534 26880
rect 15657 26877 15669 26880
rect 15703 26877 15715 26911
rect 15764 26908 15792 27004
rect 17402 26976 17408 26988
rect 17363 26948 17408 26976
rect 17402 26936 17408 26948
rect 17460 26936 17466 26988
rect 18064 26976 18092 27016
rect 21818 27004 21824 27056
rect 21876 27044 21882 27056
rect 21876 27016 22094 27044
rect 21876 27004 21882 27016
rect 18322 26976 18328 26988
rect 18064 26948 18328 26976
rect 18064 26917 18092 26948
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 19058 26936 19064 26988
rect 19116 26976 19122 26988
rect 19797 26979 19855 26985
rect 19797 26976 19809 26979
rect 19116 26948 19809 26976
rect 19116 26936 19122 26948
rect 19797 26945 19809 26948
rect 19843 26945 19855 26979
rect 22066 26976 22094 27016
rect 22830 27004 22836 27056
rect 22888 27044 22894 27056
rect 22888 27016 29132 27044
rect 22888 27004 22894 27016
rect 23109 26979 23167 26985
rect 23109 26976 23121 26979
rect 22066 26948 23121 26976
rect 19797 26939 19855 26945
rect 23109 26945 23121 26948
rect 23155 26945 23167 26979
rect 23109 26939 23167 26945
rect 24673 26979 24731 26985
rect 24673 26945 24685 26979
rect 24719 26976 24731 26979
rect 24762 26976 24768 26988
rect 24719 26948 24768 26976
rect 24719 26945 24731 26948
rect 24673 26939 24731 26945
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 29104 26985 29132 27016
rect 29089 26979 29147 26985
rect 29089 26945 29101 26979
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 32493 26979 32551 26985
rect 32493 26945 32505 26979
rect 32539 26976 32551 26979
rect 36998 26976 37004 26988
rect 32539 26948 37004 26976
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 36998 26936 37004 26948
rect 37056 26936 37062 26988
rect 15841 26911 15899 26917
rect 15841 26908 15853 26911
rect 15764 26880 15853 26908
rect 15657 26871 15715 26877
rect 15841 26877 15853 26880
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 18049 26911 18107 26917
rect 18049 26877 18061 26911
rect 18095 26877 18107 26911
rect 18230 26908 18236 26920
rect 18191 26880 18236 26908
rect 18049 26871 18107 26877
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 20254 26908 20260 26920
rect 20215 26880 20260 26908
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 20714 26868 20720 26920
rect 20772 26908 20778 26920
rect 20901 26911 20959 26917
rect 20901 26908 20913 26911
rect 20772 26880 20913 26908
rect 20772 26868 20778 26880
rect 20901 26877 20913 26880
rect 20947 26877 20959 26911
rect 20901 26871 20959 26877
rect 22005 26911 22063 26917
rect 22005 26877 22017 26911
rect 22051 26877 22063 26911
rect 22186 26908 22192 26920
rect 22147 26880 22192 26908
rect 22005 26871 22063 26877
rect 7006 26800 7012 26852
rect 7064 26800 7070 26852
rect 12158 26840 12164 26852
rect 8312 26812 8892 26840
rect 5718 26732 5724 26784
rect 5776 26772 5782 26784
rect 8312 26772 8340 26812
rect 8754 26772 8760 26784
rect 5776 26744 8340 26772
rect 8715 26744 8760 26772
rect 5776 26732 5782 26744
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 8864 26772 8892 26812
rect 10520 26812 12164 26840
rect 10520 26772 10548 26812
rect 12158 26800 12164 26812
rect 12216 26800 12222 26852
rect 12250 26800 12256 26852
rect 12308 26840 12314 26852
rect 12345 26843 12403 26849
rect 12345 26840 12357 26843
rect 12308 26812 12357 26840
rect 12308 26800 12314 26812
rect 12345 26809 12357 26812
rect 12391 26809 12403 26843
rect 12345 26803 12403 26809
rect 12728 26812 13032 26840
rect 10962 26772 10968 26784
rect 8864 26744 10548 26772
rect 10923 26744 10968 26772
rect 10962 26732 10968 26744
rect 11020 26772 11026 26784
rect 12728 26772 12756 26812
rect 12894 26772 12900 26784
rect 11020 26744 12756 26772
rect 12855 26744 12900 26772
rect 11020 26732 11026 26744
rect 12894 26732 12900 26744
rect 12952 26732 12958 26784
rect 13004 26772 13032 26812
rect 13464 26812 13952 26840
rect 13464 26772 13492 26812
rect 13630 26772 13636 26784
rect 13004 26744 13492 26772
rect 13591 26744 13636 26772
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 13924 26772 13952 26812
rect 13998 26800 14004 26852
rect 14056 26840 14062 26852
rect 16025 26843 16083 26849
rect 16025 26840 16037 26843
rect 14056 26812 16037 26840
rect 14056 26800 14062 26812
rect 16025 26809 16037 26812
rect 16071 26840 16083 26843
rect 16758 26840 16764 26852
rect 16071 26812 16764 26840
rect 16071 26809 16083 26812
rect 16025 26803 16083 26809
rect 16758 26800 16764 26812
rect 16816 26800 16822 26852
rect 17586 26800 17592 26852
rect 17644 26840 17650 26852
rect 19978 26840 19984 26852
rect 17644 26812 19984 26840
rect 17644 26800 17650 26812
rect 19978 26800 19984 26812
rect 20036 26840 20042 26852
rect 22020 26840 22048 26871
rect 22186 26868 22192 26880
rect 22244 26868 22250 26920
rect 23290 26908 23296 26920
rect 23251 26880 23296 26908
rect 23290 26868 23296 26880
rect 23348 26868 23354 26920
rect 24486 26908 24492 26920
rect 24447 26880 24492 26908
rect 24486 26868 24492 26880
rect 24544 26868 24550 26920
rect 31754 26840 31760 26852
rect 20036 26812 21036 26840
rect 22020 26812 31760 26840
rect 20036 26800 20042 26812
rect 17310 26772 17316 26784
rect 13924 26744 17316 26772
rect 17310 26732 17316 26744
rect 17368 26732 17374 26784
rect 17494 26772 17500 26784
rect 17455 26744 17500 26772
rect 17494 26732 17500 26744
rect 17552 26732 17558 26784
rect 19613 26775 19671 26781
rect 19613 26741 19625 26775
rect 19659 26772 19671 26775
rect 20898 26772 20904 26784
rect 19659 26744 20904 26772
rect 19659 26741 19671 26744
rect 19613 26735 19671 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 21008 26772 21036 26812
rect 31754 26800 31760 26812
rect 31812 26800 31818 26852
rect 22373 26775 22431 26781
rect 22373 26772 22385 26775
rect 21008 26744 22385 26772
rect 22373 26741 22385 26744
rect 22419 26741 22431 26775
rect 22373 26735 22431 26741
rect 23753 26775 23811 26781
rect 23753 26741 23765 26775
rect 23799 26772 23811 26775
rect 24026 26772 24032 26784
rect 23799 26744 24032 26772
rect 23799 26741 23811 26744
rect 23753 26735 23811 26741
rect 24026 26732 24032 26744
rect 24084 26732 24090 26784
rect 32582 26772 32588 26784
rect 32543 26744 32588 26772
rect 32582 26732 32588 26744
rect 32640 26732 32646 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1844 26571 1902 26577
rect 1844 26537 1856 26571
rect 1890 26568 1902 26571
rect 5718 26568 5724 26580
rect 1890 26540 5724 26568
rect 1890 26537 1902 26540
rect 1844 26531 1902 26537
rect 5718 26528 5724 26540
rect 5776 26528 5782 26580
rect 7088 26571 7146 26577
rect 7088 26537 7100 26571
rect 7134 26568 7146 26571
rect 10962 26568 10968 26580
rect 7134 26540 10968 26568
rect 7134 26537 7146 26540
rect 7088 26531 7146 26537
rect 10962 26528 10968 26540
rect 11020 26528 11026 26580
rect 11609 26571 11667 26577
rect 11609 26537 11621 26571
rect 11655 26568 11667 26571
rect 12526 26568 12532 26580
rect 11655 26540 12532 26568
rect 11655 26537 11667 26540
rect 11609 26531 11667 26537
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 15105 26571 15163 26577
rect 15105 26537 15117 26571
rect 15151 26568 15163 26571
rect 18414 26568 18420 26580
rect 15151 26540 18420 26568
rect 15151 26537 15163 26540
rect 15105 26531 15163 26537
rect 18414 26528 18420 26540
rect 18472 26568 18478 26580
rect 19518 26568 19524 26580
rect 18472 26540 19524 26568
rect 18472 26528 18478 26540
rect 19518 26528 19524 26540
rect 19576 26528 19582 26580
rect 23290 26528 23296 26580
rect 23348 26568 23354 26580
rect 25869 26571 25927 26577
rect 25869 26568 25881 26571
rect 23348 26540 25881 26568
rect 23348 26528 23354 26540
rect 25869 26537 25881 26540
rect 25915 26537 25927 26571
rect 25869 26531 25927 26537
rect 34885 26571 34943 26577
rect 34885 26537 34897 26571
rect 34931 26568 34943 26571
rect 38010 26568 38016 26580
rect 34931 26540 38016 26568
rect 34931 26537 34943 26540
rect 34885 26531 34943 26537
rect 38010 26528 38016 26540
rect 38068 26528 38074 26580
rect 3329 26503 3387 26509
rect 3329 26469 3341 26503
rect 3375 26500 3387 26503
rect 3602 26500 3608 26512
rect 3375 26472 3608 26500
rect 3375 26469 3387 26472
rect 3329 26463 3387 26469
rect 3602 26460 3608 26472
rect 3660 26460 3666 26512
rect 6273 26503 6331 26509
rect 6273 26469 6285 26503
rect 6319 26500 6331 26503
rect 8573 26503 8631 26509
rect 6319 26472 6960 26500
rect 6319 26469 6331 26472
rect 6273 26463 6331 26469
rect 3970 26432 3976 26444
rect 1596 26404 3976 26432
rect 1596 26376 1624 26404
rect 3970 26392 3976 26404
rect 4028 26392 4034 26444
rect 4249 26435 4307 26441
rect 4249 26401 4261 26435
rect 4295 26432 4307 26435
rect 5810 26432 5816 26444
rect 4295 26404 5816 26432
rect 4295 26401 4307 26404
rect 4249 26395 4307 26401
rect 5810 26392 5816 26404
rect 5868 26392 5874 26444
rect 6822 26432 6828 26444
rect 6783 26404 6828 26432
rect 6822 26392 6828 26404
rect 6880 26392 6886 26444
rect 6932 26432 6960 26472
rect 8573 26469 8585 26503
rect 8619 26500 8631 26503
rect 9398 26500 9404 26512
rect 8619 26472 9404 26500
rect 8619 26469 8631 26472
rect 8573 26463 8631 26469
rect 9398 26460 9404 26472
rect 9456 26460 9462 26512
rect 9582 26460 9588 26512
rect 9640 26500 9646 26512
rect 11330 26500 11336 26512
rect 9640 26472 11336 26500
rect 9640 26460 9646 26472
rect 11330 26460 11336 26472
rect 11388 26500 11394 26512
rect 12250 26500 12256 26512
rect 11388 26472 12256 26500
rect 11388 26460 11394 26472
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 12897 26503 12955 26509
rect 12897 26469 12909 26503
rect 12943 26500 12955 26503
rect 16758 26500 16764 26512
rect 12943 26472 14780 26500
rect 12943 26469 12955 26472
rect 12897 26463 12955 26469
rect 9493 26435 9551 26441
rect 9493 26432 9505 26435
rect 6932 26404 9505 26432
rect 9493 26401 9505 26404
rect 9539 26401 9551 26435
rect 9493 26395 9551 26401
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26432 10195 26435
rect 14366 26432 14372 26444
rect 10183 26404 14372 26432
rect 10183 26401 10195 26404
rect 10137 26395 10195 26401
rect 14366 26392 14372 26404
rect 14424 26392 14430 26444
rect 14642 26432 14648 26444
rect 14603 26404 14648 26432
rect 14642 26392 14648 26404
rect 14700 26392 14706 26444
rect 14752 26432 14780 26472
rect 15396 26472 16436 26500
rect 16719 26472 16764 26500
rect 15396 26432 15424 26472
rect 14752 26404 15424 26432
rect 16408 26432 16436 26472
rect 16758 26460 16764 26472
rect 16816 26460 16822 26512
rect 17497 26503 17555 26509
rect 17497 26469 17509 26503
rect 17543 26469 17555 26503
rect 17497 26463 17555 26469
rect 18141 26503 18199 26509
rect 18141 26469 18153 26503
rect 18187 26500 18199 26503
rect 18690 26500 18696 26512
rect 18187 26472 18696 26500
rect 18187 26469 18199 26472
rect 18141 26463 18199 26469
rect 16470 26435 16528 26441
rect 16470 26432 16482 26435
rect 16408 26404 16482 26432
rect 16470 26401 16482 26404
rect 16516 26401 16528 26435
rect 17512 26432 17540 26463
rect 18690 26460 18696 26472
rect 18748 26460 18754 26512
rect 21358 26460 21364 26512
rect 21416 26500 21422 26512
rect 26326 26500 26332 26512
rect 21416 26472 22600 26500
rect 21416 26460 21422 26472
rect 17512 26404 22140 26432
rect 16470 26395 16528 26401
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 6178 26364 6184 26376
rect 6139 26336 6184 26364
rect 6178 26324 6184 26336
rect 6236 26324 6242 26376
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 2866 26256 2872 26308
rect 2924 26256 2930 26308
rect 3878 26256 3884 26308
rect 3936 26296 3942 26308
rect 3936 26268 4200 26296
rect 3936 26256 3942 26268
rect 4172 26228 4200 26268
rect 4356 26268 4738 26296
rect 4356 26228 4384 26268
rect 5626 26256 5632 26308
rect 5684 26296 5690 26308
rect 5684 26268 7590 26296
rect 8404 26268 9444 26296
rect 5684 26256 5690 26268
rect 4172 26200 4384 26228
rect 4522 26188 4528 26240
rect 4580 26228 4586 26240
rect 7098 26228 7104 26240
rect 4580 26200 7104 26228
rect 4580 26188 4586 26200
rect 7098 26188 7104 26200
rect 7156 26188 7162 26240
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 8404 26228 8432 26268
rect 7800 26200 8432 26228
rect 9416 26228 9444 26268
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 9585 26299 9643 26305
rect 9585 26296 9597 26299
rect 9548 26268 9597 26296
rect 9548 26256 9554 26268
rect 9585 26265 9597 26268
rect 9631 26265 9643 26299
rect 10980 26296 11008 26327
rect 11238 26324 11244 26376
rect 11296 26364 11302 26376
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 11296 26336 11805 26364
rect 11296 26324 11302 26336
rect 11793 26333 11805 26336
rect 11839 26333 11851 26367
rect 11793 26327 11851 26333
rect 12066 26324 12072 26376
rect 12124 26364 12130 26376
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 12124 26336 12265 26364
rect 12124 26324 12130 26336
rect 12253 26333 12265 26336
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26364 13139 26367
rect 13170 26364 13176 26376
rect 13127 26336 13176 26364
rect 13127 26333 13139 26336
rect 13081 26327 13139 26333
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 13722 26364 13728 26376
rect 13683 26336 13728 26364
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 14274 26324 14280 26376
rect 14332 26364 14338 26376
rect 14461 26367 14519 26373
rect 14461 26364 14473 26367
rect 14332 26336 14473 26364
rect 14332 26324 14338 26336
rect 14461 26333 14473 26336
rect 14507 26333 14519 26367
rect 14461 26327 14519 26333
rect 15562 26324 15568 26376
rect 15620 26364 15626 26376
rect 15657 26367 15715 26373
rect 15657 26364 15669 26367
rect 15620 26336 15669 26364
rect 15620 26324 15626 26336
rect 15657 26333 15669 26336
rect 15703 26364 15715 26367
rect 16206 26364 16212 26376
rect 15703 26336 16212 26364
rect 15703 26333 15715 26336
rect 15657 26327 15715 26333
rect 16206 26324 16212 26336
rect 16264 26324 16270 26376
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26364 16359 26367
rect 16408 26364 16528 26366
rect 16666 26364 16672 26376
rect 16347 26338 16672 26364
rect 16347 26336 16436 26338
rect 16500 26336 16672 26338
rect 16347 26333 16359 26336
rect 16301 26327 16359 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17310 26324 17316 26376
rect 17368 26364 17374 26376
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 17368 26336 17693 26364
rect 17368 26324 17374 26336
rect 17681 26333 17693 26336
rect 17727 26364 17739 26367
rect 18046 26364 18052 26376
rect 17727 26336 18052 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 18322 26364 18328 26376
rect 18283 26336 18328 26364
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 22112 26373 22140 26404
rect 22572 26373 22600 26472
rect 23400 26472 26332 26500
rect 23400 26441 23428 26472
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 23385 26435 23443 26441
rect 23385 26401 23397 26435
rect 23431 26401 23443 26435
rect 23566 26432 23572 26444
rect 23527 26404 23572 26432
rect 23385 26395 23443 26401
rect 23566 26392 23572 26404
rect 23624 26392 23630 26444
rect 23750 26392 23756 26444
rect 23808 26432 23814 26444
rect 23808 26404 24900 26432
rect 23808 26392 23814 26404
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 20404 26336 20821 26364
rect 20404 26324 20410 26336
rect 20809 26333 20821 26336
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22097 26327 22155 26333
rect 22557 26367 22615 26373
rect 22557 26333 22569 26367
rect 22603 26333 22615 26367
rect 22557 26327 22615 26333
rect 23474 26324 23480 26376
rect 23532 26364 23538 26376
rect 24765 26367 24823 26373
rect 24765 26364 24777 26367
rect 23532 26336 24777 26364
rect 23532 26324 23538 26336
rect 24765 26333 24777 26336
rect 24811 26333 24823 26367
rect 24872 26364 24900 26404
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 24872 26336 25421 26364
rect 24765 26327 24823 26333
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26333 26111 26367
rect 26053 26327 26111 26333
rect 9585 26259 9643 26265
rect 9692 26268 11008 26296
rect 11057 26299 11115 26305
rect 9692 26228 9720 26268
rect 11057 26265 11069 26299
rect 11103 26296 11115 26299
rect 15749 26299 15807 26305
rect 11103 26268 14504 26296
rect 11103 26265 11115 26268
rect 11057 26259 11115 26265
rect 14476 26240 14504 26268
rect 15749 26265 15761 26299
rect 15795 26296 15807 26299
rect 19518 26296 19524 26308
rect 15795 26268 19380 26296
rect 19479 26268 19524 26296
rect 15795 26265 15807 26268
rect 15749 26259 15807 26265
rect 9416 26200 9720 26228
rect 12345 26231 12403 26237
rect 7800 26188 7806 26200
rect 12345 26197 12357 26231
rect 12391 26228 12403 26231
rect 13170 26228 13176 26240
rect 12391 26200 13176 26228
rect 12391 26197 12403 26200
rect 12345 26191 12403 26197
rect 13170 26188 13176 26200
rect 13228 26188 13234 26240
rect 13538 26228 13544 26240
rect 13499 26200 13544 26228
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 14458 26188 14464 26240
rect 14516 26188 14522 26240
rect 15654 26188 15660 26240
rect 15712 26228 15718 26240
rect 17310 26228 17316 26240
rect 15712 26200 17316 26228
rect 15712 26188 15718 26200
rect 17310 26188 17316 26200
rect 17368 26188 17374 26240
rect 19352 26228 19380 26268
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 19613 26299 19671 26305
rect 19613 26265 19625 26299
rect 19659 26265 19671 26299
rect 19613 26259 19671 26265
rect 20165 26299 20223 26305
rect 20165 26265 20177 26299
rect 20211 26296 20223 26299
rect 21450 26296 21456 26308
rect 20211 26268 21456 26296
rect 20211 26265 20223 26268
rect 20165 26259 20223 26265
rect 19628 26228 19656 26259
rect 21450 26256 21456 26268
rect 21508 26256 21514 26308
rect 24029 26299 24087 26305
rect 24029 26265 24041 26299
rect 24075 26296 24087 26299
rect 24946 26296 24952 26308
rect 24075 26268 24952 26296
rect 24075 26265 24087 26268
rect 24029 26259 24087 26265
rect 24946 26256 24952 26268
rect 25004 26256 25010 26308
rect 26068 26296 26096 26327
rect 34514 26324 34520 26376
rect 34572 26364 34578 26376
rect 35069 26367 35127 26373
rect 35069 26364 35081 26367
rect 34572 26336 35081 26364
rect 34572 26324 34578 26336
rect 35069 26333 35081 26336
rect 35115 26333 35127 26367
rect 35069 26327 35127 26333
rect 25240 26268 26096 26296
rect 20622 26228 20628 26240
rect 19352 26200 19656 26228
rect 20583 26200 20628 26228
rect 20622 26188 20628 26200
rect 20680 26188 20686 26240
rect 20806 26188 20812 26240
rect 20864 26228 20870 26240
rect 21269 26231 21327 26237
rect 21269 26228 21281 26231
rect 20864 26200 21281 26228
rect 20864 26188 20870 26200
rect 21269 26197 21281 26200
rect 21315 26197 21327 26231
rect 21910 26228 21916 26240
rect 21871 26200 21916 26228
rect 21269 26191 21327 26197
rect 21910 26188 21916 26200
rect 21968 26188 21974 26240
rect 22646 26228 22652 26240
rect 22607 26200 22652 26228
rect 22646 26188 22652 26200
rect 22704 26188 22710 26240
rect 24118 26188 24124 26240
rect 24176 26228 24182 26240
rect 25240 26237 25268 26268
rect 24581 26231 24639 26237
rect 24581 26228 24593 26231
rect 24176 26200 24593 26228
rect 24176 26188 24182 26200
rect 24581 26197 24593 26200
rect 24627 26197 24639 26231
rect 24581 26191 24639 26197
rect 25225 26231 25283 26237
rect 25225 26197 25237 26231
rect 25271 26197 25283 26231
rect 25225 26191 25283 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 4522 26024 4528 26036
rect 4264 25996 4528 26024
rect 4264 25956 4292 25996
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 4706 25984 4712 26036
rect 4764 26024 4770 26036
rect 12158 26024 12164 26036
rect 4764 25996 12164 26024
rect 4764 25984 4770 25996
rect 12158 25984 12164 25996
rect 12216 25984 12222 26036
rect 13173 26027 13231 26033
rect 13173 25993 13185 26027
rect 13219 26024 13231 26027
rect 15194 26024 15200 26036
rect 13219 25996 15200 26024
rect 13219 25993 13231 25996
rect 13173 25987 13231 25993
rect 15194 25984 15200 25996
rect 15252 26024 15258 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15252 25996 15853 26024
rect 15252 25984 15258 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 15841 25987 15899 25993
rect 16945 26027 17003 26033
rect 16945 25993 16957 26027
rect 16991 26024 17003 26027
rect 18322 26024 18328 26036
rect 16991 25996 18328 26024
rect 16991 25993 17003 25996
rect 16945 25987 17003 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 18969 26027 19027 26033
rect 18969 25993 18981 26027
rect 19015 26024 19027 26027
rect 20346 26024 20352 26036
rect 19015 25996 20352 26024
rect 19015 25993 19027 25996
rect 18969 25987 19027 25993
rect 20346 25984 20352 25996
rect 20404 25984 20410 26036
rect 20714 26024 20720 26036
rect 20456 25996 20720 26024
rect 3082 25928 4292 25956
rect 4341 25959 4399 25965
rect 4341 25925 4353 25959
rect 4387 25956 4399 25959
rect 4614 25956 4620 25968
rect 4387 25928 4620 25956
rect 4387 25925 4399 25928
rect 4341 25919 4399 25925
rect 4614 25916 4620 25928
rect 4672 25916 4678 25968
rect 5074 25916 5080 25968
rect 5132 25916 5138 25968
rect 5902 25916 5908 25968
rect 5960 25956 5966 25968
rect 8481 25959 8539 25965
rect 8481 25956 8493 25959
rect 5960 25928 8493 25956
rect 5960 25916 5966 25928
rect 8481 25925 8493 25928
rect 8527 25925 8539 25959
rect 8481 25919 8539 25925
rect 8938 25916 8944 25968
rect 8996 25916 9002 25968
rect 10980 25928 13584 25956
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4065 25891 4123 25897
rect 4065 25888 4077 25891
rect 4028 25860 4077 25888
rect 4028 25848 4034 25860
rect 4065 25857 4077 25860
rect 4111 25857 4123 25891
rect 4065 25851 4123 25857
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 10980 25897 11008 25928
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 6972 25860 8217 25888
rect 6972 25848 6978 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 10965 25891 11023 25897
rect 10965 25857 10977 25891
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 12066 25888 12072 25900
rect 11756 25860 12072 25888
rect 11756 25848 11762 25860
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 12158 25848 12164 25900
rect 12216 25888 12222 25900
rect 12713 25891 12771 25897
rect 12216 25860 12664 25888
rect 12216 25848 12222 25860
rect 1578 25820 1584 25832
rect 1539 25792 1584 25820
rect 1578 25780 1584 25792
rect 1636 25780 1642 25832
rect 1857 25823 1915 25829
rect 1857 25789 1869 25823
rect 1903 25820 1915 25823
rect 3602 25820 3608 25832
rect 1903 25792 3464 25820
rect 3563 25792 3608 25820
rect 1903 25789 1915 25792
rect 1857 25783 1915 25789
rect 3436 25752 3464 25792
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 5810 25820 5816 25832
rect 5771 25792 5816 25820
rect 5810 25780 5816 25792
rect 5868 25780 5874 25832
rect 7098 25820 7104 25832
rect 7059 25792 7104 25820
rect 7098 25780 7104 25792
rect 7156 25780 7162 25832
rect 7285 25823 7343 25829
rect 7285 25789 7297 25823
rect 7331 25820 7343 25823
rect 7466 25820 7472 25832
rect 7331 25792 7472 25820
rect 7331 25789 7343 25792
rect 7285 25783 7343 25789
rect 7466 25780 7472 25792
rect 7524 25780 7530 25832
rect 11057 25823 11115 25829
rect 11057 25820 11069 25823
rect 7668 25792 11069 25820
rect 3436 25724 4108 25752
rect 1486 25644 1492 25696
rect 1544 25684 1550 25696
rect 3970 25684 3976 25696
rect 1544 25656 3976 25684
rect 1544 25644 1550 25656
rect 3970 25644 3976 25656
rect 4028 25644 4034 25696
rect 4080 25684 4108 25724
rect 5442 25712 5448 25764
rect 5500 25752 5506 25764
rect 7668 25752 7696 25792
rect 11057 25789 11069 25792
rect 11103 25789 11115 25823
rect 12529 25823 12587 25829
rect 12529 25820 12541 25823
rect 11057 25783 11115 25789
rect 12406 25792 12541 25820
rect 10778 25752 10784 25764
rect 5500 25724 7696 25752
rect 9876 25724 10784 25752
rect 5500 25712 5506 25724
rect 4706 25684 4712 25696
rect 4080 25656 4712 25684
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 7745 25687 7803 25693
rect 7745 25653 7757 25687
rect 7791 25684 7803 25687
rect 9876 25684 9904 25724
rect 10778 25712 10784 25724
rect 10836 25712 10842 25764
rect 10870 25712 10876 25764
rect 10928 25752 10934 25764
rect 12406 25752 12434 25792
rect 12529 25789 12541 25792
rect 12575 25789 12587 25823
rect 12529 25783 12587 25789
rect 10928 25724 12434 25752
rect 12636 25752 12664 25860
rect 12713 25857 12725 25891
rect 12759 25888 12771 25891
rect 12894 25888 12900 25900
rect 12759 25860 12900 25888
rect 12759 25857 12771 25860
rect 12713 25851 12771 25857
rect 12894 25848 12900 25860
rect 12952 25848 12958 25900
rect 13556 25888 13584 25928
rect 13630 25916 13636 25968
rect 13688 25956 13694 25968
rect 19426 25956 19432 25968
rect 13688 25928 15424 25956
rect 13688 25916 13694 25928
rect 13998 25888 14004 25900
rect 13556 25860 14004 25888
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14553 25891 14611 25897
rect 14148 25860 14193 25888
rect 14148 25848 14154 25860
rect 14553 25857 14565 25891
rect 14599 25888 14611 25891
rect 15286 25888 15292 25900
rect 14599 25860 15292 25888
rect 14599 25857 14611 25860
rect 14553 25851 14611 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15396 25897 15424 25928
rect 17788 25928 19432 25956
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15470 25848 15476 25900
rect 15528 25888 15534 25900
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 15528 25860 17141 25888
rect 15528 25848 15534 25860
rect 17129 25857 17141 25860
rect 17175 25888 17187 25891
rect 17402 25888 17408 25900
rect 17175 25860 17408 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 17586 25848 17592 25900
rect 17644 25888 17650 25900
rect 17788 25897 17816 25928
rect 19426 25916 19432 25928
rect 19484 25916 19490 25968
rect 17773 25891 17831 25897
rect 17773 25888 17785 25891
rect 17644 25860 17785 25888
rect 17644 25848 17650 25860
rect 17773 25857 17785 25860
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 18417 25891 18475 25897
rect 18417 25857 18429 25891
rect 18463 25857 18475 25891
rect 19150 25888 19156 25900
rect 19111 25860 19156 25888
rect 18417 25851 18475 25857
rect 15197 25823 15255 25829
rect 15197 25789 15209 25823
rect 15243 25820 15255 25823
rect 17034 25820 17040 25832
rect 15243 25792 17040 25820
rect 15243 25789 15255 25792
rect 15197 25783 15255 25789
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 18432 25820 18460 25851
rect 19150 25848 19156 25860
rect 19208 25848 19214 25900
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25888 19671 25891
rect 20456 25888 20484 25996
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 24397 26027 24455 26033
rect 24397 26024 24409 26027
rect 22756 25996 24409 26024
rect 20806 25956 20812 25968
rect 20767 25928 20812 25956
rect 20806 25916 20812 25928
rect 20864 25916 20870 25968
rect 20898 25916 20904 25968
rect 20956 25956 20962 25968
rect 21450 25956 21456 25968
rect 20956 25928 21001 25956
rect 21411 25928 21456 25956
rect 20956 25916 20962 25928
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 22756 25965 22784 25996
rect 24397 25993 24409 25996
rect 24443 25993 24455 26027
rect 24397 25987 24455 25993
rect 22741 25959 22799 25965
rect 22741 25925 22753 25959
rect 22787 25925 22799 25959
rect 22741 25919 22799 25925
rect 23106 25916 23112 25968
rect 23164 25956 23170 25968
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 23164 25928 23305 25956
rect 23164 25916 23170 25928
rect 23293 25925 23305 25928
rect 23339 25956 23351 25959
rect 26602 25956 26608 25968
rect 23339 25928 26608 25956
rect 23339 25925 23351 25928
rect 23293 25919 23351 25925
rect 26602 25916 26608 25928
rect 26660 25916 26666 25968
rect 23750 25888 23756 25900
rect 19659 25860 20484 25888
rect 23711 25860 23756 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 23750 25848 23756 25860
rect 23808 25848 23814 25900
rect 24578 25888 24584 25900
rect 24539 25860 24584 25888
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25888 27583 25891
rect 34609 25891 34667 25897
rect 34609 25888 34621 25891
rect 27571 25860 34621 25888
rect 27571 25857 27583 25860
rect 27525 25851 27583 25857
rect 34609 25857 34621 25860
rect 34655 25857 34667 25891
rect 34609 25851 34667 25857
rect 17604 25792 18460 25820
rect 19797 25823 19855 25829
rect 14645 25755 14703 25761
rect 12636 25724 14596 25752
rect 10928 25712 10934 25724
rect 7791 25656 9904 25684
rect 7791 25653 7803 25656
rect 7745 25647 7803 25653
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 10008 25656 10053 25684
rect 10008 25644 10014 25656
rect 11238 25644 11244 25696
rect 11296 25684 11302 25696
rect 11885 25687 11943 25693
rect 11885 25684 11897 25687
rect 11296 25656 11897 25684
rect 11296 25644 11302 25656
rect 11885 25653 11897 25656
rect 11931 25653 11943 25687
rect 11885 25647 11943 25653
rect 12526 25644 12532 25696
rect 12584 25684 12590 25696
rect 13262 25684 13268 25696
rect 12584 25656 13268 25684
rect 12584 25644 12590 25656
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 13909 25687 13967 25693
rect 13909 25653 13921 25687
rect 13955 25684 13967 25687
rect 14090 25684 14096 25696
rect 13955 25656 14096 25684
rect 13955 25653 13967 25656
rect 13909 25647 13967 25653
rect 14090 25644 14096 25656
rect 14148 25644 14154 25696
rect 14568 25684 14596 25724
rect 14645 25721 14657 25755
rect 14691 25752 14703 25755
rect 17218 25752 17224 25764
rect 14691 25724 17224 25752
rect 14691 25721 14703 25724
rect 14645 25715 14703 25721
rect 17218 25712 17224 25724
rect 17276 25712 17282 25764
rect 17604 25761 17632 25792
rect 19797 25789 19809 25823
rect 19843 25820 19855 25823
rect 21910 25820 21916 25832
rect 19843 25792 21916 25820
rect 19843 25789 19855 25792
rect 19797 25783 19855 25789
rect 21910 25780 21916 25792
rect 21968 25780 21974 25832
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 25041 25823 25099 25829
rect 25041 25820 25053 25823
rect 22695 25808 23244 25820
rect 23492 25808 25053 25820
rect 22695 25792 25053 25808
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 23216 25780 23520 25792
rect 25041 25789 25053 25792
rect 25087 25789 25099 25823
rect 25041 25783 25099 25789
rect 17589 25755 17647 25761
rect 17589 25721 17601 25755
rect 17635 25721 17647 25755
rect 19978 25752 19984 25764
rect 19939 25724 19984 25752
rect 17589 25715 17647 25721
rect 19978 25712 19984 25724
rect 20036 25712 20042 25764
rect 21726 25712 21732 25764
rect 21784 25752 21790 25764
rect 23106 25752 23112 25764
rect 21784 25724 23112 25752
rect 21784 25712 21790 25724
rect 23106 25712 23112 25724
rect 23164 25712 23170 25764
rect 27448 25752 27476 25851
rect 23676 25724 27476 25752
rect 16114 25684 16120 25696
rect 14568 25656 16120 25684
rect 16114 25644 16120 25656
rect 16172 25644 16178 25696
rect 18230 25684 18236 25696
rect 18191 25656 18236 25684
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 21450 25644 21456 25696
rect 21508 25684 21514 25696
rect 23676 25684 23704 25724
rect 23842 25684 23848 25696
rect 21508 25656 23704 25684
rect 23803 25656 23848 25684
rect 21508 25644 21514 25656
rect 23842 25644 23848 25656
rect 23900 25644 23906 25696
rect 34425 25687 34483 25693
rect 34425 25653 34437 25687
rect 34471 25684 34483 25687
rect 38010 25684 38016 25696
rect 34471 25656 38016 25684
rect 34471 25653 34483 25656
rect 34425 25647 34483 25653
rect 38010 25644 38016 25656
rect 38068 25644 38074 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1844 25483 1902 25489
rect 1844 25449 1856 25483
rect 1890 25480 1902 25483
rect 3970 25480 3976 25492
rect 1890 25452 3648 25480
rect 3931 25452 3976 25480
rect 1890 25449 1902 25452
rect 1844 25443 1902 25449
rect 3620 25424 3648 25452
rect 3970 25440 3976 25452
rect 4028 25440 4034 25492
rect 5534 25480 5540 25492
rect 5495 25452 5540 25480
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 6825 25483 6883 25489
rect 6825 25449 6837 25483
rect 6871 25480 6883 25483
rect 7190 25480 7196 25492
rect 6871 25452 7196 25480
rect 6871 25449 6883 25452
rect 6825 25443 6883 25449
rect 7190 25440 7196 25452
rect 7248 25440 7254 25492
rect 7466 25480 7472 25492
rect 7427 25452 7472 25480
rect 7466 25440 7472 25452
rect 7524 25440 7530 25492
rect 12345 25483 12403 25489
rect 7576 25452 11284 25480
rect 3602 25372 3608 25424
rect 3660 25412 3666 25424
rect 7576 25412 7604 25452
rect 3660 25384 7604 25412
rect 9309 25415 9367 25421
rect 3660 25372 3666 25384
rect 9309 25381 9321 25415
rect 9355 25381 9367 25415
rect 9309 25375 9367 25381
rect 10137 25415 10195 25421
rect 10137 25381 10149 25415
rect 10183 25412 10195 25415
rect 11146 25412 11152 25424
rect 10183 25384 11152 25412
rect 10183 25381 10195 25384
rect 10137 25375 10195 25381
rect 1578 25344 1584 25356
rect 1491 25316 1584 25344
rect 1578 25304 1584 25316
rect 1636 25344 1642 25356
rect 2498 25344 2504 25356
rect 1636 25316 2504 25344
rect 1636 25304 1642 25316
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 5166 25304 5172 25356
rect 5224 25344 5230 25356
rect 8113 25347 8171 25353
rect 8113 25344 8125 25347
rect 5224 25316 8125 25344
rect 5224 25304 5230 25316
rect 8113 25313 8125 25316
rect 8159 25313 8171 25347
rect 9324 25344 9352 25375
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 11256 25412 11284 25452
rect 12345 25449 12357 25483
rect 12391 25480 12403 25483
rect 16574 25480 16580 25492
rect 12391 25452 16160 25480
rect 16535 25452 16580 25480
rect 12391 25449 12403 25452
rect 12345 25443 12403 25449
rect 11256 25384 16068 25412
rect 13538 25344 13544 25356
rect 9324 25316 10364 25344
rect 8113 25307 8171 25313
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 3970 25208 3976 25220
rect 3082 25180 3976 25208
rect 3970 25168 3976 25180
rect 4028 25168 4034 25220
rect 4172 25208 4200 25239
rect 4338 25236 4344 25288
rect 4396 25276 4402 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4396 25248 4905 25276
rect 4396 25236 4402 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 5718 25276 5724 25288
rect 4893 25239 4951 25245
rect 5000 25248 5580 25276
rect 5679 25248 5724 25276
rect 5000 25208 5028 25248
rect 4172 25180 5028 25208
rect 5552 25208 5580 25248
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5902 25236 5908 25288
rect 5960 25276 5966 25288
rect 6733 25279 6791 25285
rect 6733 25276 6745 25279
rect 5960 25248 6745 25276
rect 5960 25236 5966 25248
rect 6733 25245 6745 25248
rect 6779 25245 6791 25279
rect 7374 25276 7380 25288
rect 7287 25248 7380 25276
rect 6733 25239 6791 25245
rect 7374 25236 7380 25248
rect 7432 25276 7438 25288
rect 8021 25279 8079 25285
rect 7432 25248 7972 25276
rect 7432 25236 7438 25248
rect 6638 25208 6644 25220
rect 5552 25180 6644 25208
rect 6638 25168 6644 25180
rect 6696 25168 6702 25220
rect 2682 25100 2688 25152
rect 2740 25140 2746 25152
rect 3329 25143 3387 25149
rect 3329 25140 3341 25143
rect 2740 25112 3341 25140
rect 2740 25100 2746 25112
rect 3329 25109 3341 25112
rect 3375 25109 3387 25143
rect 4982 25140 4988 25152
rect 4943 25112 4988 25140
rect 3329 25103 3387 25109
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 7944 25140 7972 25248
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8036 25208 8064 25239
rect 9214 25236 9220 25288
rect 9272 25276 9278 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 9272 25248 9505 25276
rect 9272 25236 9278 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 9582 25236 9588 25288
rect 9640 25276 9646 25288
rect 10336 25285 10364 25316
rect 12544 25316 13544 25344
rect 10321 25279 10379 25285
rect 9640 25248 10088 25276
rect 9640 25236 9646 25248
rect 9950 25208 9956 25220
rect 8036 25180 9956 25208
rect 9950 25168 9956 25180
rect 10008 25168 10014 25220
rect 10060 25208 10088 25248
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10321 25239 10379 25245
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11241 25279 11299 25285
rect 11241 25276 11253 25279
rect 11112 25248 11253 25276
rect 11112 25236 11118 25248
rect 11241 25245 11253 25248
rect 11287 25245 11299 25279
rect 11241 25239 11299 25245
rect 11330 25236 11336 25288
rect 11388 25276 11394 25288
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 11388 25248 11713 25276
rect 11388 25236 11394 25248
rect 11701 25245 11713 25248
rect 11747 25276 11759 25279
rect 11790 25276 11796 25288
rect 11747 25248 11796 25276
rect 11747 25245 11759 25248
rect 11701 25239 11759 25245
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 12544 25285 12572 25316
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 14366 25304 14372 25356
rect 14424 25344 14430 25356
rect 14645 25347 14703 25353
rect 14645 25344 14657 25347
rect 14424 25316 14657 25344
rect 14424 25304 14430 25316
rect 14645 25313 14657 25316
rect 14691 25344 14703 25347
rect 15102 25344 15108 25356
rect 14691 25316 15108 25344
rect 14691 25313 14703 25316
rect 14645 25307 14703 25313
rect 15102 25304 15108 25316
rect 15160 25304 15166 25356
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 15930 25276 15936 25288
rect 15891 25248 15936 25276
rect 12529 25239 12587 25245
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 16040 25276 16068 25384
rect 16132 25353 16160 25452
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 17310 25440 17316 25492
rect 17368 25480 17374 25492
rect 17405 25483 17463 25489
rect 17405 25480 17417 25483
rect 17368 25452 17417 25480
rect 17368 25440 17374 25452
rect 17405 25449 17417 25452
rect 17451 25480 17463 25483
rect 17586 25480 17592 25492
rect 17451 25452 17592 25480
rect 17451 25449 17463 25452
rect 17405 25443 17463 25449
rect 17586 25440 17592 25452
rect 17644 25440 17650 25492
rect 18138 25440 18144 25492
rect 18196 25480 18202 25492
rect 18601 25483 18659 25489
rect 18601 25480 18613 25483
rect 18196 25452 18613 25480
rect 18196 25440 18202 25452
rect 18601 25449 18613 25452
rect 18647 25480 18659 25483
rect 18874 25480 18880 25492
rect 18647 25452 18880 25480
rect 18647 25449 18659 25452
rect 18601 25443 18659 25449
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 20901 25483 20959 25489
rect 20901 25449 20913 25483
rect 20947 25480 20959 25483
rect 20990 25480 20996 25492
rect 20947 25452 20996 25480
rect 20947 25449 20959 25452
rect 20901 25443 20959 25449
rect 20990 25440 20996 25452
rect 21048 25440 21054 25492
rect 22281 25483 22339 25489
rect 22281 25449 22293 25483
rect 22327 25480 22339 25483
rect 22738 25480 22744 25492
rect 22327 25452 22744 25480
rect 22327 25449 22339 25452
rect 22281 25443 22339 25449
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 23477 25483 23535 25489
rect 23477 25449 23489 25483
rect 23523 25480 23535 25483
rect 23658 25480 23664 25492
rect 23523 25452 23664 25480
rect 23523 25449 23535 25452
rect 23477 25443 23535 25449
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 23750 25412 23756 25424
rect 16224 25384 23756 25412
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25313 16175 25347
rect 16117 25307 16175 25313
rect 16224 25276 16252 25384
rect 23750 25372 23756 25384
rect 23808 25412 23814 25424
rect 24762 25412 24768 25424
rect 23808 25384 24768 25412
rect 23808 25372 23814 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 17218 25344 17224 25356
rect 17179 25316 17224 25344
rect 17218 25304 17224 25316
rect 17276 25304 17282 25356
rect 17494 25304 17500 25356
rect 17552 25344 17558 25356
rect 18417 25347 18475 25353
rect 18417 25344 18429 25347
rect 17552 25316 18429 25344
rect 17552 25304 17558 25316
rect 18417 25313 18429 25316
rect 18463 25313 18475 25347
rect 20254 25344 20260 25356
rect 20215 25316 20260 25344
rect 18417 25307 18475 25313
rect 20254 25304 20260 25316
rect 20312 25304 20318 25356
rect 20441 25347 20499 25353
rect 20441 25313 20453 25347
rect 20487 25344 20499 25347
rect 20622 25344 20628 25356
rect 20487 25316 20628 25344
rect 20487 25313 20499 25316
rect 20441 25307 20499 25313
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 21821 25347 21879 25353
rect 21821 25313 21833 25347
rect 21867 25344 21879 25347
rect 22646 25344 22652 25356
rect 21867 25316 22652 25344
rect 21867 25313 21879 25316
rect 21821 25307 21879 25313
rect 22646 25304 22652 25316
rect 22704 25304 22710 25356
rect 23017 25347 23075 25353
rect 23017 25313 23029 25347
rect 23063 25344 23075 25347
rect 24118 25344 24124 25356
rect 23063 25316 24124 25344
rect 23063 25313 23075 25316
rect 23017 25307 23075 25313
rect 24118 25304 24124 25316
rect 24176 25304 24182 25356
rect 17034 25276 17040 25288
rect 16040 25248 16252 25276
rect 16947 25248 17040 25276
rect 17034 25236 17040 25248
rect 17092 25276 17098 25288
rect 17862 25276 17868 25288
rect 17092 25248 17868 25276
rect 17092 25236 17098 25248
rect 17862 25236 17868 25248
rect 17920 25236 17926 25288
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25276 18291 25279
rect 19334 25276 19340 25288
rect 18279 25248 19340 25276
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 19334 25236 19340 25248
rect 19392 25236 19398 25288
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 19484 25248 19625 25276
rect 19484 25236 19490 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 21542 25236 21548 25288
rect 21600 25276 21606 25288
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 21600 25248 21649 25276
rect 21600 25236 21606 25248
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 22833 25279 22891 25285
rect 22833 25276 22845 25279
rect 21637 25239 21695 25245
rect 22066 25248 22845 25276
rect 13078 25208 13084 25220
rect 10060 25180 12434 25208
rect 13039 25180 13084 25208
rect 9030 25140 9036 25152
rect 7944 25112 9036 25140
rect 9030 25100 9036 25112
rect 9088 25100 9094 25152
rect 10042 25100 10048 25152
rect 10100 25140 10106 25152
rect 10226 25140 10232 25152
rect 10100 25112 10232 25140
rect 10100 25100 10106 25112
rect 10226 25100 10232 25112
rect 10284 25100 10290 25152
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11606 25140 11612 25152
rect 11103 25112 11612 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 11790 25140 11796 25152
rect 11751 25112 11796 25140
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 12406 25140 12434 25180
rect 13078 25168 13084 25180
rect 13136 25168 13142 25220
rect 13170 25168 13176 25220
rect 13228 25208 13234 25220
rect 13722 25208 13728 25220
rect 13228 25180 13273 25208
rect 13683 25180 13728 25208
rect 13228 25168 13234 25180
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 13998 25168 14004 25220
rect 14056 25208 14062 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 14056 25180 14381 25208
rect 14056 25168 14062 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 14458 25168 14464 25220
rect 14516 25208 14522 25220
rect 14516 25180 14561 25208
rect 14516 25168 14522 25180
rect 14826 25168 14832 25220
rect 14884 25208 14890 25220
rect 18966 25208 18972 25220
rect 14884 25180 18972 25208
rect 14884 25168 14890 25180
rect 18966 25168 18972 25180
rect 19024 25168 19030 25220
rect 21174 25168 21180 25220
rect 21232 25208 21238 25220
rect 22066 25208 22094 25248
rect 22833 25245 22845 25248
rect 22879 25245 22891 25279
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 22833 25239 22891 25245
rect 24578 25236 24584 25248
rect 24636 25276 24642 25288
rect 25866 25276 25872 25288
rect 24636 25248 25872 25276
rect 24636 25236 24642 25248
rect 25866 25236 25872 25248
rect 25924 25236 25930 25288
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 21232 25180 22094 25208
rect 21232 25168 21238 25180
rect 15378 25140 15384 25152
rect 12406 25112 15384 25140
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 20806 25140 20812 25152
rect 19475 25112 20812 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 20806 25100 20812 25112
rect 20864 25100 20870 25152
rect 24670 25140 24676 25152
rect 24631 25112 24676 25140
rect 24670 25100 24676 25112
rect 24728 25100 24734 25152
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 2406 24896 2412 24948
rect 2464 24936 2470 24948
rect 12158 24936 12164 24948
rect 2464 24908 12164 24936
rect 2464 24896 2470 24908
rect 12158 24896 12164 24908
rect 12216 24896 12222 24948
rect 13357 24939 13415 24945
rect 13357 24905 13369 24939
rect 13403 24936 13415 24939
rect 15930 24936 15936 24948
rect 13403 24908 15936 24936
rect 13403 24905 13415 24908
rect 13357 24899 13415 24905
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 3510 24828 3516 24880
rect 3568 24828 3574 24880
rect 5810 24828 5816 24880
rect 5868 24868 5874 24880
rect 12250 24868 12256 24880
rect 5868 24840 12256 24868
rect 5868 24828 5874 24840
rect 12250 24828 12256 24840
rect 12308 24828 12314 24880
rect 13078 24828 13084 24880
rect 13136 24868 13142 24880
rect 14826 24868 14832 24880
rect 13136 24840 14832 24868
rect 13136 24828 13142 24840
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 15289 24871 15347 24877
rect 15289 24868 15301 24871
rect 15028 24840 15301 24868
rect 1762 24800 1768 24812
rect 1723 24772 1768 24800
rect 1762 24760 1768 24772
rect 1820 24760 1826 24812
rect 2498 24800 2504 24812
rect 2459 24772 2504 24800
rect 2498 24760 2504 24772
rect 2556 24760 2562 24812
rect 4062 24760 4068 24812
rect 4120 24760 4126 24812
rect 5074 24800 5080 24812
rect 5035 24772 5080 24800
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5534 24800 5540 24812
rect 5495 24772 5540 24800
rect 5534 24760 5540 24772
rect 5592 24760 5598 24812
rect 6546 24800 6552 24812
rect 6507 24772 6552 24800
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 6638 24760 6644 24812
rect 6696 24800 6702 24812
rect 7653 24803 7711 24809
rect 6696 24772 6741 24800
rect 6696 24760 6702 24772
rect 7653 24769 7665 24803
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24800 8815 24803
rect 9214 24800 9220 24812
rect 8803 24772 9220 24800
rect 8803 24769 8815 24772
rect 8757 24763 8815 24769
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 4080 24732 4108 24760
rect 2823 24704 4108 24732
rect 4249 24735 4307 24741
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 4249 24701 4261 24735
rect 4295 24732 4307 24735
rect 4706 24732 4712 24744
rect 4295 24704 4712 24732
rect 4295 24701 4307 24704
rect 4249 24695 4307 24701
rect 4706 24692 4712 24704
rect 4764 24692 4770 24744
rect 5629 24735 5687 24741
rect 5629 24701 5641 24735
rect 5675 24732 5687 24735
rect 7098 24732 7104 24744
rect 5675 24704 7104 24732
rect 5675 24701 5687 24704
rect 5629 24695 5687 24701
rect 7098 24692 7104 24704
rect 7156 24692 7162 24744
rect 4338 24664 4344 24676
rect 3804 24636 4344 24664
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 3804 24596 3832 24636
rect 4338 24624 4344 24636
rect 4396 24624 4402 24676
rect 4890 24664 4896 24676
rect 4851 24636 4896 24664
rect 4890 24624 4896 24636
rect 4948 24624 4954 24676
rect 7668 24664 7696 24763
rect 9214 24760 9220 24772
rect 9272 24760 9278 24812
rect 9398 24800 9404 24812
rect 9359 24772 9404 24800
rect 9398 24760 9404 24772
rect 9456 24760 9462 24812
rect 9490 24760 9496 24812
rect 9548 24800 9554 24812
rect 9548 24772 9593 24800
rect 9548 24760 9554 24772
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 10192 24772 10517 24800
rect 10192 24760 10198 24772
rect 10505 24769 10517 24772
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 10594 24760 10600 24812
rect 10652 24800 10658 24812
rect 11149 24803 11207 24809
rect 11149 24800 11161 24803
rect 10652 24772 11161 24800
rect 10652 24760 10658 24772
rect 11149 24769 11161 24772
rect 11195 24800 11207 24803
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11195 24772 12081 24800
rect 11195 24769 11207 24772
rect 11149 24763 11207 24769
rect 12069 24769 12081 24772
rect 12115 24769 12127 24803
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12069 24763 12127 24769
rect 12176 24772 12909 24800
rect 12176 24732 12204 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 15028 24800 15056 24840
rect 15289 24837 15301 24840
rect 15335 24837 15347 24871
rect 15289 24831 15347 24837
rect 23293 24871 23351 24877
rect 23293 24837 23305 24871
rect 23339 24868 23351 24871
rect 24670 24868 24676 24880
rect 23339 24840 24676 24868
rect 23339 24837 23351 24840
rect 23293 24831 23351 24837
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 12897 24763 12955 24769
rect 13004 24772 15056 24800
rect 17313 24803 17371 24809
rect 13004 24732 13032 24772
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 18506 24800 18512 24812
rect 17359 24772 18368 24800
rect 18467 24772 18512 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 13998 24732 14004 24744
rect 11256 24720 12204 24732
rect 11072 24704 12204 24720
rect 12636 24704 13032 24732
rect 13959 24704 14004 24732
rect 11072 24692 11284 24704
rect 7668 24636 8984 24664
rect 7742 24596 7748 24608
rect 1627 24568 3832 24596
rect 7703 24568 7748 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 8846 24596 8852 24608
rect 8807 24568 8852 24596
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 8956 24596 8984 24636
rect 9582 24624 9588 24676
rect 9640 24664 9646 24676
rect 10321 24667 10379 24673
rect 10321 24664 10333 24667
rect 9640 24636 10333 24664
rect 9640 24624 9646 24636
rect 10321 24633 10333 24636
rect 10367 24633 10379 24667
rect 10321 24627 10379 24633
rect 10965 24667 11023 24673
rect 10965 24633 10977 24667
rect 11011 24664 11023 24667
rect 11072 24664 11100 24692
rect 11011 24636 11100 24664
rect 12161 24667 12219 24673
rect 11011 24633 11023 24636
rect 10965 24627 11023 24633
rect 12161 24633 12173 24667
rect 12207 24664 12219 24667
rect 12636 24664 12664 24704
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 14182 24732 14188 24744
rect 14143 24704 14188 24732
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 15194 24732 15200 24744
rect 15155 24704 15200 24732
rect 15194 24692 15200 24704
rect 15252 24692 15258 24744
rect 15841 24735 15899 24741
rect 15841 24701 15853 24735
rect 15887 24732 15899 24735
rect 16390 24732 16396 24744
rect 15887 24704 16396 24732
rect 15887 24701 15899 24704
rect 15841 24695 15899 24701
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 17494 24732 17500 24744
rect 17455 24704 17500 24732
rect 17494 24692 17500 24704
rect 17552 24692 17558 24744
rect 18340 24732 18368 24772
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 18690 24800 18696 24812
rect 18651 24772 18696 24800
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 19484 24772 19901 24800
rect 19484 24760 19490 24772
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 20806 24760 20812 24812
rect 20864 24800 20870 24812
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 20864 24772 21189 24800
rect 20864 24760 20870 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 22465 24803 22523 24809
rect 22465 24769 22477 24803
rect 22511 24800 22523 24803
rect 22511 24772 23060 24800
rect 22511 24769 22523 24772
rect 22465 24763 22523 24769
rect 18340 24704 20116 24732
rect 12207 24636 12664 24664
rect 12713 24667 12771 24673
rect 12207 24633 12219 24636
rect 12161 24627 12219 24633
rect 12713 24633 12725 24667
rect 12759 24664 12771 24667
rect 17678 24664 17684 24676
rect 12759 24636 15700 24664
rect 17639 24636 17684 24664
rect 12759 24633 12771 24636
rect 12713 24627 12771 24633
rect 11882 24596 11888 24608
rect 8956 24568 11888 24596
rect 11882 24556 11888 24568
rect 11940 24556 11946 24608
rect 13906 24556 13912 24608
rect 13964 24596 13970 24608
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 13964 24568 14381 24596
rect 13964 24556 13970 24568
rect 14369 24565 14381 24568
rect 14415 24565 14427 24599
rect 15672 24596 15700 24636
rect 17678 24624 17684 24636
rect 17736 24624 17742 24676
rect 18874 24664 18880 24676
rect 18835 24636 18880 24664
rect 18874 24624 18880 24636
rect 18932 24624 18938 24676
rect 20088 24664 20116 24704
rect 20162 24692 20168 24744
rect 20220 24732 20226 24744
rect 20349 24735 20407 24741
rect 20349 24732 20361 24735
rect 20220 24704 20361 24732
rect 20220 24692 20226 24704
rect 20349 24701 20361 24704
rect 20395 24701 20407 24735
rect 20349 24695 20407 24701
rect 21358 24664 21364 24676
rect 20088 24636 21364 24664
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 16022 24596 16028 24608
rect 15672 24568 16028 24596
rect 14369 24559 14427 24565
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 19705 24599 19763 24605
rect 19705 24565 19717 24599
rect 19751 24596 19763 24599
rect 20530 24596 20536 24608
rect 19751 24568 20536 24596
rect 19751 24565 19763 24568
rect 19705 24559 19763 24565
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 20990 24596 20996 24608
rect 20951 24568 20996 24596
rect 20990 24556 20996 24568
rect 21048 24556 21054 24608
rect 22278 24596 22284 24608
rect 22239 24568 22284 24596
rect 22278 24556 22284 24568
rect 22336 24556 22342 24608
rect 23032 24596 23060 24772
rect 24394 24760 24400 24812
rect 24452 24800 24458 24812
rect 24489 24803 24547 24809
rect 24489 24800 24501 24803
rect 24452 24772 24501 24800
rect 24452 24760 24458 24772
rect 24489 24769 24501 24772
rect 24535 24800 24547 24803
rect 24949 24803 25007 24809
rect 24949 24800 24961 24803
rect 24535 24772 24961 24800
rect 24535 24769 24547 24772
rect 24489 24763 24547 24769
rect 24949 24769 24961 24772
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24800 25835 24803
rect 26326 24800 26332 24812
rect 25823 24772 26332 24800
rect 25823 24769 25835 24772
rect 25777 24763 25835 24769
rect 26326 24760 26332 24772
rect 26384 24760 26390 24812
rect 27522 24800 27528 24812
rect 27483 24772 27528 24800
rect 27522 24760 27528 24772
rect 27580 24760 27586 24812
rect 27617 24803 27675 24809
rect 27617 24769 27629 24803
rect 27663 24800 27675 24803
rect 34514 24800 34520 24812
rect 27663 24772 34520 24800
rect 27663 24769 27675 24772
rect 27617 24763 27675 24769
rect 34514 24760 34520 24772
rect 34572 24760 34578 24812
rect 23201 24735 23259 24741
rect 23201 24701 23213 24735
rect 23247 24732 23259 24735
rect 23658 24732 23664 24744
rect 23247 24704 23664 24732
rect 23247 24701 23259 24704
rect 23201 24695 23259 24701
rect 23658 24692 23664 24704
rect 23716 24692 23722 24744
rect 23750 24664 23756 24676
rect 23711 24636 23756 24664
rect 23750 24624 23756 24636
rect 23808 24624 23814 24676
rect 24305 24599 24363 24605
rect 24305 24596 24317 24599
rect 23032 24568 24317 24596
rect 24305 24565 24317 24568
rect 24351 24565 24363 24599
rect 24305 24559 24363 24565
rect 24394 24556 24400 24608
rect 24452 24596 24458 24608
rect 25041 24599 25099 24605
rect 25041 24596 25053 24599
rect 24452 24568 25053 24596
rect 24452 24556 24458 24568
rect 25041 24565 25053 24568
rect 25087 24565 25099 24599
rect 25590 24596 25596 24608
rect 25551 24568 25596 24596
rect 25041 24559 25099 24565
rect 25590 24556 25596 24568
rect 25648 24556 25654 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 2406 24392 2412 24404
rect 2367 24364 2412 24392
rect 2406 24352 2412 24364
rect 2464 24352 2470 24404
rect 3050 24392 3056 24404
rect 3011 24364 3056 24392
rect 3050 24352 3056 24364
rect 3108 24352 3114 24404
rect 4062 24392 4068 24404
rect 4023 24364 4068 24392
rect 4062 24352 4068 24364
rect 4120 24352 4126 24404
rect 5074 24352 5080 24404
rect 5132 24392 5138 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 5132 24364 5733 24392
rect 5132 24352 5138 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 5994 24352 6000 24404
rect 6052 24392 6058 24404
rect 6733 24395 6791 24401
rect 6733 24392 6745 24395
rect 6052 24364 6745 24392
rect 6052 24352 6058 24364
rect 6733 24361 6745 24364
rect 6779 24361 6791 24395
rect 6733 24355 6791 24361
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 9674 24392 9680 24404
rect 8536 24364 9680 24392
rect 8536 24352 8542 24364
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 9950 24392 9956 24404
rect 9911 24364 9956 24392
rect 9950 24352 9956 24364
rect 10008 24392 10014 24404
rect 11333 24395 11391 24401
rect 11333 24392 11345 24395
rect 10008 24364 11345 24392
rect 10008 24352 10014 24364
rect 11333 24361 11345 24364
rect 11379 24361 11391 24395
rect 11333 24355 11391 24361
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 12989 24395 13047 24401
rect 12400 24364 12940 24392
rect 12400 24352 12434 24364
rect 1394 24284 1400 24336
rect 1452 24324 1458 24336
rect 1452 24296 4660 24324
rect 1452 24284 1458 24296
rect 3326 24256 3332 24268
rect 1596 24228 3332 24256
rect 1596 24197 1624 24228
rect 3326 24216 3332 24228
rect 3384 24216 3390 24268
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 1581 24151 1639 24157
rect 2317 24191 2375 24197
rect 2317 24157 2329 24191
rect 2363 24157 2375 24191
rect 2317 24151 2375 24157
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3234 24188 3240 24200
rect 3007 24160 3240 24188
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 2332 24120 2360 24151
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 3694 24148 3700 24200
rect 3752 24188 3758 24200
rect 4632 24197 4660 24296
rect 9398 24284 9404 24336
rect 9456 24324 9462 24336
rect 9456 24296 11376 24324
rect 9456 24284 9462 24296
rect 11348 24268 11376 24296
rect 4798 24216 4804 24268
rect 4856 24256 4862 24268
rect 4856 24228 6960 24256
rect 4856 24216 4862 24228
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 3752 24160 3985 24188
rect 3752 24148 3758 24160
rect 3973 24157 3985 24160
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 5902 24188 5908 24200
rect 5863 24160 5908 24188
rect 4617 24151 4675 24157
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 6932 24197 6960 24228
rect 8846 24216 8852 24268
rect 8904 24256 8910 24268
rect 9769 24259 9827 24265
rect 9769 24256 9781 24259
rect 8904 24228 9781 24256
rect 8904 24216 8910 24228
rect 9769 24225 9781 24228
rect 9815 24225 9827 24259
rect 9769 24219 9827 24225
rect 10686 24216 10692 24268
rect 10744 24256 10750 24268
rect 10744 24228 11100 24256
rect 10744 24216 10750 24228
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24157 6975 24191
rect 7558 24188 7564 24200
rect 7519 24160 7564 24188
rect 6917 24151 6975 24157
rect 7558 24148 7564 24160
rect 7616 24148 7622 24200
rect 9585 24191 9643 24197
rect 9585 24157 9597 24191
rect 9631 24188 9643 24191
rect 10410 24188 10416 24200
rect 9631 24160 10416 24188
rect 9631 24157 9643 24160
rect 9585 24151 9643 24157
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 10965 24191 11023 24197
rect 10965 24157 10977 24191
rect 11011 24157 11023 24191
rect 11072 24188 11100 24228
rect 11146 24216 11152 24268
rect 11204 24256 11210 24268
rect 11204 24228 11249 24256
rect 11204 24216 11210 24228
rect 11330 24216 11336 24268
rect 11388 24216 11394 24268
rect 11698 24216 11704 24268
rect 11756 24256 11762 24268
rect 11974 24256 11980 24268
rect 11756 24228 11980 24256
rect 11756 24216 11762 24228
rect 11974 24216 11980 24228
rect 12032 24216 12038 24268
rect 12406 24256 12434 24352
rect 12084 24228 12434 24256
rect 12084 24188 12112 24228
rect 12250 24188 12256 24200
rect 11072 24160 12112 24188
rect 12211 24160 12256 24188
rect 10965 24151 11023 24157
rect 3712 24120 3740 24148
rect 2332 24092 3740 24120
rect 4709 24123 4767 24129
rect 4709 24089 4721 24123
rect 4755 24120 4767 24123
rect 10042 24120 10048 24132
rect 4755 24092 10048 24120
rect 4755 24089 4767 24092
rect 4709 24083 4767 24089
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 10980 24120 11008 24151
rect 12250 24148 12256 24160
rect 12308 24148 12314 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12912 24197 12940 24364
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 14182 24392 14188 24404
rect 13035 24364 14188 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 14553 24395 14611 24401
rect 14553 24361 14565 24395
rect 14599 24392 14611 24395
rect 17494 24392 17500 24404
rect 14599 24364 17500 24392
rect 14599 24361 14611 24364
rect 14553 24355 14611 24361
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 19702 24392 19708 24404
rect 19352 24364 19708 24392
rect 13354 24284 13360 24336
rect 13412 24324 13418 24336
rect 16298 24324 16304 24336
rect 13412 24296 16304 24324
rect 13412 24284 13418 24296
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 16390 24284 16396 24336
rect 16448 24324 16454 24336
rect 16485 24327 16543 24333
rect 16485 24324 16497 24327
rect 16448 24296 16497 24324
rect 16448 24284 16454 24296
rect 16485 24293 16497 24296
rect 16531 24293 16543 24327
rect 16485 24287 16543 24293
rect 17126 24284 17132 24336
rect 17184 24324 17190 24336
rect 19352 24324 19380 24364
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 23661 24395 23719 24401
rect 23661 24361 23673 24395
rect 23707 24392 23719 24395
rect 23934 24392 23940 24404
rect 23707 24364 23940 24392
rect 23707 24361 23719 24364
rect 23661 24355 23719 24361
rect 23934 24352 23940 24364
rect 23992 24352 23998 24404
rect 24946 24392 24952 24404
rect 24907 24364 24952 24392
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 26326 24392 26332 24404
rect 26287 24364 26332 24392
rect 26326 24352 26332 24364
rect 26384 24352 26390 24404
rect 17184 24296 19380 24324
rect 17184 24284 17190 24296
rect 19426 24284 19432 24336
rect 19484 24324 19490 24336
rect 24302 24324 24308 24336
rect 19484 24296 24308 24324
rect 19484 24284 19490 24296
rect 24302 24284 24308 24296
rect 24360 24324 24366 24336
rect 24360 24296 26556 24324
rect 24360 24284 24366 24296
rect 13446 24216 13452 24268
rect 13504 24216 13510 24268
rect 23201 24259 23259 24265
rect 13740 24228 15240 24256
rect 12897 24191 12955 24197
rect 12400 24160 12848 24188
rect 12400 24148 12406 24160
rect 11974 24120 11980 24132
rect 10980 24092 11980 24120
rect 11974 24080 11980 24092
rect 12032 24080 12038 24132
rect 12066 24080 12072 24132
rect 12124 24120 12130 24132
rect 12268 24120 12296 24148
rect 12124 24092 12296 24120
rect 12820 24120 12848 24160
rect 12897 24157 12909 24191
rect 12943 24157 12955 24191
rect 13464 24188 13492 24216
rect 13740 24197 13768 24228
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 13464 24160 13737 24188
rect 12897 24151 12955 24157
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 15212 24197 15240 24228
rect 15764 24228 21220 24256
rect 14737 24191 14795 24197
rect 14737 24188 14749 24191
rect 14148 24160 14749 24188
rect 14148 24148 14154 24160
rect 14737 24157 14749 24160
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15764 24120 15792 24228
rect 16850 24148 16856 24200
rect 16908 24188 16914 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 16908 24160 17877 24188
rect 16908 24148 16914 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24157 18107 24191
rect 19702 24188 19708 24200
rect 19663 24160 19708 24188
rect 18049 24151 18107 24157
rect 12820 24092 15792 24120
rect 15933 24123 15991 24129
rect 12124 24080 12130 24092
rect 15933 24089 15945 24123
rect 15979 24089 15991 24123
rect 15933 24083 15991 24089
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 7653 24055 7711 24061
rect 7653 24021 7665 24055
rect 7699 24052 7711 24055
rect 11514 24052 11520 24064
rect 7699 24024 11520 24052
rect 7699 24021 7711 24024
rect 7653 24015 7711 24021
rect 11514 24012 11520 24024
rect 11572 24012 11578 24064
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 14182 24052 14188 24064
rect 13587 24024 14188 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 15286 24052 15292 24064
rect 15247 24024 15292 24052
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 15948 24052 15976 24083
rect 16022 24080 16028 24132
rect 16080 24120 16086 24132
rect 16080 24092 16125 24120
rect 16080 24080 16086 24092
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 18064 24120 18092 24151
rect 19702 24148 19708 24160
rect 19760 24148 19766 24200
rect 20530 24188 20536 24200
rect 20491 24160 20536 24188
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 21192 24197 21220 24228
rect 23201 24225 23213 24259
rect 23247 24256 23259 24259
rect 23842 24256 23848 24268
rect 23247 24228 23848 24256
rect 23247 24225 23259 24228
rect 23201 24219 23259 24225
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 24486 24216 24492 24268
rect 24544 24256 24550 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24544 24228 24593 24256
rect 24544 24216 24550 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 24765 24259 24823 24265
rect 24765 24225 24777 24259
rect 24811 24256 24823 24259
rect 25590 24256 25596 24268
rect 24811 24228 25596 24256
rect 24811 24225 24823 24228
rect 24765 24219 24823 24225
rect 25590 24216 25596 24228
rect 25648 24216 25654 24268
rect 21177 24191 21235 24197
rect 21177 24157 21189 24191
rect 21223 24188 21235 24191
rect 21821 24191 21879 24197
rect 21821 24188 21833 24191
rect 21223 24160 21833 24188
rect 21223 24157 21235 24160
rect 21177 24151 21235 24157
rect 21821 24157 21833 24160
rect 21867 24157 21879 24191
rect 21821 24151 21879 24157
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24188 23075 24191
rect 24504 24188 24532 24216
rect 25866 24188 25872 24200
rect 23063 24160 24532 24188
rect 25827 24160 25872 24188
rect 23063 24157 23075 24160
rect 23017 24151 23075 24157
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 26528 24197 26556 24296
rect 26513 24191 26571 24197
rect 26513 24157 26525 24191
rect 26559 24157 26571 24191
rect 26513 24151 26571 24157
rect 26602 24148 26608 24200
rect 26660 24188 26666 24200
rect 28813 24191 28871 24197
rect 28813 24188 28825 24191
rect 26660 24160 28825 24188
rect 26660 24148 26666 24160
rect 28813 24157 28825 24160
rect 28859 24157 28871 24191
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 28813 24151 28871 24157
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 16724 24092 18092 24120
rect 16724 24080 16730 24092
rect 18138 24080 18144 24132
rect 18196 24120 18202 24132
rect 27522 24120 27528 24132
rect 18196 24092 27528 24120
rect 18196 24080 18202 24092
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 16574 24052 16580 24064
rect 15948 24024 16580 24052
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 17221 24055 17279 24061
rect 17221 24021 17233 24055
rect 17267 24052 17279 24055
rect 17770 24052 17776 24064
rect 17267 24024 17776 24052
rect 17267 24021 17279 24024
rect 17221 24015 17279 24021
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 18506 24052 18512 24064
rect 18467 24024 18512 24052
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 19978 24052 19984 24064
rect 19843 24024 19984 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20346 24052 20352 24064
rect 20307 24024 20352 24052
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 20993 24055 21051 24061
rect 20993 24021 21005 24055
rect 21039 24052 21051 24055
rect 21450 24052 21456 24064
rect 21039 24024 21456 24052
rect 21039 24021 21051 24024
rect 20993 24015 21051 24021
rect 21450 24012 21456 24024
rect 21508 24012 21514 24064
rect 21913 24055 21971 24061
rect 21913 24021 21925 24055
rect 21959 24052 21971 24055
rect 22738 24052 22744 24064
rect 21959 24024 22744 24052
rect 21959 24021 21971 24024
rect 21913 24015 21971 24021
rect 22738 24012 22744 24024
rect 22796 24012 22802 24064
rect 25682 24052 25688 24064
rect 25643 24024 25688 24052
rect 25682 24012 25688 24024
rect 25740 24012 25746 24064
rect 28905 24055 28963 24061
rect 28905 24021 28917 24055
rect 28951 24052 28963 24055
rect 30190 24052 30196 24064
rect 28951 24024 30196 24052
rect 28951 24021 28963 24024
rect 28905 24015 28963 24021
rect 30190 24012 30196 24024
rect 30248 24012 30254 24064
rect 38102 24052 38108 24064
rect 38063 24024 38108 24052
rect 38102 24012 38108 24024
rect 38160 24012 38166 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 2130 23808 2136 23860
rect 2188 23848 2194 23860
rect 2317 23851 2375 23857
rect 2317 23848 2329 23851
rect 2188 23820 2329 23848
rect 2188 23808 2194 23820
rect 2317 23817 2329 23820
rect 2363 23817 2375 23851
rect 2317 23811 2375 23817
rect 2961 23851 3019 23857
rect 2961 23817 2973 23851
rect 3007 23848 3019 23851
rect 5626 23848 5632 23860
rect 3007 23820 5632 23848
rect 3007 23817 3019 23820
rect 2961 23811 3019 23817
rect 5626 23808 5632 23820
rect 5684 23808 5690 23860
rect 8573 23851 8631 23857
rect 8573 23817 8585 23851
rect 8619 23848 8631 23851
rect 8619 23820 11836 23848
rect 8619 23817 8631 23820
rect 8573 23811 8631 23817
rect 3602 23780 3608 23792
rect 3563 23752 3608 23780
rect 3602 23740 3608 23752
rect 3660 23740 3666 23792
rect 8021 23783 8079 23789
rect 8021 23749 8033 23783
rect 8067 23780 8079 23783
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 8067 23752 9413 23780
rect 8067 23749 8079 23752
rect 8021 23743 8079 23749
rect 9401 23749 9413 23752
rect 9447 23749 9459 23783
rect 9401 23743 9459 23749
rect 9953 23783 10011 23789
rect 9953 23749 9965 23783
rect 9999 23780 10011 23783
rect 9999 23752 11560 23780
rect 9999 23749 10011 23752
rect 9953 23743 10011 23749
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23712 1639 23715
rect 1946 23712 1952 23724
rect 1627 23684 1952 23712
rect 1627 23681 1639 23684
rect 1581 23675 1639 23681
rect 1946 23672 1952 23684
rect 2004 23712 2010 23724
rect 2225 23715 2283 23721
rect 2225 23712 2237 23715
rect 2004 23684 2237 23712
rect 2004 23672 2010 23684
rect 2225 23681 2237 23684
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2240 23644 2268 23675
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 2869 23715 2927 23721
rect 2869 23712 2881 23715
rect 2832 23684 2881 23712
rect 2832 23672 2838 23684
rect 2869 23681 2881 23684
rect 2915 23681 2927 23715
rect 2869 23675 2927 23681
rect 3513 23715 3571 23721
rect 3513 23681 3525 23715
rect 3559 23681 3571 23715
rect 6730 23712 6736 23724
rect 6691 23684 6736 23712
rect 3513 23675 3571 23681
rect 3528 23644 3556 23675
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 7006 23672 7012 23724
rect 7064 23712 7070 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7064 23684 7941 23712
rect 7064 23672 7070 23684
rect 7929 23681 7941 23684
rect 7975 23712 7987 23715
rect 8570 23712 8576 23724
rect 7975 23684 8576 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 8570 23672 8576 23684
rect 8628 23672 8634 23724
rect 8754 23712 8760 23724
rect 8715 23684 8760 23712
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 11146 23712 11152 23724
rect 11059 23684 11152 23712
rect 11146 23672 11152 23684
rect 11204 23712 11210 23724
rect 11330 23712 11336 23724
rect 11204 23684 11336 23712
rect 11204 23672 11210 23684
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 2240 23616 3556 23644
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 9309 23647 9367 23653
rect 9309 23644 9321 23647
rect 6871 23616 9321 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 9309 23613 9321 23616
rect 9355 23613 9367 23647
rect 11532 23644 11560 23752
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 11808 23712 11836 23820
rect 11974 23808 11980 23860
rect 12032 23848 12038 23860
rect 13814 23848 13820 23860
rect 12032 23820 13820 23848
rect 12032 23808 12038 23820
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 15286 23808 15292 23860
rect 15344 23848 15350 23860
rect 18046 23848 18052 23860
rect 15344 23820 18052 23848
rect 15344 23808 15350 23820
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18417 23851 18475 23857
rect 18417 23817 18429 23851
rect 18463 23848 18475 23851
rect 18506 23848 18512 23860
rect 18463 23820 18512 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 20809 23851 20867 23857
rect 20809 23817 20821 23851
rect 20855 23848 20867 23851
rect 21082 23848 21088 23860
rect 20855 23820 21088 23848
rect 20855 23817 20867 23820
rect 20809 23811 20867 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 24394 23848 24400 23860
rect 22296 23820 24400 23848
rect 12342 23740 12348 23792
rect 12400 23780 12406 23792
rect 14829 23783 14887 23789
rect 14829 23780 14841 23783
rect 12400 23752 14841 23780
rect 12400 23740 12406 23752
rect 14829 23749 14841 23752
rect 14875 23749 14887 23783
rect 14829 23743 14887 23749
rect 15010 23740 15016 23792
rect 15068 23780 15074 23792
rect 20438 23780 20444 23792
rect 15068 23752 20444 23780
rect 15068 23740 15074 23752
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 22296 23789 22324 23820
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 22281 23783 22339 23789
rect 22281 23749 22293 23783
rect 22327 23749 22339 23783
rect 22830 23780 22836 23792
rect 22791 23752 22836 23780
rect 22281 23743 22339 23749
rect 22830 23740 22836 23752
rect 22888 23740 22894 23792
rect 25041 23783 25099 23789
rect 25041 23780 25053 23783
rect 23308 23752 25053 23780
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11808 23684 11897 23712
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 11974 23672 11980 23724
rect 12032 23712 12038 23724
rect 13354 23712 13360 23724
rect 12032 23684 13360 23712
rect 12032 23672 12038 23684
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 13538 23712 13544 23724
rect 13499 23684 13544 23712
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 14182 23712 14188 23724
rect 14143 23684 14188 23712
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17313 23715 17371 23721
rect 17313 23712 17325 23715
rect 17184 23684 17325 23712
rect 17184 23672 17190 23684
rect 17313 23681 17325 23684
rect 17359 23681 17371 23715
rect 17770 23712 17776 23724
rect 17731 23684 17776 23712
rect 17313 23675 17371 23681
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 17957 23715 18015 23721
rect 17957 23681 17969 23715
rect 18003 23712 18015 23715
rect 18230 23712 18236 23724
rect 18003 23684 18236 23712
rect 18003 23681 18015 23684
rect 17957 23675 18015 23681
rect 18230 23672 18236 23684
rect 18288 23672 18294 23724
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18340 23684 19073 23712
rect 12710 23644 12716 23656
rect 9309 23607 9367 23613
rect 9646 23616 11376 23644
rect 11532 23616 12716 23644
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23576 1731 23579
rect 8294 23576 8300 23588
rect 1719 23548 8300 23576
rect 1719 23545 1731 23548
rect 1673 23539 1731 23545
rect 8294 23536 8300 23548
rect 8352 23536 8358 23588
rect 8754 23536 8760 23588
rect 8812 23576 8818 23588
rect 9646 23576 9674 23616
rect 8812 23548 9674 23576
rect 8812 23536 8818 23548
rect 11348 23520 11376 23616
rect 12710 23604 12716 23616
rect 12768 23644 12774 23656
rect 13262 23644 13268 23656
rect 12768 23616 13268 23644
rect 12768 23604 12774 23616
rect 13262 23604 13268 23616
rect 13320 23604 13326 23656
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23644 14795 23647
rect 15010 23644 15016 23656
rect 14783 23616 15016 23644
rect 14783 23613 14795 23616
rect 14737 23607 14795 23613
rect 15010 23604 15016 23616
rect 15068 23604 15074 23656
rect 15286 23644 15292 23656
rect 15247 23616 15292 23644
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 18340 23644 18368 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 20990 23712 20996 23724
rect 20395 23684 20996 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 21450 23712 21456 23724
rect 21411 23684 21456 23712
rect 21450 23672 21456 23684
rect 21508 23672 21514 23724
rect 23308 23721 23336 23752
rect 25041 23749 25053 23752
rect 25087 23749 25099 23783
rect 25041 23743 25099 23749
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23681 23351 23715
rect 23934 23712 23940 23724
rect 23895 23684 23940 23712
rect 23293 23675 23351 23681
rect 23934 23672 23940 23684
rect 23992 23672 23998 23724
rect 24578 23712 24584 23724
rect 24539 23684 24584 23712
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 16632 23616 18368 23644
rect 18877 23647 18935 23653
rect 16632 23604 16638 23616
rect 18877 23613 18889 23647
rect 18923 23613 18935 23647
rect 18877 23607 18935 23613
rect 20165 23647 20223 23653
rect 20165 23613 20177 23647
rect 20211 23644 20223 23647
rect 20254 23644 20260 23656
rect 20211 23616 20260 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 11572 23548 12173 23576
rect 11572 23536 11578 23548
rect 12161 23545 12173 23548
rect 12207 23545 12219 23579
rect 15470 23576 15476 23588
rect 12161 23539 12219 23545
rect 12268 23548 15476 23576
rect 8662 23468 8668 23520
rect 8720 23508 8726 23520
rect 10965 23511 11023 23517
rect 10965 23508 10977 23511
rect 8720 23480 10977 23508
rect 8720 23468 8726 23480
rect 10965 23477 10977 23480
rect 11011 23477 11023 23511
rect 10965 23471 11023 23477
rect 11330 23468 11336 23520
rect 11388 23508 11394 23520
rect 12268 23508 12296 23548
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 17218 23536 17224 23588
rect 17276 23576 17282 23588
rect 18892 23576 18920 23607
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 22189 23647 22247 23653
rect 22189 23613 22201 23647
rect 22235 23644 22247 23647
rect 22370 23644 22376 23656
rect 22235 23616 22376 23644
rect 22235 23613 22247 23616
rect 22189 23607 22247 23613
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23523 23616 24440 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 24412 23585 24440 23616
rect 24397 23579 24455 23585
rect 17276 23548 18000 23576
rect 18892 23548 22094 23576
rect 17276 23536 17282 23548
rect 13354 23508 13360 23520
rect 11388 23480 12296 23508
rect 13315 23480 13360 23508
rect 11388 23468 11394 23480
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 14001 23511 14059 23517
rect 14001 23477 14013 23511
rect 14047 23508 14059 23511
rect 17034 23508 17040 23520
rect 14047 23480 17040 23508
rect 14047 23477 14059 23480
rect 14001 23471 14059 23477
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 17129 23511 17187 23517
rect 17129 23477 17141 23511
rect 17175 23508 17187 23511
rect 17862 23508 17868 23520
rect 17175 23480 17868 23508
rect 17175 23477 17187 23480
rect 17129 23471 17187 23477
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 17972 23508 18000 23548
rect 19245 23511 19303 23517
rect 19245 23508 19257 23511
rect 17972 23480 19257 23508
rect 19245 23477 19257 23480
rect 19291 23477 19303 23511
rect 19245 23471 19303 23477
rect 20898 23468 20904 23520
rect 20956 23508 20962 23520
rect 21269 23511 21327 23517
rect 21269 23508 21281 23511
rect 20956 23480 21281 23508
rect 20956 23468 20962 23480
rect 21269 23477 21281 23480
rect 21315 23477 21327 23511
rect 22066 23508 22094 23548
rect 22848 23548 24348 23576
rect 22848 23508 22876 23548
rect 22066 23480 22876 23508
rect 24320 23508 24348 23548
rect 24397 23545 24409 23579
rect 24443 23545 24455 23579
rect 24397 23539 24455 23545
rect 32582 23508 32588 23520
rect 24320 23480 32588 23508
rect 21269 23471 21327 23477
rect 32582 23468 32588 23480
rect 32640 23468 32646 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 2590 23304 2596 23316
rect 1627 23276 2596 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 2961 23307 3019 23313
rect 2961 23273 2973 23307
rect 3007 23304 3019 23307
rect 6086 23304 6092 23316
rect 3007 23276 6092 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 6086 23264 6092 23276
rect 6144 23264 6150 23316
rect 8389 23307 8447 23313
rect 8389 23273 8401 23307
rect 8435 23304 8447 23307
rect 11054 23304 11060 23316
rect 8435 23276 11060 23304
rect 8435 23273 8447 23276
rect 8389 23267 8447 23273
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 11514 23304 11520 23316
rect 11475 23276 11520 23304
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 12158 23264 12164 23316
rect 12216 23304 12222 23316
rect 16301 23307 16359 23313
rect 12216 23276 15608 23304
rect 12216 23264 12222 23276
rect 6362 23196 6368 23248
rect 6420 23236 6426 23248
rect 6420 23208 9812 23236
rect 6420 23196 6426 23208
rect 4982 23128 4988 23180
rect 5040 23168 5046 23180
rect 9401 23171 9459 23177
rect 9401 23168 9413 23171
rect 5040 23140 9413 23168
rect 5040 23128 5046 23140
rect 9401 23137 9413 23140
rect 9447 23137 9459 23171
rect 9401 23131 9459 23137
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 9585 23171 9643 23177
rect 9585 23168 9597 23171
rect 9548 23140 9597 23168
rect 9548 23128 9554 23140
rect 9585 23137 9597 23140
rect 9631 23137 9643 23171
rect 9585 23131 9643 23137
rect 1670 23060 1676 23112
rect 1728 23100 1734 23112
rect 1765 23103 1823 23109
rect 1765 23100 1777 23103
rect 1728 23072 1777 23100
rect 1728 23060 1734 23072
rect 1765 23069 1777 23072
rect 1811 23069 1823 23103
rect 1765 23063 1823 23069
rect 1946 23060 1952 23112
rect 2004 23100 2010 23112
rect 2225 23103 2283 23109
rect 2225 23100 2237 23103
rect 2004 23072 2237 23100
rect 2004 23060 2010 23072
rect 2225 23069 2237 23072
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 5258 23100 5264 23112
rect 2915 23072 5264 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 7101 23103 7159 23109
rect 7101 23069 7113 23103
rect 7147 23100 7159 23103
rect 8573 23103 8631 23109
rect 8573 23100 8585 23103
rect 7147 23072 8585 23100
rect 7147 23069 7159 23072
rect 7101 23063 7159 23069
rect 8573 23069 8585 23072
rect 8619 23069 8631 23103
rect 9784 23100 9812 23208
rect 9950 23196 9956 23248
rect 10008 23236 10014 23248
rect 11977 23239 12035 23245
rect 11977 23236 11989 23239
rect 10008 23208 11989 23236
rect 10008 23196 10014 23208
rect 11977 23205 11989 23208
rect 12023 23205 12035 23239
rect 11977 23199 12035 23205
rect 13265 23239 13323 23245
rect 13265 23205 13277 23239
rect 13311 23236 13323 23239
rect 14737 23239 14795 23245
rect 14737 23236 14749 23239
rect 13311 23208 14749 23236
rect 13311 23205 13323 23208
rect 13265 23199 13323 23205
rect 14737 23205 14749 23208
rect 14783 23236 14795 23239
rect 14918 23236 14924 23248
rect 14783 23208 14924 23236
rect 14783 23205 14795 23208
rect 14737 23199 14795 23205
rect 14918 23196 14924 23208
rect 14976 23196 14982 23248
rect 9858 23128 9864 23180
rect 9916 23168 9922 23180
rect 10870 23168 10876 23180
rect 9916 23140 10876 23168
rect 9916 23128 9922 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 11848 23140 12817 23168
rect 11848 23128 11854 23140
rect 12805 23137 12817 23140
rect 12851 23137 12863 23171
rect 12805 23131 12863 23137
rect 13354 23128 13360 23180
rect 13412 23168 13418 23180
rect 14553 23171 14611 23177
rect 14553 23168 14565 23171
rect 13412 23140 14565 23168
rect 13412 23128 13418 23140
rect 14553 23137 14565 23140
rect 14599 23137 14611 23171
rect 15580 23168 15608 23276
rect 16301 23273 16313 23307
rect 16347 23304 16359 23307
rect 16574 23304 16580 23316
rect 16347 23276 16580 23304
rect 16347 23273 16359 23276
rect 16301 23267 16359 23273
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 24578 23304 24584 23316
rect 24539 23276 24584 23304
rect 24578 23264 24584 23276
rect 24636 23264 24642 23316
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 16666 23236 16672 23248
rect 15703 23208 16672 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 16666 23196 16672 23208
rect 16724 23196 16730 23248
rect 16850 23196 16856 23248
rect 16908 23236 16914 23248
rect 18877 23239 18935 23245
rect 16908 23208 18276 23236
rect 16908 23196 16914 23208
rect 17589 23171 17647 23177
rect 15580 23140 16252 23168
rect 14553 23131 14611 23137
rect 10042 23100 10048 23112
rect 9784 23072 10048 23100
rect 8573 23063 8631 23069
rect 2314 23032 2320 23044
rect 2275 23004 2320 23032
rect 2314 22992 2320 23004
rect 2372 22992 2378 23044
rect 7193 23035 7251 23041
rect 7193 23001 7205 23035
rect 7239 23032 7251 23035
rect 8110 23032 8116 23044
rect 7239 23004 8116 23032
rect 7239 23001 7251 23004
rect 7193 22995 7251 23001
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 8588 23032 8616 23063
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 10686 23100 10692 23112
rect 10244 23072 10692 23100
rect 10244 23032 10272 23072
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 11054 23100 11060 23112
rect 11015 23072 11060 23100
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 12066 23060 12072 23112
rect 12124 23100 12130 23112
rect 12161 23103 12219 23109
rect 12161 23100 12173 23103
rect 12124 23072 12173 23100
rect 12124 23060 12130 23072
rect 12161 23069 12173 23072
rect 12207 23069 12219 23103
rect 12161 23063 12219 23069
rect 12342 23060 12348 23112
rect 12400 23100 12406 23112
rect 12621 23103 12679 23109
rect 12621 23100 12633 23103
rect 12400 23072 12633 23100
rect 12400 23060 12406 23072
rect 12621 23069 12633 23072
rect 12667 23069 12679 23103
rect 14366 23100 14372 23112
rect 14327 23072 14372 23100
rect 12621 23063 12679 23069
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 15562 23100 15568 23112
rect 15523 23072 15568 23100
rect 15562 23060 15568 23072
rect 15620 23060 15626 23112
rect 16224 23109 16252 23140
rect 17589 23137 17601 23171
rect 17635 23168 17647 23171
rect 18138 23168 18144 23180
rect 17635 23140 18144 23168
rect 17635 23137 17647 23140
rect 17589 23131 17647 23137
rect 18138 23128 18144 23140
rect 18196 23128 18202 23180
rect 18248 23177 18276 23208
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 20257 23239 20315 23245
rect 20257 23236 20269 23239
rect 18923 23208 20269 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 20257 23205 20269 23208
rect 20303 23236 20315 23239
rect 20806 23236 20812 23248
rect 20303 23208 20812 23236
rect 20303 23205 20315 23208
rect 20257 23199 20315 23205
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 21174 23196 21180 23248
rect 21232 23196 21238 23248
rect 24946 23236 24952 23248
rect 23400 23208 24952 23236
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23137 18291 23171
rect 18233 23131 18291 23137
rect 20073 23171 20131 23177
rect 20073 23137 20085 23171
rect 20119 23168 20131 23171
rect 20346 23168 20352 23180
rect 20119 23140 20352 23168
rect 20119 23137 20131 23140
rect 20073 23131 20131 23137
rect 20346 23128 20352 23140
rect 20404 23128 20410 23180
rect 20993 23171 21051 23177
rect 20993 23137 21005 23171
rect 21039 23168 21051 23171
rect 21192 23168 21220 23196
rect 22830 23168 22836 23180
rect 21039 23140 21220 23168
rect 22791 23140 22836 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 23400 23177 23428 23208
rect 24946 23196 24952 23208
rect 25004 23196 25010 23248
rect 23385 23171 23443 23177
rect 23385 23137 23397 23171
rect 23431 23137 23443 23171
rect 23842 23168 23848 23180
rect 23803 23140 23848 23168
rect 23385 23131 23443 23137
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 16209 23103 16267 23109
rect 16209 23069 16221 23103
rect 16255 23100 16267 23103
rect 16666 23100 16672 23112
rect 16255 23072 16672 23100
rect 16255 23069 16267 23072
rect 16209 23063 16267 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 18414 23100 18420 23112
rect 18375 23072 18420 23100
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20162 23100 20168 23112
rect 19935 23072 20168 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20162 23060 20168 23072
rect 20220 23060 20226 23112
rect 21174 23100 21180 23112
rect 21135 23072 21180 23100
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 24762 23100 24768 23112
rect 24723 23072 24768 23100
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 8588 23004 10272 23032
rect 10318 22992 10324 23044
rect 10376 23032 10382 23044
rect 13538 23032 13544 23044
rect 10376 23004 13544 23032
rect 10376 22992 10382 23004
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 16942 23032 16948 23044
rect 16903 23004 16948 23032
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 17034 22992 17040 23044
rect 17092 23032 17098 23044
rect 17092 23004 17137 23032
rect 17092 22992 17098 23004
rect 21266 22992 21272 23044
rect 21324 23032 21330 23044
rect 22189 23035 22247 23041
rect 22189 23032 22201 23035
rect 21324 23004 22201 23032
rect 21324 22992 21330 23004
rect 22189 23001 22201 23004
rect 22235 23001 22247 23035
rect 22189 22995 22247 23001
rect 22278 22992 22284 23044
rect 22336 23032 22342 23044
rect 23477 23035 23535 23041
rect 22336 23004 22381 23032
rect 22336 22992 22342 23004
rect 23477 23001 23489 23035
rect 23523 23001 23535 23035
rect 23477 22995 23535 23001
rect 7742 22964 7748 22976
rect 7703 22936 7748 22964
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 10045 22967 10103 22973
rect 10045 22933 10057 22967
rect 10091 22964 10103 22967
rect 12342 22964 12348 22976
rect 10091 22936 12348 22964
rect 10091 22933 10103 22936
rect 10045 22927 10103 22933
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 16850 22964 16856 22976
rect 12860 22936 16856 22964
rect 12860 22924 12866 22936
rect 16850 22924 16856 22936
rect 16908 22924 16914 22976
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 19426 22964 19432 22976
rect 17184 22936 19432 22964
rect 17184 22924 17190 22936
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 21634 22964 21640 22976
rect 21595 22936 21640 22964
rect 21634 22924 21640 22936
rect 21692 22924 21698 22976
rect 22738 22924 22744 22976
rect 22796 22964 22802 22976
rect 23492 22964 23520 22995
rect 22796 22936 23520 22964
rect 22796 22924 22802 22936
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 6730 22760 6736 22772
rect 1627 22732 6736 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 8481 22763 8539 22769
rect 8481 22729 8493 22763
rect 8527 22760 8539 22763
rect 11054 22760 11060 22772
rect 8527 22732 11060 22760
rect 8527 22729 8539 22732
rect 8481 22723 8539 22729
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 11606 22720 11612 22772
rect 11664 22760 11670 22772
rect 13081 22763 13139 22769
rect 11664 22732 11836 22760
rect 11664 22720 11670 22732
rect 7742 22652 7748 22704
rect 7800 22692 7806 22704
rect 7800 22664 11560 22692
rect 7800 22652 7806 22664
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7377 22627 7435 22633
rect 7377 22624 7389 22627
rect 7340 22596 7389 22624
rect 7340 22584 7346 22596
rect 7377 22593 7389 22596
rect 7423 22624 7435 22627
rect 7834 22624 7840 22636
rect 7423 22596 7840 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22624 8447 22627
rect 9677 22627 9735 22633
rect 8435 22596 9628 22624
rect 8435 22593 8447 22596
rect 8389 22587 8447 22593
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22556 9091 22559
rect 9490 22556 9496 22568
rect 9079 22528 9496 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 9600 22488 9628 22596
rect 9677 22593 9689 22627
rect 9723 22624 9735 22627
rect 10042 22624 10048 22636
rect 9723 22596 10048 22624
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 10505 22627 10563 22633
rect 10505 22593 10517 22627
rect 10551 22624 10563 22627
rect 11054 22624 11060 22636
rect 10551 22596 11060 22624
rect 10551 22593 10563 22596
rect 10505 22587 10563 22593
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22624 11207 22627
rect 11330 22624 11336 22636
rect 11195 22596 11336 22624
rect 11195 22593 11207 22596
rect 11149 22587 11207 22593
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 9769 22559 9827 22565
rect 9769 22525 9781 22559
rect 9815 22556 9827 22559
rect 11422 22556 11428 22568
rect 9815 22528 11428 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 11422 22516 11428 22528
rect 11480 22516 11486 22568
rect 11532 22544 11560 22664
rect 11808 22624 11836 22732
rect 13081 22729 13093 22763
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13725 22763 13783 22769
rect 13725 22729 13737 22763
rect 13771 22760 13783 22763
rect 16206 22760 16212 22772
rect 13771 22732 16212 22760
rect 13771 22729 13783 22732
rect 13725 22723 13783 22729
rect 13096 22692 13124 22723
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 17681 22763 17739 22769
rect 17681 22729 17693 22763
rect 17727 22760 17739 22763
rect 21082 22760 21088 22772
rect 17727 22732 18552 22760
rect 17727 22729 17739 22732
rect 17681 22723 17739 22729
rect 13096 22664 14596 22692
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 11808 22596 11897 22624
rect 11885 22593 11897 22596
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 14568 22633 14596 22664
rect 15378 22652 15384 22704
rect 15436 22692 15442 22704
rect 17129 22695 17187 22701
rect 15436 22664 16344 22692
rect 15436 22652 15442 22664
rect 13265 22627 13323 22633
rect 13265 22624 13277 22627
rect 12216 22596 13277 22624
rect 12216 22584 12222 22596
rect 13265 22593 13277 22596
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22593 14611 22627
rect 15470 22624 15476 22636
rect 15431 22596 15476 22624
rect 14553 22587 14611 22593
rect 15470 22584 15476 22596
rect 15528 22584 15534 22636
rect 16316 22633 16344 22664
rect 17129 22661 17141 22695
rect 17175 22692 17187 22695
rect 18414 22692 18420 22704
rect 17175 22664 18420 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 18524 22701 18552 22732
rect 19628 22732 21088 22760
rect 19628 22701 19656 22732
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21174 22720 21180 22772
rect 21232 22760 21238 22772
rect 22097 22763 22155 22769
rect 22097 22760 22109 22763
rect 21232 22732 22109 22760
rect 21232 22720 21238 22732
rect 22097 22729 22109 22732
rect 22143 22729 22155 22763
rect 22097 22723 22155 22729
rect 23937 22763 23995 22769
rect 23937 22729 23949 22763
rect 23983 22760 23995 22763
rect 24026 22760 24032 22772
rect 23983 22732 24032 22760
rect 23983 22729 23995 22732
rect 23937 22723 23995 22729
rect 24026 22720 24032 22732
rect 24084 22720 24090 22772
rect 18509 22695 18567 22701
rect 18509 22661 18521 22695
rect 18555 22661 18567 22695
rect 18509 22655 18567 22661
rect 19613 22695 19671 22701
rect 19613 22661 19625 22695
rect 19659 22661 19671 22695
rect 19613 22655 19671 22661
rect 19705 22695 19763 22701
rect 19705 22661 19717 22695
rect 19751 22692 19763 22695
rect 19978 22692 19984 22704
rect 19751 22664 19984 22692
rect 19751 22661 19763 22664
rect 19705 22655 19763 22661
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 20898 22692 20904 22704
rect 20859 22664 20904 22692
rect 20898 22652 20904 22664
rect 20956 22652 20962 22704
rect 21453 22695 21511 22701
rect 21453 22661 21465 22695
rect 21499 22692 21511 22695
rect 23842 22692 23848 22704
rect 21499 22664 23848 22692
rect 21499 22661 21511 22664
rect 21453 22655 21511 22661
rect 23842 22652 23848 22664
rect 23900 22652 23906 22704
rect 25682 22692 25688 22704
rect 24596 22664 25688 22692
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22593 16359 22627
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 16301 22587 16359 22593
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 17862 22624 17868 22636
rect 17823 22596 17868 22624
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 24596 22633 24624 22664
rect 25682 22652 25688 22664
rect 25740 22652 25746 22704
rect 38102 22692 38108 22704
rect 31726 22664 38108 22692
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 24581 22627 24639 22633
rect 24581 22593 24593 22627
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 11699 22559 11757 22565
rect 11699 22544 11711 22559
rect 11532 22525 11711 22544
rect 11745 22525 11757 22559
rect 11532 22519 11757 22525
rect 11532 22516 11744 22519
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 12345 22559 12403 22565
rect 12345 22556 12357 22559
rect 12308 22528 12357 22556
rect 12308 22516 12314 22528
rect 12345 22525 12357 22528
rect 12391 22525 12403 22559
rect 12345 22519 12403 22525
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 14369 22559 14427 22565
rect 14369 22556 14381 22559
rect 14240 22528 14381 22556
rect 14240 22516 14246 22528
rect 14369 22525 14381 22528
rect 14415 22556 14427 22559
rect 18417 22559 18475 22565
rect 14415 22528 17724 22556
rect 14415 22525 14427 22528
rect 14369 22519 14427 22525
rect 10134 22488 10140 22500
rect 9600 22460 10140 22488
rect 10134 22448 10140 22460
rect 10192 22448 10198 22500
rect 10318 22488 10324 22500
rect 10279 22460 10324 22488
rect 10318 22448 10324 22460
rect 10376 22448 10382 22500
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 14737 22491 14795 22497
rect 14737 22488 14749 22491
rect 10468 22460 14749 22488
rect 10468 22448 10474 22460
rect 14737 22457 14749 22460
rect 14783 22457 14795 22491
rect 14737 22451 14795 22457
rect 15565 22491 15623 22497
rect 15565 22457 15577 22491
rect 15611 22488 15623 22491
rect 16850 22488 16856 22500
rect 15611 22460 16856 22488
rect 15611 22457 15623 22460
rect 15565 22451 15623 22457
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 7193 22423 7251 22429
rect 7193 22420 7205 22423
rect 6052 22392 7205 22420
rect 6052 22380 6058 22392
rect 7193 22389 7205 22392
rect 7239 22389 7251 22423
rect 7193 22383 7251 22389
rect 8570 22380 8576 22432
rect 8628 22420 8634 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 8628 22392 10977 22420
rect 8628 22380 8634 22392
rect 10965 22389 10977 22392
rect 11011 22389 11023 22423
rect 10965 22383 11023 22389
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 12250 22420 12256 22432
rect 11112 22392 12256 22420
rect 11112 22380 11118 22392
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 16117 22423 16175 22429
rect 16117 22389 16129 22423
rect 16163 22420 16175 22423
rect 17310 22420 17316 22432
rect 16163 22392 17316 22420
rect 16163 22389 16175 22392
rect 16117 22383 16175 22389
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 17696 22420 17724 22528
rect 18417 22525 18429 22559
rect 18463 22556 18475 22559
rect 18506 22556 18512 22568
rect 18463 22528 18512 22556
rect 18463 22525 18475 22528
rect 18417 22519 18475 22525
rect 18506 22516 18512 22528
rect 18564 22516 18570 22568
rect 19889 22559 19947 22565
rect 19889 22525 19901 22559
rect 19935 22525 19947 22559
rect 20806 22556 20812 22568
rect 20767 22528 20812 22556
rect 19889 22519 19947 22525
rect 18969 22491 19027 22497
rect 18969 22457 18981 22491
rect 19015 22488 19027 22491
rect 19058 22488 19064 22500
rect 19015 22460 19064 22488
rect 19015 22457 19027 22460
rect 18969 22451 19027 22457
rect 19058 22448 19064 22460
rect 19116 22488 19122 22500
rect 19904 22488 19932 22519
rect 20806 22516 20812 22528
rect 20864 22516 20870 22568
rect 19116 22460 19932 22488
rect 19116 22448 19122 22460
rect 20162 22448 20168 22500
rect 20220 22488 20226 22500
rect 22020 22488 22048 22587
rect 24762 22584 24768 22636
rect 24820 22624 24826 22636
rect 25041 22627 25099 22633
rect 25041 22624 25053 22627
rect 24820 22596 25053 22624
rect 24820 22584 24826 22596
rect 25041 22593 25053 22596
rect 25087 22593 25099 22627
rect 25041 22587 25099 22593
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22624 30343 22627
rect 31726 22624 31754 22664
rect 38102 22652 38108 22664
rect 38160 22652 38166 22704
rect 30331 22596 31754 22624
rect 34977 22627 35035 22633
rect 30331 22593 30343 22596
rect 30285 22587 30343 22593
rect 34977 22593 34989 22627
rect 35023 22593 35035 22627
rect 34977 22587 35035 22593
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22649 22559 22707 22565
rect 22649 22556 22661 22559
rect 22152 22528 22661 22556
rect 22152 22516 22158 22528
rect 22649 22525 22661 22528
rect 22695 22525 22707 22559
rect 22649 22519 22707 22525
rect 23293 22559 23351 22565
rect 23293 22525 23305 22559
rect 23339 22556 23351 22559
rect 23382 22556 23388 22568
rect 23339 22528 23388 22556
rect 23339 22525 23351 22528
rect 23293 22519 23351 22525
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 23477 22559 23535 22565
rect 23477 22525 23489 22559
rect 23523 22556 23535 22559
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 23523 22528 25145 22556
rect 23523 22525 23535 22528
rect 23477 22519 23535 22525
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 30190 22516 30196 22568
rect 30248 22556 30254 22568
rect 34992 22556 35020 22587
rect 30248 22528 35020 22556
rect 30248 22516 30254 22528
rect 24397 22491 24455 22497
rect 24397 22488 24409 22491
rect 20220 22460 22048 22488
rect 23492 22460 24409 22488
rect 20220 22448 20226 22460
rect 23492 22432 23520 22460
rect 24397 22457 24409 22460
rect 24443 22457 24455 22491
rect 24397 22451 24455 22457
rect 20254 22420 20260 22432
rect 17696 22392 20260 22420
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 23474 22380 23480 22432
rect 23532 22380 23538 22432
rect 28258 22380 28264 22432
rect 28316 22420 28322 22432
rect 30377 22423 30435 22429
rect 30377 22420 30389 22423
rect 28316 22392 30389 22420
rect 28316 22380 28322 22392
rect 30377 22389 30389 22392
rect 30423 22389 30435 22423
rect 30377 22383 30435 22389
rect 34793 22423 34851 22429
rect 34793 22389 34805 22423
rect 34839 22420 34851 22423
rect 38010 22420 38016 22432
rect 34839 22392 38016 22420
rect 34839 22389 34851 22392
rect 34793 22383 34851 22389
rect 38010 22380 38016 22392
rect 38068 22380 38074 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3786 22176 3792 22228
rect 3844 22216 3850 22228
rect 11054 22216 11060 22228
rect 3844 22188 11060 22216
rect 3844 22176 3850 22188
rect 11054 22176 11060 22188
rect 11112 22176 11118 22228
rect 11422 22176 11428 22228
rect 11480 22216 11486 22228
rect 12066 22216 12072 22228
rect 11480 22188 12072 22216
rect 11480 22176 11486 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 12250 22176 12256 22228
rect 12308 22216 12314 22228
rect 17034 22216 17040 22228
rect 12308 22188 17040 22216
rect 12308 22176 12314 22188
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18196 22188 18552 22216
rect 18196 22176 18202 22188
rect 7377 22151 7435 22157
rect 7377 22117 7389 22151
rect 7423 22148 7435 22151
rect 7423 22120 9352 22148
rect 7423 22117 7435 22120
rect 7377 22111 7435 22117
rect 8110 22080 8116 22092
rect 8071 22052 8116 22080
rect 8110 22040 8116 22052
rect 8168 22040 8174 22092
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 9214 22080 9220 22092
rect 9171 22052 9220 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 9324 22089 9352 22120
rect 9490 22108 9496 22160
rect 9548 22148 9554 22160
rect 10318 22148 10324 22160
rect 9548 22120 10324 22148
rect 9548 22108 9554 22120
rect 10318 22108 10324 22120
rect 10376 22108 10382 22160
rect 10689 22151 10747 22157
rect 10689 22117 10701 22151
rect 10735 22117 10747 22151
rect 12342 22148 12348 22160
rect 12303 22120 12348 22148
rect 10689 22111 10747 22117
rect 9309 22083 9367 22089
rect 9309 22049 9321 22083
rect 9355 22049 9367 22083
rect 9309 22043 9367 22049
rect 9769 22083 9827 22089
rect 9769 22049 9781 22083
rect 9815 22080 9827 22083
rect 10134 22080 10140 22092
rect 9815 22052 10140 22080
rect 9815 22049 9827 22052
rect 9769 22043 9827 22049
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 10704 22024 10732 22111
rect 12342 22108 12348 22120
rect 12400 22108 12406 22160
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 15160 22120 15332 22148
rect 15160 22108 15166 22120
rect 11054 22040 11060 22092
rect 11112 22080 11118 22092
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11112 22052 11989 22080
rect 11112 22040 11118 22052
rect 11977 22049 11989 22052
rect 12023 22049 12035 22083
rect 11977 22043 12035 22049
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12124 22052 12434 22080
rect 12124 22040 12130 22052
rect 1578 21972 1584 22024
rect 1636 22012 1642 22024
rect 6641 22015 6699 22021
rect 6641 22012 6653 22015
rect 1636 21984 6653 22012
rect 1636 21972 1642 21984
rect 6641 21981 6653 21984
rect 6687 21981 6699 22015
rect 7282 22012 7288 22024
rect 7243 21984 7288 22012
rect 6641 21975 6699 21981
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7926 22012 7932 22024
rect 7887 21984 7932 22012
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 8018 21972 8024 22024
rect 8076 22012 8082 22024
rect 10318 22012 10324 22024
rect 8076 21984 10324 22012
rect 8076 21972 8082 21984
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 10686 21972 10692 22024
rect 10744 21972 10750 22024
rect 10873 22015 10931 22021
rect 10873 21981 10885 22015
rect 10919 21981 10931 22015
rect 10873 21975 10931 21981
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 21981 11391 22015
rect 11333 21975 11391 21981
rect 9398 21904 9404 21956
rect 9456 21944 9462 21956
rect 10502 21944 10508 21956
rect 9456 21916 10508 21944
rect 9456 21904 9462 21916
rect 10502 21904 10508 21916
rect 10560 21904 10566 21956
rect 10888 21944 10916 21975
rect 11348 21944 11376 21975
rect 11606 21972 11612 22024
rect 11664 22012 11670 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11664 21984 12173 22012
rect 11664 21972 11670 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12406 22012 12434 22052
rect 12802 22040 12808 22092
rect 12860 22080 12866 22092
rect 13081 22083 13139 22089
rect 13081 22080 13093 22083
rect 12860 22052 13093 22080
rect 12860 22040 12866 22052
rect 13081 22049 13093 22052
rect 13127 22049 13139 22083
rect 14918 22080 14924 22092
rect 14879 22052 14924 22080
rect 13081 22043 13139 22049
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 15304 22080 15332 22120
rect 17586 22108 17592 22160
rect 17644 22148 17650 22160
rect 18524 22157 18552 22188
rect 18509 22151 18567 22157
rect 17644 22120 18368 22148
rect 17644 22108 17650 22120
rect 16761 22083 16819 22089
rect 16761 22080 16773 22083
rect 15304 22052 16773 22080
rect 16761 22049 16773 22052
rect 16807 22049 16819 22083
rect 16761 22043 16819 22049
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22080 17463 22083
rect 18230 22080 18236 22092
rect 17451 22052 18236 22080
rect 17451 22049 17463 22052
rect 17405 22043 17463 22049
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 18340 22080 18368 22120
rect 18509 22117 18521 22151
rect 18555 22117 18567 22151
rect 19797 22151 19855 22157
rect 19797 22148 19809 22151
rect 18509 22111 18567 22117
rect 19352 22120 19809 22148
rect 19352 22080 19380 22120
rect 19797 22117 19809 22120
rect 19843 22117 19855 22151
rect 19797 22111 19855 22117
rect 20254 22108 20260 22160
rect 20312 22148 20318 22160
rect 20312 22120 23520 22148
rect 20312 22108 20318 22120
rect 18340 22052 19380 22080
rect 19429 22083 19487 22089
rect 19429 22049 19441 22083
rect 19475 22080 19487 22083
rect 20809 22083 20867 22089
rect 19475 22052 20576 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12406 21984 13277 22012
rect 12161 21975 12219 21981
rect 13265 21981 13277 21984
rect 13311 21981 13323 22015
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 13265 21975 13323 21981
rect 15672 21984 16221 22012
rect 10888 21916 11376 21944
rect 6730 21876 6736 21888
rect 6691 21848 6736 21876
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21876 8631 21879
rect 10594 21876 10600 21888
rect 8619 21848 10600 21876
rect 8619 21845 8631 21848
rect 8573 21839 8631 21845
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 11348 21876 11376 21916
rect 11425 21947 11483 21953
rect 11425 21913 11437 21947
rect 11471 21944 11483 21947
rect 15013 21947 15071 21953
rect 15013 21944 15025 21947
rect 11471 21916 15025 21944
rect 11471 21913 11483 21916
rect 11425 21907 11483 21913
rect 15013 21913 15025 21916
rect 15059 21913 15071 21947
rect 15562 21944 15568 21956
rect 15523 21916 15568 21944
rect 15013 21907 15071 21913
rect 15562 21904 15568 21916
rect 15620 21904 15626 21956
rect 12618 21876 12624 21888
rect 11348 21848 12624 21876
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 13354 21836 13360 21888
rect 13412 21876 13418 21888
rect 13725 21879 13783 21885
rect 13725 21876 13737 21879
rect 13412 21848 13737 21876
rect 13412 21836 13418 21848
rect 13725 21845 13737 21848
rect 13771 21845 13783 21879
rect 13725 21839 13783 21845
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15672 21876 15700 21984
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 16850 21904 16856 21956
rect 16908 21944 16914 21956
rect 17954 21944 17960 21956
rect 16908 21916 16953 21944
rect 17915 21916 17960 21944
rect 16908 21904 16914 21916
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 18046 21904 18052 21956
rect 18104 21944 18110 21956
rect 18104 21916 18149 21944
rect 18104 21904 18110 21916
rect 16022 21876 16028 21888
rect 15252 21848 15700 21876
rect 15983 21848 16028 21876
rect 15252 21836 15258 21848
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 19628 21876 19656 21975
rect 20548 21944 20576 22052
rect 20809 22049 20821 22083
rect 20855 22080 20867 22083
rect 21545 22083 21603 22089
rect 21545 22080 21557 22083
rect 20855 22052 21557 22080
rect 20855 22049 20867 22052
rect 20809 22043 20867 22049
rect 21545 22049 21557 22052
rect 21591 22049 21603 22083
rect 23492 22080 23520 22120
rect 31297 22083 31355 22089
rect 31297 22080 31309 22083
rect 23492 22052 31309 22080
rect 21545 22043 21603 22049
rect 31297 22049 31309 22052
rect 31343 22049 31355 22083
rect 31297 22043 31355 22049
rect 20714 22012 20720 22024
rect 20675 21984 20720 22012
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 21358 22012 21364 22024
rect 21319 21984 21364 22012
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 31205 22015 31263 22021
rect 31205 21981 31217 22015
rect 31251 22012 31263 22015
rect 38286 22012 38292 22024
rect 31251 21984 35894 22012
rect 38247 21984 38292 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 21450 21944 21456 21956
rect 20548 21916 21456 21944
rect 21450 21904 21456 21916
rect 21508 21904 21514 21956
rect 22005 21947 22063 21953
rect 22005 21913 22017 21947
rect 22051 21944 22063 21947
rect 22646 21944 22652 21956
rect 22051 21916 22652 21944
rect 22051 21913 22063 21916
rect 22005 21907 22063 21913
rect 22646 21904 22652 21916
rect 22704 21944 22710 21956
rect 23017 21947 23075 21953
rect 23017 21944 23029 21947
rect 22704 21916 23029 21944
rect 22704 21904 22710 21916
rect 23017 21913 23029 21916
rect 23063 21913 23075 21947
rect 23017 21907 23075 21913
rect 23109 21947 23167 21953
rect 23109 21913 23121 21947
rect 23155 21944 23167 21947
rect 23474 21944 23480 21956
rect 23155 21916 23480 21944
rect 23155 21913 23167 21916
rect 23109 21907 23167 21913
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23661 21947 23719 21953
rect 23661 21913 23673 21947
rect 23707 21944 23719 21947
rect 23750 21944 23756 21956
rect 23707 21916 23756 21944
rect 23707 21913 23719 21916
rect 23661 21907 23719 21913
rect 23750 21904 23756 21916
rect 23808 21904 23814 21956
rect 17184 21848 19656 21876
rect 35866 21876 35894 21984
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 35866 21848 38117 21876
rect 17184 21836 17190 21848
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 8389 21675 8447 21681
rect 8389 21641 8401 21675
rect 8435 21672 8447 21675
rect 9398 21672 9404 21684
rect 8435 21644 9404 21672
rect 8435 21641 8447 21644
rect 8389 21635 8447 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 9677 21675 9735 21681
rect 9677 21641 9689 21675
rect 9723 21672 9735 21675
rect 10410 21672 10416 21684
rect 9723 21644 10416 21672
rect 9723 21641 9735 21644
rect 9677 21635 9735 21641
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 10502 21632 10508 21684
rect 10560 21672 10566 21684
rect 11146 21672 11152 21684
rect 10560 21644 11152 21672
rect 10560 21632 10566 21644
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 17126 21672 17132 21684
rect 17087 21644 17132 21672
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18417 21675 18475 21681
rect 18417 21672 18429 21675
rect 18012 21644 18429 21672
rect 18012 21632 18018 21644
rect 18417 21641 18429 21644
rect 18463 21641 18475 21675
rect 18417 21635 18475 21641
rect 21453 21675 21511 21681
rect 21453 21641 21465 21675
rect 21499 21672 21511 21675
rect 21634 21672 21640 21684
rect 21499 21644 21640 21672
rect 21499 21641 21511 21644
rect 21453 21635 21511 21641
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 22646 21672 22652 21684
rect 22607 21644 22652 21672
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 6788 21576 11744 21604
rect 6788 21564 6794 21576
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 8478 21536 8484 21548
rect 7791 21508 8484 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 8478 21496 8484 21508
rect 8536 21496 8542 21548
rect 8573 21539 8631 21545
rect 8573 21505 8585 21539
rect 8619 21536 8631 21539
rect 8662 21536 8668 21548
rect 8619 21508 8668 21536
rect 8619 21505 8631 21508
rect 8573 21499 8631 21505
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 10502 21536 10508 21548
rect 10463 21508 10508 21536
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 10962 21536 10968 21548
rect 10923 21508 10968 21536
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11716 21545 11744 21576
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 14550 21604 14556 21616
rect 12400 21576 13492 21604
rect 14511 21576 14556 21604
rect 12400 21564 12406 21576
rect 11701 21539 11759 21545
rect 11701 21505 11713 21539
rect 11747 21505 11759 21539
rect 11701 21499 11759 21505
rect 12066 21496 12072 21548
rect 12124 21536 12130 21548
rect 13354 21536 13360 21548
rect 12124 21508 13360 21536
rect 12124 21496 12130 21508
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 7098 21468 7104 21480
rect 7059 21440 7104 21468
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 9033 21471 9091 21477
rect 9033 21468 9045 21471
rect 7208 21440 9045 21468
rect 5534 21360 5540 21412
rect 5592 21400 5598 21412
rect 7208 21400 7236 21440
rect 9033 21437 9045 21440
rect 9079 21437 9091 21471
rect 9214 21468 9220 21480
rect 9175 21440 9220 21468
rect 9033 21431 9091 21437
rect 9214 21428 9220 21440
rect 9272 21428 9278 21480
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 9876 21440 11897 21468
rect 5592 21372 7236 21400
rect 7837 21403 7895 21409
rect 5592 21360 5598 21372
rect 7837 21369 7849 21403
rect 7883 21400 7895 21403
rect 9876 21400 9904 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 12989 21471 13047 21477
rect 12989 21437 13001 21471
rect 13035 21437 13047 21471
rect 13170 21468 13176 21480
rect 13131 21440 13176 21468
rect 12989 21431 13047 21437
rect 7883 21372 9904 21400
rect 10321 21403 10379 21409
rect 7883 21369 7895 21372
rect 7837 21363 7895 21369
rect 10321 21369 10333 21403
rect 10367 21400 10379 21403
rect 12894 21400 12900 21412
rect 10367 21372 12900 21400
rect 10367 21369 10379 21372
rect 10321 21363 10379 21369
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 13004 21400 13032 21431
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 13078 21400 13084 21412
rect 13004 21372 13084 21400
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 13372 21409 13400 21496
rect 13464 21468 13492 21576
rect 14550 21564 14556 21576
rect 14608 21564 14614 21616
rect 16482 21564 16488 21616
rect 16540 21604 16546 21616
rect 18690 21604 18696 21616
rect 16540 21576 18696 21604
rect 16540 21564 16546 21576
rect 18690 21564 18696 21576
rect 18748 21604 18754 21616
rect 18748 21576 19104 21604
rect 18748 21564 18754 21576
rect 16022 21496 16028 21548
rect 16080 21536 16086 21548
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 16080 21508 16313 21536
rect 16080 21496 16086 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 17310 21536 17316 21548
rect 17271 21508 17316 21536
rect 16301 21499 16359 21505
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 19076 21545 19104 21576
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 24210 21604 24216 21616
rect 20772 21576 24216 21604
rect 20772 21564 20778 21576
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 19061 21539 19119 21545
rect 17819 21508 18092 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 14461 21471 14519 21477
rect 14461 21468 14473 21471
rect 13464 21440 14473 21468
rect 14461 21437 14473 21440
rect 14507 21437 14519 21471
rect 17788 21468 17816 21499
rect 14461 21431 14519 21437
rect 14568 21440 17816 21468
rect 17957 21471 18015 21477
rect 13357 21403 13415 21409
rect 13357 21369 13369 21403
rect 13403 21369 13415 21403
rect 13357 21363 13415 21369
rect 13446 21360 13452 21412
rect 13504 21400 13510 21412
rect 13630 21400 13636 21412
rect 13504 21372 13636 21400
rect 13504 21360 13510 21372
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 13998 21360 14004 21412
rect 14056 21400 14062 21412
rect 14568 21400 14596 21440
rect 17957 21437 17969 21471
rect 18003 21437 18015 21471
rect 18064 21468 18092 21508
rect 19061 21505 19073 21539
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19484 21508 19533 21536
rect 19484 21496 19490 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22094 21536 22100 21548
rect 22051 21508 22100 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22094 21496 22100 21508
rect 22152 21496 22158 21548
rect 23308 21545 23336 21576
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21505 23995 21539
rect 23937 21499 23995 21505
rect 19242 21468 19248 21480
rect 18064 21440 19248 21468
rect 17957 21431 18015 21437
rect 14056 21372 14596 21400
rect 15013 21403 15071 21409
rect 14056 21360 14062 21372
rect 15013 21369 15025 21403
rect 15059 21369 15071 21403
rect 15013 21363 15071 21369
rect 16117 21403 16175 21409
rect 16117 21369 16129 21403
rect 16163 21400 16175 21403
rect 17972 21400 18000 21431
rect 19242 21428 19248 21440
rect 19300 21428 19306 21480
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 19705 21471 19763 21477
rect 19705 21468 19717 21471
rect 19392 21440 19717 21468
rect 19392 21428 19398 21440
rect 19705 21437 19717 21440
rect 19751 21437 19763 21471
rect 20806 21468 20812 21480
rect 20767 21440 20812 21468
rect 19705 21431 19763 21437
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 20990 21468 20996 21480
rect 20951 21440 20996 21468
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 22189 21471 22247 21477
rect 22189 21437 22201 21471
rect 22235 21468 22247 21471
rect 23952 21468 23980 21499
rect 22235 21440 22968 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 16163 21372 18000 21400
rect 18877 21403 18935 21409
rect 16163 21369 16175 21372
rect 16117 21363 16175 21369
rect 18877 21369 18889 21403
rect 18923 21400 18935 21403
rect 22830 21400 22836 21412
rect 18923 21372 22836 21400
rect 18923 21369 18935 21372
rect 18877 21363 18935 21369
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 9582 21332 9588 21344
rect 8536 21304 9588 21332
rect 8536 21292 8542 21304
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 9674 21292 9680 21344
rect 9732 21332 9738 21344
rect 10962 21332 10968 21344
rect 9732 21304 10968 21332
rect 9732 21292 9738 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 12342 21332 12348 21344
rect 11112 21304 11157 21332
rect 12303 21304 12348 21332
rect 11112 21292 11118 21304
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 15028 21332 15056 21363
rect 22830 21360 22836 21372
rect 22888 21360 22894 21412
rect 15562 21332 15568 21344
rect 15028 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21332 15626 21344
rect 19518 21332 19524 21344
rect 15620 21304 19524 21332
rect 15620 21292 15626 21304
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 20165 21335 20223 21341
rect 20165 21301 20177 21335
rect 20211 21332 20223 21335
rect 20254 21332 20260 21344
rect 20211 21304 20260 21332
rect 20211 21301 20223 21304
rect 20165 21295 20223 21301
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 22940 21332 22968 21440
rect 23124 21440 23980 21468
rect 23124 21409 23152 21440
rect 23109 21403 23167 21409
rect 23109 21369 23121 21403
rect 23155 21369 23167 21403
rect 23109 21363 23167 21369
rect 23753 21335 23811 21341
rect 23753 21332 23765 21335
rect 22940 21304 23765 21332
rect 23753 21301 23765 21304
rect 23799 21301 23811 21335
rect 23753 21295 23811 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 6549 21131 6607 21137
rect 6549 21097 6561 21131
rect 6595 21128 6607 21131
rect 9214 21128 9220 21140
rect 6595 21100 9220 21128
rect 6595 21097 6607 21100
rect 6549 21091 6607 21097
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 10778 21128 10784 21140
rect 10739 21100 10784 21128
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11698 21128 11704 21140
rect 11659 21100 11704 21128
rect 11698 21088 11704 21100
rect 11756 21088 11762 21140
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 16577 21131 16635 21137
rect 16577 21128 16589 21131
rect 12400 21100 16589 21128
rect 12400 21088 12406 21100
rect 16577 21097 16589 21100
rect 16623 21128 16635 21131
rect 16942 21128 16948 21140
rect 16623 21100 16948 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17954 21088 17960 21140
rect 18012 21128 18018 21140
rect 18049 21131 18107 21137
rect 18049 21128 18061 21131
rect 18012 21100 18061 21128
rect 18012 21088 18018 21100
rect 18049 21097 18061 21100
rect 18095 21097 18107 21131
rect 18049 21091 18107 21097
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 22925 21131 22983 21137
rect 22925 21128 22937 21131
rect 21048 21100 22937 21128
rect 21048 21088 21054 21100
rect 22925 21097 22937 21100
rect 22971 21097 22983 21131
rect 22925 21091 22983 21097
rect 23014 21088 23020 21140
rect 23072 21128 23078 21140
rect 23072 21100 23796 21128
rect 23072 21088 23078 21100
rect 8018 21060 8024 21072
rect 7024 21032 8024 21060
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20924 6515 20927
rect 7024 20924 7052 21032
rect 8018 21020 8024 21032
rect 8076 21020 8082 21072
rect 8294 21020 8300 21072
rect 8352 21060 8358 21072
rect 13078 21060 13084 21072
rect 8352 21032 10272 21060
rect 8352 21020 8358 21032
rect 7098 20952 7104 21004
rect 7156 20992 7162 21004
rect 10137 20995 10195 21001
rect 10137 20992 10149 20995
rect 7156 20964 10149 20992
rect 7156 20952 7162 20964
rect 10137 20961 10149 20964
rect 10183 20961 10195 20995
rect 10244 20992 10272 21032
rect 10520 21032 13084 21060
rect 10321 20995 10379 21001
rect 10321 20992 10333 20995
rect 10244 20964 10333 20992
rect 10137 20955 10195 20961
rect 10321 20961 10333 20964
rect 10367 20961 10379 20995
rect 10321 20955 10379 20961
rect 6503 20896 7052 20924
rect 7285 20927 7343 20933
rect 6503 20893 6515 20896
rect 6457 20887 6515 20893
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7374 20924 7380 20936
rect 7331 20896 7380 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7374 20884 7380 20896
rect 7432 20924 7438 20936
rect 7834 20924 7840 20936
rect 7432 20896 7840 20924
rect 7432 20884 7438 20896
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 8570 20924 8576 20936
rect 8531 20896 8576 20924
rect 8570 20884 8576 20896
rect 8628 20884 8634 20936
rect 9674 20924 9680 20936
rect 9635 20896 9680 20924
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 10520 20924 10548 21032
rect 13078 21020 13084 21032
rect 13136 21020 13142 21072
rect 14277 21063 14335 21069
rect 14277 21029 14289 21063
rect 14323 21060 14335 21063
rect 19889 21063 19947 21069
rect 14323 21032 16436 21060
rect 14323 21029 14335 21032
rect 14277 21023 14335 21029
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 13170 20992 13176 21004
rect 11388 20964 13176 20992
rect 11388 20952 11394 20964
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 13446 20992 13452 21004
rect 13407 20964 13452 20992
rect 13446 20952 13452 20964
rect 13504 20992 13510 21004
rect 13722 20992 13728 21004
rect 13504 20964 13728 20992
rect 13504 20952 13510 20964
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 15562 20992 15568 21004
rect 14476 20964 15568 20992
rect 10336 20896 10548 20924
rect 7745 20859 7803 20865
rect 7745 20825 7757 20859
rect 7791 20856 7803 20859
rect 10336 20856 10364 20896
rect 10686 20884 10692 20936
rect 10744 20924 10750 20936
rect 14476 20933 14504 20964
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 16206 20992 16212 21004
rect 16167 20964 16212 20992
rect 16206 20952 16212 20964
rect 16264 20952 16270 21004
rect 16408 21001 16436 21032
rect 19889 21029 19901 21063
rect 19935 21060 19947 21063
rect 19935 21032 23152 21060
rect 19935 21029 19947 21032
rect 19889 21023 19947 21029
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20961 16451 20995
rect 16393 20955 16451 20961
rect 21177 20995 21235 21001
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 21266 20992 21272 21004
rect 21223 20964 21272 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 21634 20952 21640 21004
rect 21692 20992 21698 21004
rect 21821 20995 21879 21001
rect 21821 20992 21833 20995
rect 21692 20964 21833 20992
rect 21692 20952 21698 20964
rect 21821 20961 21833 20964
rect 21867 20961 21879 20995
rect 21821 20955 21879 20961
rect 11885 20927 11943 20933
rect 11885 20924 11897 20927
rect 10744 20896 11897 20924
rect 10744 20884 10750 20896
rect 11885 20893 11897 20896
rect 11931 20893 11943 20927
rect 12529 20927 12587 20933
rect 12529 20924 12541 20927
rect 11885 20887 11943 20893
rect 12406 20896 12541 20924
rect 7791 20828 10364 20856
rect 7791 20825 7803 20828
rect 7745 20819 7803 20825
rect 10502 20816 10508 20868
rect 10560 20856 10566 20868
rect 12406 20856 12434 20896
rect 12529 20893 12541 20896
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 15194 20924 15200 20936
rect 14967 20896 15200 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 13078 20856 13084 20868
rect 10560 20828 12434 20856
rect 13039 20828 13084 20856
rect 10560 20816 10566 20828
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 13173 20859 13231 20865
rect 13173 20825 13185 20859
rect 13219 20825 13231 20859
rect 13173 20819 13231 20825
rect 7101 20791 7159 20797
rect 7101 20757 7113 20791
rect 7147 20788 7159 20791
rect 7650 20788 7656 20800
rect 7147 20760 7656 20788
rect 7147 20757 7159 20760
rect 7101 20751 7159 20757
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 9398 20788 9404 20800
rect 8435 20760 9404 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 10410 20788 10416 20800
rect 9539 20760 10416 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 12158 20748 12164 20800
rect 12216 20788 12222 20800
rect 12345 20791 12403 20797
rect 12345 20788 12357 20791
rect 12216 20760 12357 20788
rect 12216 20748 12222 20760
rect 12345 20757 12357 20760
rect 12391 20757 12403 20791
rect 12345 20751 12403 20757
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 13188 20788 13216 20819
rect 12952 20760 13216 20788
rect 12952 20748 12958 20760
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 14936 20788 14964 20887
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15470 20884 15476 20936
rect 15528 20924 15534 20936
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 15528 20896 15761 20924
rect 15528 20884 15534 20896
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 17678 20924 17684 20936
rect 17639 20896 17684 20924
rect 15749 20887 15807 20893
rect 17678 20884 17684 20896
rect 17736 20884 17742 20936
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 15013 20859 15071 20865
rect 15013 20825 15025 20859
rect 15059 20856 15071 20859
rect 17880 20856 17908 20887
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 20073 20927 20131 20933
rect 20073 20924 20085 20927
rect 19484 20896 20085 20924
rect 19484 20884 19490 20896
rect 20073 20893 20085 20896
rect 20119 20924 20131 20927
rect 20162 20924 20168 20936
rect 20119 20896 20168 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20530 20924 20536 20936
rect 20491 20896 20536 20924
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 22554 20924 22560 20936
rect 22511 20896 22560 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 23124 20933 23152 21032
rect 23768 20933 23796 21100
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 23753 20927 23811 20933
rect 23753 20893 23765 20927
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 25038 20924 25044 20936
rect 24811 20896 25044 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 38010 20924 38016 20936
rect 37971 20896 38016 20924
rect 38010 20884 38016 20896
rect 38068 20884 38074 20936
rect 15059 20828 17908 20856
rect 21913 20859 21971 20865
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 21913 20825 21925 20859
rect 21959 20856 21971 20859
rect 21959 20828 22094 20856
rect 21959 20825 21971 20828
rect 21913 20819 21971 20825
rect 13412 20760 14964 20788
rect 15565 20791 15623 20797
rect 13412 20748 13418 20760
rect 15565 20757 15577 20791
rect 15611 20788 15623 20791
rect 16758 20788 16764 20800
rect 15611 20760 16764 20788
rect 15611 20757 15623 20760
rect 15565 20751 15623 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 20162 20788 20168 20800
rect 19576 20760 20168 20788
rect 19576 20748 19582 20760
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 22066 20788 22094 20828
rect 22572 20828 23612 20856
rect 22572 20788 22600 20828
rect 23584 20797 23612 20828
rect 22066 20760 22600 20788
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20757 23627 20791
rect 23569 20751 23627 20757
rect 24026 20748 24032 20800
rect 24084 20788 24090 20800
rect 24581 20791 24639 20797
rect 24581 20788 24593 20791
rect 24084 20760 24593 20788
rect 24084 20748 24090 20760
rect 24581 20757 24593 20760
rect 24627 20757 24639 20791
rect 38194 20788 38200 20800
rect 38155 20760 38200 20788
rect 24581 20751 24639 20757
rect 38194 20748 38200 20760
rect 38252 20748 38258 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5534 20584 5540 20596
rect 5307 20556 5540 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 8294 20584 8300 20596
rect 7791 20556 8300 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 9033 20587 9091 20593
rect 9033 20553 9045 20587
rect 9079 20584 9091 20587
rect 13078 20584 13084 20596
rect 9079 20556 13084 20584
rect 9079 20553 9091 20556
rect 9033 20547 9091 20553
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 16853 20587 16911 20593
rect 13228 20556 16804 20584
rect 13228 20544 13234 20556
rect 7193 20519 7251 20525
rect 7193 20485 7205 20519
rect 7239 20516 7251 20519
rect 7239 20488 11468 20516
rect 7239 20485 7251 20488
rect 7193 20479 7251 20485
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 5169 20451 5227 20457
rect 5169 20448 5181 20451
rect 1636 20420 5181 20448
rect 1636 20408 1642 20420
rect 5169 20417 5181 20420
rect 5215 20417 5227 20451
rect 5994 20448 6000 20460
rect 5955 20420 6000 20448
rect 5169 20411 5227 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7116 20380 7144 20411
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7708 20420 7941 20448
rect 7708 20408 7714 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 8570 20448 8576 20460
rect 8531 20420 8576 20448
rect 7929 20411 7987 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 9858 20448 9864 20460
rect 9771 20420 9864 20448
rect 9858 20408 9864 20420
rect 9916 20448 9922 20460
rect 10318 20448 10324 20460
rect 9916 20420 10324 20448
rect 9916 20408 9922 20420
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20417 10563 20451
rect 11330 20448 11336 20460
rect 10505 20411 10563 20417
rect 10612 20420 11336 20448
rect 9030 20380 9036 20392
rect 7116 20352 9036 20380
rect 9030 20340 9036 20352
rect 9088 20380 9094 20392
rect 9398 20380 9404 20392
rect 9088 20352 9404 20380
rect 9088 20340 9094 20352
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 10520 20380 10548 20411
rect 9692 20352 10548 20380
rect 9692 20321 9720 20352
rect 9677 20315 9735 20321
rect 9677 20281 9689 20315
rect 9723 20281 9735 20315
rect 10612 20312 10640 20420
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 11440 20380 11468 20488
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 11793 20519 11851 20525
rect 11793 20516 11805 20519
rect 11572 20488 11805 20516
rect 11572 20476 11578 20488
rect 11793 20485 11805 20488
rect 11839 20485 11851 20519
rect 11793 20479 11851 20485
rect 11882 20476 11888 20528
rect 11940 20516 11946 20528
rect 11940 20488 11985 20516
rect 11940 20476 11946 20488
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 16114 20516 16120 20528
rect 13044 20488 16120 20516
rect 13044 20476 13050 20488
rect 16114 20476 16120 20488
rect 16172 20476 16178 20528
rect 16776 20516 16804 20556
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 16899 20556 19012 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 18874 20516 18880 20528
rect 16776 20488 18880 20516
rect 18874 20476 18880 20488
rect 18932 20476 18938 20528
rect 18984 20525 19012 20556
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 20864 20556 22017 20584
rect 20864 20544 20870 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 25038 20584 25044 20596
rect 24999 20556 25044 20584
rect 22005 20547 22063 20553
rect 25038 20544 25044 20556
rect 25096 20544 25102 20596
rect 18969 20519 19027 20525
rect 18969 20485 18981 20519
rect 19015 20485 19027 20519
rect 20346 20516 20352 20528
rect 20307 20488 20352 20516
rect 18969 20479 19027 20485
rect 20346 20476 20352 20488
rect 20404 20476 20410 20528
rect 22830 20516 22836 20528
rect 22791 20488 22836 20516
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 24026 20516 24032 20528
rect 23987 20488 24032 20516
rect 24026 20476 24032 20488
rect 24084 20476 24090 20528
rect 14461 20451 14519 20457
rect 14461 20448 14473 20451
rect 13096 20420 14473 20448
rect 11882 20380 11888 20392
rect 11440 20352 11888 20380
rect 10965 20343 11023 20349
rect 9677 20275 9735 20281
rect 10152 20284 10640 20312
rect 5813 20247 5871 20253
rect 5813 20213 5825 20247
rect 5859 20244 5871 20247
rect 7098 20244 7104 20256
rect 5859 20216 7104 20244
rect 5859 20213 5871 20216
rect 5813 20207 5871 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 8389 20247 8447 20253
rect 8389 20213 8401 20247
rect 8435 20244 8447 20247
rect 10152 20244 10180 20284
rect 8435 20216 10180 20244
rect 10321 20247 10379 20253
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 10321 20213 10333 20247
rect 10367 20244 10379 20247
rect 10870 20244 10876 20256
rect 10367 20216 10876 20244
rect 10367 20213 10379 20216
rect 10321 20207 10379 20213
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 10980 20244 11008 20343
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 13096 20380 13124 20420
rect 14461 20417 14473 20420
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 15470 20408 15476 20460
rect 15528 20448 15534 20460
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15528 20420 15577 20448
rect 15528 20408 15534 20420
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16816 20420 17049 20448
rect 16816 20408 16822 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 18322 20448 18328 20460
rect 18283 20420 18328 20448
rect 17037 20411 17095 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 25225 20451 25283 20457
rect 25225 20448 25237 20451
rect 24636 20420 25237 20448
rect 24636 20408 24642 20420
rect 25225 20417 25237 20420
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 11992 20352 13124 20380
rect 13173 20383 13231 20389
rect 11146 20272 11152 20324
rect 11204 20312 11210 20324
rect 11992 20312 12020 20352
rect 13173 20349 13185 20383
rect 13219 20349 13231 20383
rect 13354 20380 13360 20392
rect 13315 20352 13360 20380
rect 13173 20343 13231 20349
rect 11204 20284 12020 20312
rect 12345 20315 12403 20321
rect 11204 20272 11210 20284
rect 12345 20281 12357 20315
rect 12391 20312 12403 20315
rect 12894 20312 12900 20324
rect 12391 20284 12900 20312
rect 12391 20281 12403 20284
rect 12345 20275 12403 20281
rect 12894 20272 12900 20284
rect 12952 20272 12958 20324
rect 12986 20272 12992 20324
rect 13044 20312 13050 20324
rect 13188 20312 13216 20343
rect 13354 20340 13360 20352
rect 13412 20340 13418 20392
rect 13630 20340 13636 20392
rect 13688 20340 13694 20392
rect 13722 20340 13728 20392
rect 13780 20380 13786 20392
rect 14274 20380 14280 20392
rect 13780 20352 14280 20380
rect 13780 20340 13786 20352
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 15381 20383 15439 20389
rect 15381 20349 15393 20383
rect 15427 20380 15439 20383
rect 17218 20380 17224 20392
rect 15427 20352 17224 20380
rect 15427 20349 15439 20352
rect 15381 20343 15439 20349
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20380 17555 20383
rect 18877 20383 18935 20389
rect 18877 20380 18889 20383
rect 17543 20352 18889 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 18877 20349 18889 20352
rect 18923 20349 18935 20383
rect 20254 20380 20260 20392
rect 20215 20352 20260 20380
rect 18877 20343 18935 20349
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 22738 20380 22744 20392
rect 22699 20352 22744 20380
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 23934 20380 23940 20392
rect 23895 20352 23940 20380
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 13044 20284 13216 20312
rect 13648 20312 13676 20340
rect 17586 20312 17592 20324
rect 13648 20284 17592 20312
rect 13044 20272 13050 20284
rect 17586 20272 17592 20284
rect 17644 20272 17650 20324
rect 18141 20315 18199 20321
rect 18141 20281 18153 20315
rect 18187 20312 18199 20315
rect 19334 20312 19340 20324
rect 18187 20284 19340 20312
rect 18187 20281 18199 20284
rect 18141 20275 18199 20281
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 19429 20315 19487 20321
rect 19429 20281 19441 20315
rect 19475 20281 19487 20315
rect 19429 20275 19487 20281
rect 20809 20315 20867 20321
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 22554 20312 22560 20324
rect 20855 20284 22560 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 13630 20244 13636 20256
rect 10980 20216 13636 20244
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 14642 20244 14648 20256
rect 14603 20216 14648 20244
rect 14642 20204 14648 20216
rect 14700 20204 14706 20256
rect 15746 20244 15752 20256
rect 15707 20216 15752 20244
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19444 20244 19472 20275
rect 22554 20272 22560 20284
rect 22612 20272 22618 20324
rect 23293 20315 23351 20321
rect 23293 20281 23305 20315
rect 23339 20312 23351 20315
rect 24486 20312 24492 20324
rect 23339 20284 24492 20312
rect 23339 20281 23351 20284
rect 23293 20275 23351 20281
rect 24486 20272 24492 20284
rect 24544 20272 24550 20324
rect 26326 20244 26332 20256
rect 18288 20216 26332 20244
rect 18288 20204 18294 20216
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 5905 20043 5963 20049
rect 5905 20009 5917 20043
rect 5951 20040 5963 20043
rect 7926 20040 7932 20052
rect 5951 20012 7932 20040
rect 5951 20009 5963 20012
rect 5905 20003 5963 20009
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 9140 20012 10916 20040
rect 6454 19932 6460 19984
rect 6512 19972 6518 19984
rect 6512 19944 8064 19972
rect 6512 19932 6518 19944
rect 7098 19864 7104 19916
rect 7156 19904 7162 19916
rect 7929 19907 7987 19913
rect 7929 19904 7941 19907
rect 7156 19876 7941 19904
rect 7156 19864 7162 19876
rect 7929 19873 7941 19876
rect 7975 19873 7987 19907
rect 7929 19867 7987 19873
rect 5810 19836 5816 19848
rect 5771 19808 5816 19836
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 7190 19836 7196 19848
rect 6687 19808 7196 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 7190 19796 7196 19808
rect 7248 19796 7254 19848
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8036 19836 8064 19944
rect 9140 19913 9168 20012
rect 10778 19972 10784 19984
rect 10520 19944 10784 19972
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 10318 19904 10324 19916
rect 9272 19876 10324 19904
rect 9272 19864 9278 19876
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 10520 19913 10548 19944
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 10888 19972 10916 20012
rect 10962 20000 10968 20052
rect 11020 20040 11026 20052
rect 13354 20040 13360 20052
rect 11020 20012 13360 20040
rect 11020 20000 11026 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 15289 20043 15347 20049
rect 15289 20040 15301 20043
rect 13872 20012 15301 20040
rect 13872 20000 13878 20012
rect 15289 20009 15301 20012
rect 15335 20009 15347 20043
rect 15289 20003 15347 20009
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17218 20040 17224 20052
rect 16807 20012 17224 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 20346 20040 20352 20052
rect 18831 20012 20352 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20533 20043 20591 20049
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 21266 20040 21272 20052
rect 20579 20012 21272 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21542 20040 21548 20052
rect 21503 20012 21548 20040
rect 21542 20000 21548 20012
rect 21600 20040 21606 20052
rect 22465 20043 22523 20049
rect 22465 20040 22477 20043
rect 21600 20012 22477 20040
rect 21600 20000 21606 20012
rect 22465 20009 22477 20012
rect 22511 20009 22523 20043
rect 22465 20003 22523 20009
rect 22830 20000 22836 20052
rect 22888 20040 22894 20052
rect 24673 20043 24731 20049
rect 24673 20040 24685 20043
rect 22888 20012 24685 20040
rect 22888 20000 22894 20012
rect 24673 20009 24685 20012
rect 24719 20009 24731 20043
rect 24673 20003 24731 20009
rect 13170 19972 13176 19984
rect 10888 19944 13176 19972
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 13262 19932 13268 19984
rect 13320 19972 13326 19984
rect 13449 19975 13507 19981
rect 13449 19972 13461 19975
rect 13320 19944 13461 19972
rect 13320 19932 13326 19944
rect 13449 19941 13461 19944
rect 13495 19941 13507 19975
rect 13449 19935 13507 19941
rect 14369 19975 14427 19981
rect 14369 19941 14381 19975
rect 14415 19972 14427 19975
rect 17865 19975 17923 19981
rect 14415 19944 17448 19972
rect 14415 19941 14427 19944
rect 14369 19935 14427 19941
rect 10505 19907 10563 19913
rect 10505 19873 10517 19907
rect 10551 19873 10563 19907
rect 10505 19867 10563 19873
rect 10870 19864 10876 19916
rect 10928 19904 10934 19916
rect 15105 19907 15163 19913
rect 15105 19904 15117 19907
rect 10928 19876 15117 19904
rect 10928 19864 10934 19876
rect 15105 19873 15117 19876
rect 15151 19873 15163 19907
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 15105 19867 15163 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 17420 19913 17448 19944
rect 17865 19941 17877 19975
rect 17911 19972 17923 19975
rect 20254 19972 20260 19984
rect 17911 19944 20260 19972
rect 17911 19941 17923 19944
rect 17865 19935 17923 19941
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 20364 19944 21496 19972
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 20364 19904 20392 19944
rect 17644 19876 20392 19904
rect 20993 19907 21051 19913
rect 17644 19864 17650 19876
rect 20993 19873 21005 19907
rect 21039 19904 21051 19907
rect 21358 19904 21364 19916
rect 21039 19876 21364 19904
rect 21039 19873 21051 19876
rect 20993 19867 21051 19873
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 7791 19808 8064 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 7300 19768 7328 19799
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 9232 19836 9260 19864
rect 9950 19836 9956 19848
rect 8352 19808 9260 19836
rect 9911 19808 9956 19836
rect 8352 19796 8358 19808
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11296 19808 11652 19836
rect 11296 19796 11302 19808
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 6472 19740 7328 19768
rect 8312 19740 10609 19768
rect 6472 19709 6500 19740
rect 6457 19703 6515 19709
rect 6457 19669 6469 19703
rect 6503 19669 6515 19703
rect 6457 19663 6515 19669
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 8312 19700 8340 19740
rect 10597 19737 10609 19740
rect 10643 19737 10655 19771
rect 10597 19731 10655 19737
rect 11149 19771 11207 19777
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11514 19768 11520 19780
rect 11195 19740 11520 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 11624 19768 11652 19808
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12345 19839 12403 19845
rect 12345 19836 12357 19839
rect 12308 19808 12357 19836
rect 12308 19796 12314 19808
rect 12345 19805 12357 19808
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 12710 19796 12716 19848
rect 12768 19796 12774 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 13596 19808 14289 19836
rect 13596 19796 13602 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 14826 19836 14832 19848
rect 14323 19808 14832 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 12728 19768 12756 19796
rect 12897 19771 12955 19777
rect 12897 19768 12909 19771
rect 11624 19740 12664 19768
rect 12728 19740 12909 19768
rect 7147 19672 8340 19700
rect 8389 19703 8447 19709
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 8389 19669 8401 19703
rect 8435 19700 8447 19703
rect 9674 19700 9680 19712
rect 8435 19672 9680 19700
rect 8435 19669 8447 19672
rect 8389 19663 8447 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 11054 19700 11060 19712
rect 9815 19672 11060 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 12161 19703 12219 19709
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 12434 19700 12440 19712
rect 12207 19672 12440 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 12636 19700 12664 19740
rect 12897 19737 12909 19740
rect 12943 19737 12955 19771
rect 12897 19731 12955 19737
rect 12989 19771 13047 19777
rect 12989 19737 13001 19771
rect 13035 19768 13047 19771
rect 13035 19740 13124 19768
rect 13035 19737 13047 19740
rect 12989 19731 13047 19737
rect 13096 19700 13124 19740
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14936 19768 14964 19799
rect 16316 19768 16344 19799
rect 17126 19796 17132 19848
rect 17184 19836 17190 19848
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 17184 19808 17233 19836
rect 17184 19796 17190 19808
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 18690 19836 18696 19848
rect 18651 19808 18696 19836
rect 17221 19799 17279 19805
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 18932 19808 19901 19836
rect 18932 19796 18938 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19836 20131 19839
rect 20898 19836 20904 19848
rect 20119 19808 20904 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21174 19836 21180 19848
rect 21135 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21468 19836 21496 19944
rect 22738 19932 22744 19984
rect 22796 19972 22802 19984
rect 23569 19975 23627 19981
rect 23569 19972 23581 19975
rect 22796 19944 23581 19972
rect 22796 19932 22802 19944
rect 23569 19941 23581 19944
rect 23615 19941 23627 19975
rect 23569 19935 23627 19941
rect 22097 19907 22155 19913
rect 22097 19873 22109 19907
rect 22143 19904 22155 19907
rect 22462 19904 22468 19916
rect 22143 19876 22468 19904
rect 22143 19873 22155 19876
rect 22097 19867 22155 19873
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 22278 19836 22284 19848
rect 21468 19808 22094 19836
rect 22239 19808 22284 19836
rect 13688 19740 14964 19768
rect 15028 19740 16344 19768
rect 13688 19728 13694 19740
rect 12636 19672 13124 19700
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 15028 19700 15056 19740
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 18414 19768 18420 19780
rect 17920 19740 18420 19768
rect 17920 19728 17926 19740
rect 18414 19728 18420 19740
rect 18472 19768 18478 19780
rect 19978 19768 19984 19780
rect 18472 19740 19984 19768
rect 18472 19728 18478 19740
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 22066 19768 22094 19808
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 23198 19836 23204 19848
rect 23159 19808 23204 19836
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19836 23443 19839
rect 23474 19836 23480 19848
rect 23431 19808 23480 19836
rect 23431 19805 23443 19808
rect 23385 19799 23443 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 23290 19768 23296 19780
rect 22066 19740 23296 19768
rect 23290 19728 23296 19740
rect 23348 19728 23354 19780
rect 13596 19672 15056 19700
rect 13596 19660 13602 19672
rect 16942 19660 16948 19712
rect 17000 19700 17006 19712
rect 17678 19700 17684 19712
rect 17000 19672 17684 19700
rect 17000 19660 17006 19672
rect 17678 19660 17684 19672
rect 17736 19700 17742 19712
rect 22094 19700 22100 19712
rect 17736 19672 22100 19700
rect 17736 19660 17742 19672
rect 22094 19660 22100 19672
rect 22152 19700 22158 19712
rect 28258 19700 28264 19712
rect 22152 19672 28264 19700
rect 22152 19660 22158 19672
rect 28258 19660 28264 19672
rect 28316 19660 28322 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19465 7159 19499
rect 7101 19459 7159 19465
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 7791 19468 8524 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 7116 19428 7144 19459
rect 8496 19428 8524 19468
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 9033 19499 9091 19505
rect 9033 19496 9045 19499
rect 8628 19468 9045 19496
rect 8628 19456 8634 19468
rect 9033 19465 9045 19468
rect 9079 19465 9091 19499
rect 9033 19459 9091 19465
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 10962 19496 10968 19508
rect 9815 19468 10968 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 11112 19468 12434 19496
rect 11112 19456 11118 19468
rect 11698 19428 11704 19440
rect 7116 19400 7972 19428
rect 8496 19400 10272 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 7944 19369 7972 19400
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 7929 19363 7987 19369
rect 7331 19332 7880 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7852 19292 7880 19332
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 8294 19360 8300 19372
rect 7929 19323 7987 19329
rect 8036 19332 8300 19360
rect 8036 19292 8064 19332
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 9122 19360 9128 19372
rect 8619 19332 9128 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9858 19360 9864 19372
rect 9723 19332 9864 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 7852 19264 8064 19292
rect 9232 19292 9260 19323
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 9232 19264 9674 19292
rect 9646 19224 9674 19264
rect 9858 19224 9864 19236
rect 9646 19196 9864 19224
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 10244 19224 10272 19400
rect 10336 19400 11704 19428
rect 10336 19233 10364 19400
rect 11698 19388 11704 19400
rect 11756 19388 11762 19440
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 11808 19400 12081 19428
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10468 19332 10517 19360
rect 10468 19320 10474 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10962 19360 10968 19372
rect 10923 19332 10968 19360
rect 10505 19323 10563 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 11808 19360 11836 19400
rect 12069 19397 12081 19400
rect 12115 19397 12127 19431
rect 12406 19428 12434 19468
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 13078 19496 13084 19508
rect 12860 19468 13084 19496
rect 12860 19456 12866 19468
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13740 19468 14412 19496
rect 13740 19428 13768 19468
rect 14384 19437 14412 19468
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 16117 19499 16175 19505
rect 16117 19496 16129 19499
rect 15620 19468 16129 19496
rect 15620 19456 15626 19468
rect 16117 19465 16129 19468
rect 16163 19465 16175 19499
rect 16117 19459 16175 19465
rect 18233 19499 18291 19505
rect 18233 19465 18245 19499
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 14277 19431 14335 19437
rect 14277 19428 14289 19431
rect 12406 19400 13768 19428
rect 13924 19400 14289 19428
rect 12069 19391 12127 19397
rect 13725 19363 13783 19369
rect 13725 19360 13737 19363
rect 11072 19332 11836 19360
rect 12636 19332 13737 19360
rect 10594 19252 10600 19304
rect 10652 19292 10658 19304
rect 11072 19292 11100 19332
rect 11974 19292 11980 19304
rect 10652 19264 11100 19292
rect 11935 19264 11980 19292
rect 10652 19252 10658 19264
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 12124 19264 12265 19292
rect 12124 19252 12130 19264
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12636 19292 12664 19332
rect 13725 19329 13737 19332
rect 13771 19329 13783 19363
rect 13924 19360 13952 19400
rect 14277 19397 14289 19400
rect 14323 19397 14335 19431
rect 14277 19391 14335 19397
rect 14369 19431 14427 19437
rect 14369 19397 14381 19431
rect 14415 19397 14427 19431
rect 14369 19391 14427 19397
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 18248 19428 18276 19459
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 18877 19499 18935 19505
rect 18877 19496 18889 19499
rect 18380 19468 18889 19496
rect 18380 19456 18386 19468
rect 18877 19465 18889 19468
rect 18923 19465 18935 19499
rect 18877 19459 18935 19465
rect 19521 19499 19579 19505
rect 19521 19465 19533 19499
rect 19567 19465 19579 19499
rect 19521 19459 19579 19465
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 20530 19496 20536 19508
rect 20211 19468 20536 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 19334 19428 19340 19440
rect 14884 19400 17724 19428
rect 18248 19400 19340 19428
rect 14884 19388 14890 19400
rect 13725 19323 13783 19329
rect 13832 19332 13952 19360
rect 12492 19264 12664 19292
rect 12492 19252 12498 19264
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 13832 19292 13860 19332
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 15252 19332 16313 19360
rect 15252 19320 15258 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 16540 19332 17601 19360
rect 16540 19320 16546 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17696 19360 17724 19400
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 19536 19428 19564 19459
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 21174 19496 21180 19508
rect 20855 19468 21180 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 22738 19496 22744 19508
rect 22699 19468 22744 19496
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 23201 19499 23259 19505
rect 23201 19465 23213 19499
rect 23247 19496 23259 19499
rect 23658 19496 23664 19508
rect 23247 19468 23664 19496
rect 23247 19465 23259 19468
rect 23201 19459 23259 19465
rect 23658 19456 23664 19468
rect 23716 19456 23722 19508
rect 23845 19499 23903 19505
rect 23845 19465 23857 19499
rect 23891 19496 23903 19499
rect 23934 19496 23940 19508
rect 23891 19468 23940 19496
rect 23891 19465 23903 19468
rect 23845 19459 23903 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 19536 19400 21036 19428
rect 18414 19360 18420 19372
rect 17696 19332 18276 19360
rect 18375 19332 18420 19360
rect 17589 19323 17647 19329
rect 13228 19264 13860 19292
rect 15105 19295 15163 19301
rect 13228 19252 13234 19264
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15286 19292 15292 19304
rect 15151 19264 15292 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 10060 19196 10272 19224
rect 10321 19227 10379 19233
rect 10060 19168 10088 19196
rect 10321 19193 10333 19227
rect 10367 19193 10379 19227
rect 10321 19187 10379 19193
rect 11057 19227 11115 19233
rect 11057 19193 11069 19227
rect 11103 19224 11115 19227
rect 11146 19224 11152 19236
rect 11103 19196 11152 19224
rect 11103 19193 11115 19196
rect 11057 19187 11115 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 15010 19184 15016 19236
rect 15068 19224 15074 19236
rect 15120 19224 15148 19255
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19261 17187 19295
rect 18248 19292 18276 19332
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18524 19332 19073 19360
rect 18524 19292 18552 19332
rect 19061 19329 19073 19332
rect 19107 19360 19119 19363
rect 19426 19360 19432 19372
rect 19107 19332 19432 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 20070 19360 20076 19372
rect 19751 19332 20076 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 20070 19320 20076 19332
rect 20128 19360 20134 19372
rect 20806 19360 20812 19372
rect 20128 19332 20812 19360
rect 20128 19320 20134 19332
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 21008 19369 21036 19400
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 22152 19332 22197 19360
rect 22152 19320 22158 19332
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23348 19332 23397 19360
rect 23348 19320 23354 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 24486 19320 24492 19372
rect 24544 19360 24550 19372
rect 28813 19363 28871 19369
rect 28813 19360 28825 19363
rect 24544 19332 28825 19360
rect 24544 19320 24550 19332
rect 28813 19329 28825 19332
rect 28859 19329 28871 19363
rect 28813 19323 28871 19329
rect 28905 19363 28963 19369
rect 28905 19329 28917 19363
rect 28951 19360 28963 19363
rect 30282 19360 30288 19372
rect 28951 19332 30288 19360
rect 28951 19329 28963 19332
rect 28905 19323 28963 19329
rect 30282 19320 30288 19332
rect 30340 19320 30346 19372
rect 18248 19264 18552 19292
rect 22281 19295 22339 19301
rect 17129 19255 17187 19261
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 22922 19292 22928 19304
rect 22327 19264 22928 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 15068 19196 15148 19224
rect 15068 19184 15074 19196
rect 16114 19184 16120 19236
rect 16172 19224 16178 19236
rect 17144 19224 17172 19255
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 16172 19196 17172 19224
rect 16172 19184 16178 19196
rect 19978 19184 19984 19236
rect 20036 19224 20042 19236
rect 20438 19224 20444 19236
rect 20036 19196 20444 19224
rect 20036 19184 20042 19196
rect 20438 19184 20444 19196
rect 20496 19224 20502 19236
rect 22186 19224 22192 19236
rect 20496 19196 22192 19224
rect 20496 19184 20502 19196
rect 22186 19184 22192 19196
rect 22244 19184 22250 19236
rect 8389 19159 8447 19165
rect 8389 19125 8401 19159
rect 8435 19156 8447 19159
rect 8570 19156 8576 19168
rect 8435 19128 8576 19156
rect 8435 19125 8447 19128
rect 8389 19119 8447 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 10042 19116 10048 19168
rect 10100 19116 10106 19168
rect 11698 19116 11704 19168
rect 11756 19156 11762 19168
rect 13170 19156 13176 19168
rect 11756 19128 13176 19156
rect 11756 19116 11762 19128
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13538 19156 13544 19168
rect 13499 19128 13544 19156
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 17310 19156 17316 19168
rect 13780 19128 17316 19156
rect 13780 19116 13786 19128
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 10551 18924 15240 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 8389 18887 8447 18893
rect 8389 18853 8401 18887
rect 8435 18884 8447 18887
rect 9674 18884 9680 18896
rect 8435 18856 9680 18884
rect 8435 18853 8447 18856
rect 8389 18847 8447 18853
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 9861 18887 9919 18893
rect 9861 18853 9873 18887
rect 9907 18853 9919 18887
rect 10060 18884 10088 18912
rect 10594 18884 10600 18896
rect 10060 18856 10600 18884
rect 9861 18847 9919 18853
rect 7190 18776 7196 18828
rect 7248 18776 7254 18828
rect 9876 18816 9904 18847
rect 10594 18844 10600 18856
rect 10652 18844 10658 18896
rect 11790 18844 11796 18896
rect 11848 18884 11854 18896
rect 13449 18887 13507 18893
rect 13449 18884 13461 18887
rect 11848 18856 13461 18884
rect 11848 18844 11854 18856
rect 13449 18853 13461 18856
rect 13495 18853 13507 18887
rect 13449 18847 13507 18853
rect 9876 18788 10732 18816
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7208 18748 7236 18776
rect 7926 18748 7932 18760
rect 7147 18720 7236 18748
rect 7887 18720 7932 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 8570 18748 8576 18760
rect 8531 18720 8576 18748
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9858 18748 9864 18760
rect 9447 18720 9864 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10704 18757 10732 18788
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 10836 18788 13277 18816
rect 10836 18776 10842 18788
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 14366 18816 14372 18828
rect 14327 18788 14372 18816
rect 13265 18779 13323 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18717 12495 18751
rect 12437 18711 12495 18717
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 14182 18748 14188 18760
rect 13127 18720 14188 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 7193 18683 7251 18689
rect 7193 18649 7205 18683
rect 7239 18680 7251 18683
rect 11238 18680 11244 18692
rect 7239 18652 11100 18680
rect 11199 18652 11244 18680
rect 7239 18649 7251 18652
rect 7193 18643 7251 18649
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 8110 18612 8116 18624
rect 7791 18584 8116 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 9217 18615 9275 18621
rect 9217 18581 9229 18615
rect 9263 18612 9275 18615
rect 10042 18612 10048 18624
rect 9263 18584 10048 18612
rect 9263 18581 9275 18584
rect 9217 18575 9275 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 11072 18612 11100 18652
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 11333 18683 11391 18689
rect 11333 18649 11345 18683
rect 11379 18649 11391 18683
rect 11333 18643 11391 18649
rect 11348 18612 11376 18643
rect 11514 18640 11520 18692
rect 11572 18680 11578 18692
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 11572 18652 11897 18680
rect 11572 18640 11578 18652
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 12452 18680 12480 18711
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 13722 18680 13728 18692
rect 12452 18652 13728 18680
rect 11885 18643 11943 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 14461 18683 14519 18689
rect 14461 18649 14473 18683
rect 14507 18649 14519 18683
rect 15212 18680 15240 18924
rect 15396 18924 18276 18952
rect 15396 18825 15424 18924
rect 18138 18884 18144 18896
rect 17144 18856 18144 18884
rect 15381 18819 15439 18825
rect 15381 18785 15393 18819
rect 15427 18785 15439 18819
rect 15381 18779 15439 18785
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 16209 18751 16267 18757
rect 16209 18748 16221 18751
rect 15344 18720 16221 18748
rect 15344 18708 15350 18720
rect 16209 18717 16221 18720
rect 16255 18717 16267 18751
rect 16209 18711 16267 18717
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18748 16451 18751
rect 17144 18748 17172 18856
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 18248 18825 18276 18924
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21545 18955 21603 18961
rect 21545 18952 21557 18955
rect 20772 18924 21557 18952
rect 20772 18912 20778 18924
rect 21545 18921 21557 18924
rect 21591 18921 21603 18955
rect 22922 18952 22928 18964
rect 22883 18924 22928 18952
rect 21545 18915 21603 18921
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 23474 18952 23480 18964
rect 23435 18924 23480 18952
rect 23474 18912 23480 18924
rect 23532 18912 23538 18964
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 19610 18884 19616 18896
rect 18380 18856 19616 18884
rect 18380 18844 18386 18856
rect 19610 18844 19616 18856
rect 19668 18844 19674 18896
rect 20993 18887 21051 18893
rect 20993 18853 21005 18887
rect 21039 18884 21051 18887
rect 22278 18884 22284 18896
rect 21039 18856 22284 18884
rect 21039 18853 21051 18856
rect 20993 18847 21051 18853
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18785 18291 18819
rect 18233 18779 18291 18785
rect 16439 18720 17172 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 17402 18680 17408 18692
rect 15212 18652 16988 18680
rect 17363 18652 17408 18680
rect 14461 18643 14519 18649
rect 12526 18612 12532 18624
rect 11072 18584 11376 18612
rect 12487 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 14476 18612 14504 18643
rect 13872 18584 14504 18612
rect 13872 18572 13878 18584
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 16298 18612 16304 18624
rect 14608 18584 16304 18612
rect 14608 18572 14614 18584
rect 16298 18572 16304 18584
rect 16356 18612 16362 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16356 18584 16865 18612
rect 16356 18572 16362 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 16960 18612 16988 18652
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 17497 18683 17555 18689
rect 17497 18649 17509 18683
rect 17543 18649 17555 18683
rect 17497 18643 17555 18649
rect 17512 18612 17540 18643
rect 16960 18584 17540 18612
rect 18248 18612 18276 18779
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19392 18788 21772 18816
rect 19392 18776 19398 18788
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 21744 18757 21772 18788
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18717 21787 18751
rect 22186 18748 22192 18760
rect 22147 18720 22192 18748
rect 21729 18711 21787 18717
rect 22186 18708 22192 18720
rect 22244 18708 22250 18760
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23290 18748 23296 18760
rect 22879 18720 23296 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 23750 18708 23756 18760
rect 23808 18748 23814 18760
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 23808 18720 29745 18748
rect 23808 18708 23814 18720
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 30282 18708 30288 18760
rect 30340 18748 30346 18760
rect 35069 18751 35127 18757
rect 35069 18748 35081 18751
rect 30340 18720 35081 18748
rect 30340 18708 30346 18720
rect 35069 18717 35081 18720
rect 35115 18717 35127 18751
rect 35069 18711 35127 18717
rect 18598 18640 18604 18692
rect 18656 18680 18662 18692
rect 19521 18683 19579 18689
rect 19521 18680 19533 18683
rect 18656 18652 19533 18680
rect 18656 18640 18662 18652
rect 19521 18649 19533 18652
rect 19567 18649 19579 18683
rect 19521 18643 19579 18649
rect 19610 18640 19616 18692
rect 19668 18680 19674 18692
rect 20162 18680 20168 18692
rect 19668 18652 19713 18680
rect 20123 18652 20168 18680
rect 19668 18640 19674 18652
rect 20162 18640 20168 18652
rect 20220 18640 20226 18692
rect 34790 18680 34796 18692
rect 20272 18652 34796 18680
rect 20272 18612 20300 18652
rect 34790 18640 34796 18652
rect 34848 18640 34854 18692
rect 18248 18584 20300 18612
rect 16853 18575 16911 18581
rect 20898 18572 20904 18624
rect 20956 18612 20962 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 20956 18584 22293 18612
rect 20956 18572 20962 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 29825 18615 29883 18621
rect 29825 18581 29837 18615
rect 29871 18612 29883 18615
rect 33042 18612 33048 18624
rect 29871 18584 33048 18612
rect 29871 18581 29883 18584
rect 29825 18575 29883 18581
rect 33042 18572 33048 18584
rect 33100 18572 33106 18624
rect 34885 18615 34943 18621
rect 34885 18581 34897 18615
rect 34931 18612 34943 18615
rect 38010 18612 38016 18624
rect 34931 18584 38016 18612
rect 34931 18581 34943 18584
rect 34885 18575 34943 18581
rect 38010 18572 38016 18584
rect 38068 18572 38074 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 5810 18408 5816 18420
rect 1627 18380 5816 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18377 9275 18411
rect 9217 18371 9275 18377
rect 9861 18411 9919 18417
rect 9861 18377 9873 18411
rect 9907 18408 9919 18411
rect 10778 18408 10784 18420
rect 9907 18380 10784 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 7374 18272 7380 18284
rect 5951 18244 7380 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18241 7527 18275
rect 8110 18272 8116 18284
rect 8071 18244 8116 18272
rect 7469 18235 7527 18241
rect 7484 18204 7512 18235
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9232 18272 9260 18371
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11020 18380 11928 18408
rect 11020 18368 11026 18380
rect 11790 18340 11796 18352
rect 11751 18312 11796 18340
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 11900 18349 11928 18380
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 16298 18408 16304 18420
rect 12584 18380 15976 18408
rect 16259 18380 16304 18408
rect 12584 18368 12590 18380
rect 11885 18343 11943 18349
rect 11885 18309 11897 18343
rect 11931 18309 11943 18343
rect 15948 18340 15976 18380
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 18598 18408 18604 18420
rect 18559 18380 18604 18408
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 26234 18408 26240 18420
rect 20180 18380 26240 18408
rect 20180 18352 20208 18380
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 15948 18312 17049 18340
rect 11885 18303 11943 18309
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 17589 18343 17647 18349
rect 17589 18309 17601 18343
rect 17635 18340 17647 18343
rect 20162 18340 20168 18352
rect 17635 18312 20168 18340
rect 17635 18309 17647 18312
rect 17589 18303 17647 18309
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 20533 18343 20591 18349
rect 20533 18309 20545 18343
rect 20579 18340 20591 18343
rect 20990 18340 20996 18352
rect 20579 18312 20996 18340
rect 20579 18309 20591 18312
rect 20533 18303 20591 18309
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 22186 18340 22192 18352
rect 22147 18312 22192 18340
rect 22186 18300 22192 18312
rect 22244 18300 22250 18352
rect 9398 18272 9404 18284
rect 8803 18244 9260 18272
rect 9359 18244 9404 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 10042 18272 10048 18284
rect 10003 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 13630 18272 13636 18284
rect 12943 18244 13636 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 15838 18272 15844 18284
rect 15799 18244 15844 18272
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 18932 18244 19257 18272
rect 18932 18232 18938 18244
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 8386 18204 8392 18216
rect 7484 18176 8392 18204
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 10502 18204 10508 18216
rect 10463 18176 10508 18204
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 12066 18204 12072 18216
rect 12027 18176 12072 18204
rect 10689 18167 10747 18173
rect 7929 18139 7987 18145
rect 7929 18105 7941 18139
rect 7975 18136 7987 18139
rect 10704 18136 10732 18167
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12802 18204 12808 18216
rect 12176 18176 12808 18204
rect 12176 18136 12204 18176
rect 12802 18164 12808 18176
rect 12860 18164 12866 18216
rect 13078 18204 13084 18216
rect 13039 18176 13084 18204
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 13228 18176 14749 18204
rect 13228 18164 13234 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16758 18204 16764 18216
rect 15703 18176 16764 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 19426 18204 19432 18216
rect 19387 18176 19432 18204
rect 16945 18167 17003 18173
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 7975 18108 10732 18136
rect 11072 18108 12204 18136
rect 12406 18108 13277 18136
rect 7975 18105 7987 18108
rect 7929 18099 7987 18105
rect 5718 18068 5724 18080
rect 5679 18040 5724 18068
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 8573 18071 8631 18077
rect 8573 18037 8585 18071
rect 8619 18068 8631 18071
rect 11072 18068 11100 18108
rect 8619 18040 11100 18068
rect 11149 18071 11207 18077
rect 8619 18037 8631 18040
rect 8573 18031 8631 18037
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11238 18068 11244 18080
rect 11195 18040 11244 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11238 18028 11244 18040
rect 11296 18068 11302 18080
rect 12406 18068 12434 18108
rect 13265 18105 13277 18108
rect 13311 18105 13323 18139
rect 13265 18099 13323 18105
rect 13998 18096 14004 18148
rect 14056 18136 14062 18148
rect 16960 18136 16988 18167
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 20254 18204 20260 18216
rect 19935 18176 20260 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 20254 18164 20260 18176
rect 20312 18204 20318 18216
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 20312 18176 20453 18204
rect 20312 18164 20318 18176
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 21453 18207 21511 18213
rect 21453 18173 21465 18207
rect 21499 18173 21511 18207
rect 21453 18167 21511 18173
rect 14056 18108 16988 18136
rect 21468 18136 21496 18167
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 23106 18204 23112 18216
rect 22152 18176 22197 18204
rect 23067 18176 23112 18204
rect 22152 18164 22158 18176
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 23124 18136 23152 18164
rect 21468 18108 23152 18136
rect 14056 18096 14062 18108
rect 11296 18040 12434 18068
rect 11296 18028 11302 18040
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13170 18068 13176 18080
rect 12952 18040 13176 18068
rect 12952 18028 12958 18040
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 15194 18068 15200 18080
rect 15155 18040 15200 18068
rect 15194 18028 15200 18040
rect 15252 18068 15258 18080
rect 15746 18068 15752 18080
rect 15252 18040 15752 18068
rect 15252 18028 15258 18040
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 24118 18068 24124 18080
rect 23440 18040 24124 18068
rect 23440 18028 23446 18040
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 18049 17867 18107 17873
rect 1912 17836 18000 17864
rect 1912 17824 1918 17836
rect 9214 17756 9220 17808
rect 9272 17796 9278 17808
rect 10502 17796 10508 17808
rect 9272 17768 10508 17796
rect 9272 17756 9278 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 11057 17799 11115 17805
rect 11057 17765 11069 17799
rect 11103 17796 11115 17799
rect 11790 17796 11796 17808
rect 11103 17768 11796 17796
rect 11103 17765 11115 17768
rect 11057 17759 11115 17765
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 14642 17796 14648 17808
rect 12584 17768 14648 17796
rect 12584 17756 12590 17768
rect 14642 17756 14648 17768
rect 14700 17756 14706 17808
rect 17972 17796 18000 17836
rect 18049 17833 18061 17867
rect 18095 17864 18107 17867
rect 19426 17864 19432 17876
rect 18095 17836 19432 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22649 17867 22707 17873
rect 22649 17864 22661 17867
rect 22244 17836 22661 17864
rect 22244 17824 22250 17836
rect 22649 17833 22661 17836
rect 22695 17833 22707 17867
rect 22649 17827 22707 17833
rect 20806 17796 20812 17808
rect 17972 17768 20812 17796
rect 20806 17756 20812 17768
rect 20864 17756 20870 17808
rect 21545 17799 21603 17805
rect 21545 17765 21557 17799
rect 21591 17796 21603 17799
rect 22370 17796 22376 17808
rect 21591 17768 22376 17796
rect 21591 17765 21603 17768
rect 21545 17759 21603 17765
rect 22370 17756 22376 17768
rect 22428 17756 22434 17808
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 8527 17700 9505 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 9732 17700 11713 17728
rect 9732 17688 9738 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 11701 17691 11759 17697
rect 11808 17700 14749 17728
rect 7282 17620 7288 17672
rect 7340 17660 7346 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7340 17632 7941 17660
rect 7340 17620 7346 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 8386 17660 8392 17672
rect 8347 17632 8392 17660
rect 7929 17623 7987 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 9272 17632 9321 17660
rect 9272 17620 9278 17632
rect 9309 17629 9321 17632
rect 9355 17629 9367 17663
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 9309 17623 9367 17629
rect 9416 17632 10425 17660
rect 8018 17552 8024 17604
rect 8076 17592 8082 17604
rect 9416 17592 9444 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10413 17623 10471 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11204 17632 11529 17660
rect 11204 17620 11210 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 11808 17660 11836 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 16482 17728 16488 17740
rect 16443 17700 16488 17728
rect 14737 17691 14795 17697
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 18831 17700 19993 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21910 17728 21916 17740
rect 20947 17700 21916 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21910 17688 21916 17700
rect 21968 17688 21974 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22094 17728 22100 17740
rect 22051 17700 22100 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 18230 17660 18236 17672
rect 11517 17623 11575 17629
rect 11624 17632 11836 17660
rect 18191 17632 18236 17660
rect 9953 17595 10011 17601
rect 9953 17592 9965 17595
rect 8076 17564 9444 17592
rect 9646 17564 9965 17592
rect 8076 17552 8082 17564
rect 7745 17527 7803 17533
rect 7745 17493 7757 17527
rect 7791 17524 7803 17527
rect 8478 17524 8484 17536
rect 7791 17496 8484 17524
rect 7791 17493 7803 17496
rect 7745 17487 7803 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8938 17484 8944 17536
rect 8996 17524 9002 17536
rect 9646 17524 9674 17564
rect 9953 17561 9965 17564
rect 9999 17592 10011 17595
rect 11624 17592 11652 17632
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 20530 17660 20536 17672
rect 19843 17632 20536 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 21082 17660 21088 17672
rect 21043 17632 21088 17660
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 22830 17660 22836 17672
rect 22791 17632 22836 17660
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 27801 17663 27859 17669
rect 27801 17660 27813 17663
rect 26384 17632 27813 17660
rect 26384 17620 26390 17632
rect 27801 17629 27813 17632
rect 27847 17629 27859 17663
rect 27801 17623 27859 17629
rect 9999 17564 11652 17592
rect 12713 17595 12771 17601
rect 9999 17561 10011 17564
rect 9953 17555 10011 17561
rect 12713 17561 12725 17595
rect 12759 17561 12771 17595
rect 12713 17555 12771 17561
rect 8996 17496 9674 17524
rect 12161 17527 12219 17533
rect 8996 17484 9002 17496
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12526 17524 12532 17536
rect 12207 17496 12532 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12729 17524 12757 17555
rect 12802 17552 12808 17604
rect 12860 17592 12866 17604
rect 12860 17564 12905 17592
rect 12860 17552 12866 17564
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 13228 17564 13369 17592
rect 13228 17552 13234 17564
rect 13357 17561 13369 17564
rect 13403 17592 13415 17595
rect 13446 17592 13452 17604
rect 13403 17564 13452 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 14826 17552 14832 17604
rect 14884 17592 14890 17604
rect 15381 17595 15439 17601
rect 14884 17564 14929 17592
rect 14884 17552 14890 17564
rect 15381 17561 15393 17595
rect 15427 17561 15439 17595
rect 15381 17555 15439 17561
rect 15102 17524 15108 17536
rect 12729 17496 15108 17524
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 15396 17524 15424 17555
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 16577 17595 16635 17601
rect 16577 17592 16589 17595
rect 15528 17564 16589 17592
rect 15528 17552 15534 17564
rect 16577 17561 16589 17564
rect 16623 17561 16635 17595
rect 16577 17555 16635 17561
rect 17129 17595 17187 17601
rect 17129 17561 17141 17595
rect 17175 17592 17187 17595
rect 17218 17592 17224 17604
rect 17175 17564 17224 17592
rect 17175 17561 17187 17564
rect 17129 17555 17187 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 18046 17524 18052 17536
rect 15396 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 27893 17527 27951 17533
rect 27893 17493 27905 17527
rect 27939 17524 27951 17527
rect 34514 17524 34520 17536
rect 27939 17496 34520 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 34514 17484 34520 17496
rect 34572 17484 34578 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 11057 17323 11115 17329
rect 7984 17292 11008 17320
rect 7984 17280 7990 17292
rect 7374 17212 7380 17264
rect 7432 17252 7438 17264
rect 10413 17255 10471 17261
rect 10413 17252 10425 17255
rect 7432 17224 10425 17252
rect 7432 17212 7438 17224
rect 10413 17221 10425 17224
rect 10459 17221 10471 17255
rect 10413 17215 10471 17221
rect 8478 17184 8484 17196
rect 8439 17156 8484 17184
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 8938 17184 8944 17196
rect 8899 17156 8944 17184
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17153 9919 17187
rect 10318 17184 10324 17196
rect 10279 17156 10324 17184
rect 9861 17147 9919 17153
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 8297 17119 8355 17125
rect 8297 17116 8309 17119
rect 7064 17088 8309 17116
rect 7064 17076 7070 17088
rect 8297 17085 8309 17088
rect 8343 17085 8355 17119
rect 9876 17116 9904 17147
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10980 17193 11008 17292
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 13078 17320 13084 17332
rect 11103 17292 13084 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 13998 17320 14004 17332
rect 13959 17292 14004 17320
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 17402 17320 17408 17332
rect 16163 17292 17408 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 20533 17323 20591 17329
rect 18248 17292 19380 17320
rect 12897 17255 12955 17261
rect 12897 17221 12909 17255
rect 12943 17252 12955 17255
rect 14016 17252 14044 17280
rect 12943 17224 14044 17252
rect 15381 17255 15439 17261
rect 12943 17221 12955 17224
rect 12897 17215 12955 17221
rect 15381 17221 15393 17255
rect 15427 17252 15439 17255
rect 16482 17252 16488 17264
rect 15427 17224 16488 17252
rect 15427 17221 15439 17224
rect 15381 17215 15439 17221
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 16758 17212 16764 17264
rect 16816 17252 16822 17264
rect 18248 17252 18276 17292
rect 16816 17224 18276 17252
rect 18325 17255 18383 17261
rect 16816 17212 16822 17224
rect 18325 17221 18337 17255
rect 18371 17252 18383 17255
rect 18371 17224 19288 17252
rect 18371 17221 18383 17224
rect 18325 17215 18383 17221
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 11112 17156 13553 17184
rect 11112 17144 11118 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 10870 17116 10876 17128
rect 9876 17088 10876 17116
rect 8297 17079 8355 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 11848 17088 12265 17116
rect 11848 17076 11854 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 9677 17051 9735 17057
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 12452 17048 12480 17079
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 14274 17116 14280 17128
rect 13412 17088 14280 17116
rect 13412 17076 13418 17088
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17085 14795 17119
rect 14918 17116 14924 17128
rect 14879 17088 14924 17116
rect 14737 17079 14795 17085
rect 9723 17020 12480 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 14752 16980 14780 17079
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17116 17279 17119
rect 17862 17116 17868 17128
rect 17267 17088 17868 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 17052 17048 17080 17079
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18966 17116 18972 17128
rect 18279 17088 18972 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 18690 17048 18696 17060
rect 17052 17020 18696 17048
rect 18690 17008 18696 17020
rect 18748 17008 18754 17060
rect 18785 17051 18843 17057
rect 18785 17017 18797 17051
rect 18831 17017 18843 17051
rect 19260 17048 19288 17224
rect 19352 17193 19380 17292
rect 20533 17289 20545 17323
rect 20579 17320 20591 17323
rect 21082 17320 21088 17332
rect 20579 17292 21088 17320
rect 20579 17289 20591 17292
rect 20533 17283 20591 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 22005 17323 22063 17329
rect 22005 17289 22017 17323
rect 22051 17320 22063 17323
rect 22830 17320 22836 17332
rect 22051 17292 22836 17320
rect 22051 17289 22063 17292
rect 22005 17283 22063 17289
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 20990 17212 20996 17264
rect 21048 17252 21054 17264
rect 21177 17255 21235 17261
rect 21177 17252 21189 17255
rect 21048 17224 21189 17252
rect 21048 17212 21054 17224
rect 21177 17221 21189 17224
rect 21223 17221 21235 17255
rect 21177 17215 21235 17221
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20438 17184 20444 17196
rect 19668 17156 20444 17184
rect 19668 17144 19674 17156
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20864 17156 21097 17184
rect 20864 17144 20870 17156
rect 21085 17153 21097 17156
rect 21131 17184 21143 17187
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 21131 17156 22201 17184
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 22189 17153 22201 17156
rect 22235 17153 22247 17187
rect 38010 17184 38016 17196
rect 37971 17156 38016 17184
rect 22189 17147 22247 17153
rect 38010 17144 38016 17156
rect 38068 17144 38074 17196
rect 19518 17116 19524 17128
rect 19479 17088 19524 17116
rect 19518 17076 19524 17088
rect 19576 17076 19582 17128
rect 19886 17048 19892 17060
rect 19260 17020 19892 17048
rect 18785 17011 18843 17017
rect 10560 16952 14780 16980
rect 10560 16940 10566 16952
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 17402 16980 17408 16992
rect 15160 16952 17408 16980
rect 15160 16940 15166 16952
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 18800 16980 18828 17011
rect 19886 17008 19892 17020
rect 19944 17008 19950 17060
rect 19981 17051 20039 17057
rect 19981 17017 19993 17051
rect 20027 17048 20039 17051
rect 22370 17048 22376 17060
rect 20027 17020 22376 17048
rect 20027 17017 20039 17020
rect 19981 17011 20039 17017
rect 22370 17008 22376 17020
rect 22428 17008 22434 17060
rect 38194 17048 38200 17060
rect 38155 17020 38200 17048
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 22002 16980 22008 16992
rect 18104 16952 22008 16980
rect 18104 16940 18110 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 15194 16776 15200 16788
rect 10376 16748 15200 16776
rect 10376 16736 10382 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 17460 16748 17877 16776
rect 17460 16736 17466 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18288 16748 18613 16776
rect 18288 16736 18294 16748
rect 18601 16745 18613 16748
rect 18647 16745 18659 16779
rect 18601 16739 18659 16745
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 19576 16748 20085 16776
rect 19576 16736 19582 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 11330 16708 11336 16720
rect 10612 16680 11336 16708
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9364 16544 9505 16572
rect 9364 16532 9370 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10410 16572 10416 16584
rect 9999 16544 10416 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10612 16581 10640 16680
rect 11330 16668 11336 16680
rect 11388 16668 11394 16720
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 19242 16708 19248 16720
rect 13596 16680 14688 16708
rect 13596 16668 13602 16680
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 12526 16640 12532 16652
rect 11287 16612 12532 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 12526 16600 12532 16612
rect 12584 16640 12590 16652
rect 12986 16640 12992 16652
rect 12584 16612 12992 16640
rect 12584 16600 12590 16612
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 14458 16640 14464 16652
rect 14419 16612 14464 16640
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 14660 16649 14688 16680
rect 17512 16680 19248 16708
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15841 16643 15899 16649
rect 15841 16640 15853 16643
rect 15160 16612 15853 16640
rect 15160 16600 15166 16612
rect 15841 16609 15853 16612
rect 15887 16609 15899 16643
rect 15841 16603 15899 16609
rect 16485 16643 16543 16649
rect 16485 16609 16497 16643
rect 16531 16640 16543 16643
rect 17218 16640 17224 16652
rect 16531 16612 17224 16640
rect 16531 16609 16543 16612
rect 16485 16603 16543 16609
rect 17218 16600 17224 16612
rect 17276 16640 17282 16652
rect 17512 16649 17540 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 17497 16643 17555 16649
rect 17276 16612 17448 16640
rect 17276 16600 17282 16612
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 11054 16572 11060 16584
rect 10735 16544 11060 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12710 16572 12716 16584
rect 12492 16544 12716 16572
rect 12492 16532 12498 16544
rect 12710 16532 12716 16544
rect 12768 16572 12774 16584
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12768 16544 13093 16572
rect 12768 16532 12774 16544
rect 13081 16541 13093 16544
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 15286 16572 15292 16584
rect 13587 16544 15292 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 17420 16572 17448 16612
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17678 16640 17684 16652
rect 17639 16612 17684 16640
rect 17497 16603 17555 16609
rect 17678 16600 17684 16612
rect 17736 16600 17742 16652
rect 23566 16640 23572 16652
rect 17788 16612 23572 16640
rect 17788 16572 17816 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 35802 16640 35808 16652
rect 26292 16612 27200 16640
rect 26292 16600 26298 16612
rect 18782 16572 18788 16584
rect 17420 16544 17816 16572
rect 18743 16544 18788 16572
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19610 16572 19616 16584
rect 19571 16544 19616 16572
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16504 10103 16507
rect 10962 16504 10968 16516
rect 10091 16476 10968 16504
rect 10091 16473 10103 16476
rect 10045 16467 10103 16473
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 12912 16476 15240 16504
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9950 16436 9956 16448
rect 9355 16408 9956 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 10376 16408 11897 16436
rect 10376 16396 10382 16408
rect 11885 16405 11897 16408
rect 11931 16436 11943 16439
rect 12802 16436 12808 16448
rect 11931 16408 12808 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 12912 16445 12940 16476
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16405 12955 16439
rect 15102 16436 15108 16448
rect 15063 16408 15108 16436
rect 12897 16399 12955 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15212 16436 15240 16476
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 15933 16507 15991 16513
rect 15933 16504 15945 16507
rect 15436 16476 15945 16504
rect 15436 16464 15442 16476
rect 15933 16473 15945 16476
rect 15979 16473 15991 16507
rect 20272 16504 20300 16535
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 27172 16581 27200 16612
rect 33612 16612 35808 16640
rect 33612 16581 33640 16612
rect 35802 16600 35808 16612
rect 35860 16600 35866 16652
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20404 16544 20913 16572
rect 20404 16532 20410 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 27157 16575 27215 16581
rect 27157 16541 27169 16575
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 33597 16575 33655 16581
rect 33597 16541 33609 16575
rect 33643 16574 33655 16575
rect 33643 16546 33677 16574
rect 33643 16541 33655 16546
rect 33597 16535 33655 16541
rect 15933 16467 15991 16473
rect 19444 16476 20300 16504
rect 16298 16436 16304 16448
rect 15212 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 19444 16445 19472 16476
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 19886 16396 19892 16448
rect 19944 16436 19950 16448
rect 20717 16439 20775 16445
rect 20717 16436 20729 16439
rect 19944 16408 20729 16436
rect 19944 16396 19950 16408
rect 20717 16405 20729 16408
rect 20763 16405 20775 16439
rect 20717 16399 20775 16405
rect 27249 16439 27307 16445
rect 27249 16405 27261 16439
rect 27295 16436 27307 16439
rect 33502 16436 33508 16448
rect 27295 16408 33508 16436
rect 27295 16405 27307 16408
rect 27249 16399 27307 16405
rect 33502 16396 33508 16408
rect 33560 16396 33566 16448
rect 33686 16436 33692 16448
rect 33647 16408 33692 16436
rect 33686 16396 33692 16408
rect 33744 16396 33750 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9214 16232 9220 16244
rect 8987 16204 9220 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10594 16232 10600 16244
rect 10459 16204 10600 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 10928 16204 10977 16232
rect 10928 16192 10934 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 12802 16192 12808 16244
rect 12860 16192 12866 16244
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 15102 16232 15108 16244
rect 13587 16204 15108 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16201 17739 16235
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 17681 16195 17739 16201
rect 12820 16164 12848 16192
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 12820 16136 14105 16164
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 14093 16127 14151 16133
rect 14182 16124 14188 16176
rect 14240 16164 14246 16176
rect 15562 16164 15568 16176
rect 14240 16136 14285 16164
rect 15523 16136 15568 16164
rect 14240 16124 14246 16136
rect 15562 16124 15568 16136
rect 15620 16124 15626 16176
rect 17696 16164 17724 16195
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18966 16232 18972 16244
rect 18927 16204 18972 16232
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 33686 16232 33692 16244
rect 20588 16204 33692 16232
rect 20588 16192 20594 16204
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 35802 16192 35808 16244
rect 35860 16232 35866 16244
rect 38105 16235 38163 16241
rect 38105 16232 38117 16235
rect 35860 16204 38117 16232
rect 35860 16192 35866 16204
rect 38105 16201 38117 16204
rect 38151 16201 38163 16235
rect 38105 16195 38163 16201
rect 17696 16136 18552 16164
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 5718 16096 5724 16108
rect 1627 16068 5724 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 8846 16096 8852 16108
rect 8807 16068 8852 16096
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9493 16099 9551 16105
rect 9493 16096 9505 16099
rect 9364 16068 9505 16096
rect 9364 16056 9370 16068
rect 9493 16065 9505 16068
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9916 16068 10333 16096
rect 9916 16056 9922 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11330 16096 11336 16108
rect 11195 16068 11336 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12342 16096 12348 16108
rect 12023 16068 12348 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12342 16056 12348 16068
rect 12400 16096 12406 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12400 16068 12449 16096
rect 12400 16056 12406 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16724 16068 17049 16096
rect 16724 16056 16730 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17310 16056 17316 16108
rect 17368 16096 17374 16108
rect 18524 16105 18552 16136
rect 18690 16124 18696 16176
rect 18748 16164 18754 16176
rect 19613 16167 19671 16173
rect 19613 16164 19625 16167
rect 18748 16136 19625 16164
rect 18748 16124 18754 16136
rect 19613 16133 19625 16136
rect 19659 16133 19671 16167
rect 19613 16127 19671 16133
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17368 16068 17877 16096
rect 17368 16056 17374 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16065 18567 16099
rect 20438 16096 20444 16108
rect 20399 16068 20444 16096
rect 18509 16059 18567 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 22554 16056 22560 16108
rect 22612 16096 22618 16108
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 22612 16068 31585 16096
rect 22612 16056 22618 16068
rect 31573 16065 31585 16068
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 33502 16056 33508 16108
rect 33560 16096 33566 16108
rect 33597 16099 33655 16105
rect 33597 16096 33609 16099
rect 33560 16068 33609 16096
rect 33560 16056 33566 16068
rect 33597 16065 33609 16068
rect 33643 16065 33655 16099
rect 38286 16096 38292 16108
rect 38247 16068 38292 16096
rect 33597 16059 33655 16065
rect 38286 16056 38292 16068
rect 38344 16056 38350 16108
rect 12894 16028 12900 16040
rect 12855 16000 12900 16028
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 11698 15920 11704 15972
rect 11756 15960 11762 15972
rect 13096 15960 13124 15991
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 13228 16000 15485 16028
rect 13228 15988 13234 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 17402 16028 17408 16040
rect 16163 16000 17408 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 11756 15932 13124 15960
rect 11756 15920 11762 15932
rect 13262 15920 13268 15972
rect 13320 15960 13326 15972
rect 14182 15960 14188 15972
rect 13320 15932 14188 15960
rect 13320 15920 13326 15932
rect 14182 15920 14188 15932
rect 14240 15920 14246 15972
rect 14645 15963 14703 15969
rect 14645 15929 14657 15963
rect 14691 15960 14703 15963
rect 16132 15960 16160 15991
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 14691 15932 16160 15960
rect 14691 15929 14703 15932
rect 14645 15923 14703 15929
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9585 15895 9643 15901
rect 9585 15892 9597 15895
rect 9364 15864 9597 15892
rect 9364 15852 9370 15864
rect 9585 15861 9597 15864
rect 9631 15861 9643 15895
rect 9585 15855 9643 15861
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 13906 15892 13912 15904
rect 12299 15864 13912 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 16853 15895 16911 15901
rect 16853 15861 16865 15895
rect 16899 15892 16911 15895
rect 18230 15892 18236 15904
rect 16899 15864 18236 15892
rect 16899 15861 16911 15864
rect 16853 15855 16911 15861
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 20257 15895 20315 15901
rect 20257 15892 20269 15895
rect 19668 15864 20269 15892
rect 19668 15852 19674 15864
rect 20257 15861 20269 15864
rect 20303 15861 20315 15895
rect 20257 15855 20315 15861
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 33318 15892 33324 15904
rect 31711 15864 33324 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 33318 15852 33324 15864
rect 33376 15852 33382 15904
rect 33413 15895 33471 15901
rect 33413 15861 33425 15895
rect 33459 15892 33471 15895
rect 35342 15892 35348 15904
rect 33459 15864 35348 15892
rect 33459 15861 33471 15864
rect 33413 15855 33471 15861
rect 35342 15852 35348 15864
rect 35400 15852 35406 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 9769 15691 9827 15697
rect 9769 15657 9781 15691
rect 9815 15688 9827 15691
rect 10318 15688 10324 15700
rect 9815 15660 10324 15688
rect 9815 15657 9827 15660
rect 9769 15651 9827 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 11422 15688 11428 15700
rect 10459 15660 11428 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15688 12311 15691
rect 13538 15688 13544 15700
rect 12299 15660 13544 15688
rect 12299 15657 12311 15660
rect 12253 15651 12311 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 13814 15688 13820 15700
rect 13679 15660 13820 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 15470 15688 15476 15700
rect 14599 15660 15476 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 18417 15691 18475 15697
rect 18417 15688 18429 15691
rect 18196 15660 18429 15688
rect 18196 15648 18202 15660
rect 18417 15657 18429 15660
rect 18463 15657 18475 15691
rect 18417 15651 18475 15657
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 17512 15592 19441 15620
rect 9306 15552 9312 15564
rect 9267 15524 9312 15552
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13170 15552 13176 15564
rect 12943 15524 13176 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 15105 15555 15163 15561
rect 15105 15521 15117 15555
rect 15151 15552 15163 15555
rect 15930 15552 15936 15564
rect 15151 15524 15936 15552
rect 15151 15521 15163 15524
rect 15105 15515 15163 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16758 15512 16764 15564
rect 16816 15552 16822 15564
rect 16942 15552 16948 15564
rect 16816 15524 16948 15552
rect 16816 15512 16822 15524
rect 16942 15512 16948 15524
rect 17000 15552 17006 15564
rect 17512 15561 17540 15592
rect 19429 15589 19441 15592
rect 19475 15589 19487 15623
rect 19429 15583 19487 15589
rect 17313 15555 17371 15561
rect 17313 15552 17325 15555
rect 17000 15524 17325 15552
rect 17000 15512 17006 15524
rect 17313 15521 17325 15524
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10008 15456 10609 15484
rect 10008 15444 10014 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 11624 15416 11652 15447
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12492 15456 12537 15484
rect 12492 15444 12498 15456
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 12676 15456 13553 15484
rect 12676 15444 12682 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14424 15456 14473 15484
rect 14424 15444 14430 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 15286 15484 15292 15496
rect 15247 15456 15292 15484
rect 14461 15447 14519 15453
rect 12710 15416 12716 15428
rect 11624 15388 12716 15416
rect 12710 15376 12716 15388
rect 12768 15376 12774 15428
rect 14476 15416 14504 15447
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16209 15447 16267 15453
rect 15654 15416 15660 15428
rect 14476 15388 15660 15416
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 16224 15416 16252 15447
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18288 15456 18613 15484
rect 18288 15444 18294 15456
rect 18601 15453 18613 15456
rect 18647 15453 18659 15487
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 18601 15447 18659 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 33042 15444 33048 15496
rect 33100 15484 33106 15496
rect 35069 15487 35127 15493
rect 35069 15484 35081 15487
rect 33100 15456 35081 15484
rect 33100 15444 33106 15456
rect 35069 15453 35081 15456
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 17954 15416 17960 15428
rect 16224 15388 17960 15416
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 16022 15348 16028 15360
rect 15795 15320 16028 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 16022 15308 16028 15320
rect 16080 15348 16086 15360
rect 16853 15351 16911 15357
rect 16853 15348 16865 15351
rect 16080 15320 16865 15348
rect 16080 15308 16086 15320
rect 16853 15317 16865 15320
rect 16899 15317 16911 15351
rect 16853 15311 16911 15317
rect 34885 15351 34943 15357
rect 34885 15317 34897 15351
rect 34931 15348 34943 15351
rect 38010 15348 38016 15360
rect 34931 15320 38016 15348
rect 34931 15317 34943 15320
rect 34885 15311 34943 15317
rect 38010 15308 38016 15320
rect 38068 15308 38074 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 7653 15147 7711 15153
rect 7653 15113 7665 15147
rect 7699 15144 7711 15147
rect 11146 15144 11152 15156
rect 7699 15116 11152 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12492 15116 12909 15144
rect 12492 15104 12498 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 13541 15147 13599 15153
rect 13541 15113 13553 15147
rect 13587 15113 13599 15147
rect 13541 15107 13599 15113
rect 14277 15147 14335 15153
rect 14277 15113 14289 15147
rect 14323 15144 14335 15147
rect 14918 15144 14924 15156
rect 14323 15116 14924 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 12345 15079 12403 15085
rect 12345 15045 12357 15079
rect 12391 15076 12403 15079
rect 13262 15076 13268 15088
rect 12391 15048 13268 15076
rect 12391 15045 12403 15048
rect 12345 15039 12403 15045
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 13556 15076 13584 15107
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 16114 15144 16120 15156
rect 16075 15116 16120 15144
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 17954 15144 17960 15156
rect 17915 15116 17960 15144
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 15562 15076 15568 15088
rect 13556 15048 15568 15076
rect 15562 15036 15568 15048
rect 15620 15036 15626 15088
rect 6914 15008 6920 15020
rect 6875 14980 6920 15008
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 15008 12311 15011
rect 12299 14980 12434 15008
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 12406 14872 12434 14980
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12768 14980 13093 15008
rect 12768 14968 12774 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13096 14940 13124 14971
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 13596 14980 13737 15008
rect 13596 14968 13602 14980
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15470 15008 15476 15020
rect 15059 14980 15476 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 14200 14940 14228 14971
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 14977 15715 15011
rect 16298 15008 16304 15020
rect 16259 14980 16304 15008
rect 15657 14971 15715 14977
rect 13096 14912 14228 14940
rect 14734 14900 14740 14952
rect 14792 14940 14798 14952
rect 15672 14940 15700 14971
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 18598 15008 18604 15020
rect 18559 14980 18604 15008
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 17310 14940 17316 14952
rect 14792 14912 15700 14940
rect 17271 14912 17316 14940
rect 14792 14900 14798 14912
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 17494 14940 17500 14952
rect 17455 14912 17500 14940
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 13722 14872 13728 14884
rect 12406 14844 13728 14872
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14872 14887 14875
rect 15378 14872 15384 14884
rect 14875 14844 15384 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 15473 14875 15531 14881
rect 15473 14841 15485 14875
rect 15519 14872 15531 14875
rect 20346 14872 20352 14884
rect 15519 14844 20352 14872
rect 15519 14841 15531 14844
rect 15473 14835 15531 14841
rect 20346 14832 20352 14844
rect 20404 14832 20410 14884
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 18104 14776 18429 14804
rect 18104 14764 18110 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 8846 14600 8852 14612
rect 1627 14572 8852 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 14921 14603 14979 14609
rect 14921 14600 14933 14603
rect 14884 14572 14933 14600
rect 14884 14560 14890 14572
rect 14921 14569 14933 14572
rect 14967 14569 14979 14603
rect 15470 14600 15476 14612
rect 15431 14572 15476 14600
rect 14921 14563 14979 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16301 14603 16359 14609
rect 16301 14600 16313 14603
rect 15896 14572 16313 14600
rect 15896 14560 15902 14572
rect 16301 14569 16313 14572
rect 16347 14569 16359 14603
rect 16301 14563 16359 14569
rect 17313 14603 17371 14609
rect 17313 14569 17325 14603
rect 17359 14600 17371 14603
rect 17678 14600 17684 14612
rect 17359 14572 17684 14600
rect 17359 14569 17371 14572
rect 17313 14563 17371 14569
rect 17678 14560 17684 14572
rect 17736 14560 17742 14612
rect 17862 14600 17868 14612
rect 17823 14572 17868 14600
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 18598 14464 18604 14476
rect 10284 14436 18604 14464
rect 10284 14424 10290 14436
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 13722 14396 13728 14408
rect 13683 14368 13728 14396
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14792 14368 14841 14396
rect 14792 14356 14798 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 14829 14359 14887 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16666 14396 16672 14408
rect 16255 14368 16672 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17236 14405 17264 14436
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 28902 14464 28908 14476
rect 19300 14436 28908 14464
rect 19300 14424 19306 14436
rect 28902 14424 28908 14436
rect 28960 14424 28966 14476
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14365 17279 14399
rect 18046 14396 18052 14408
rect 18007 14368 18052 14396
rect 17221 14359 17279 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 35069 14399 35127 14405
rect 35069 14396 35081 14399
rect 34572 14368 35081 14396
rect 34572 14356 34578 14368
rect 35069 14365 35081 14368
rect 35115 14365 35127 14399
rect 35069 14359 35127 14365
rect 35342 14356 35348 14408
rect 35400 14396 35406 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 35400 14368 38025 14396
rect 35400 14356 35406 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 34885 14263 34943 14269
rect 34885 14229 34897 14263
rect 34931 14260 34943 14263
rect 37274 14260 37280 14272
rect 34931 14232 37280 14260
rect 34931 14229 34943 14232
rect 34885 14223 34943 14229
rect 37274 14220 37280 14232
rect 37332 14220 37338 14272
rect 38194 14260 38200 14272
rect 38155 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 14516 14028 14565 14056
rect 14516 14016 14522 14028
rect 14553 14025 14565 14028
rect 14599 14025 14611 14059
rect 15286 14056 15292 14068
rect 15247 14028 15292 14056
rect 14553 14019 14611 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15930 14056 15936 14068
rect 15891 14028 15936 14056
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 17129 14059 17187 14065
rect 17129 14025 17141 14059
rect 17175 14056 17187 14059
rect 17494 14056 17500 14068
rect 17175 14028 17500 14056
rect 17175 14025 17187 14028
rect 17129 14019 17187 14025
rect 17494 14016 17500 14028
rect 17552 14016 17558 14068
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 13964 13892 15485 13920
rect 13964 13880 13970 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 17034 13920 17040 13932
rect 16995 13892 17040 13920
rect 15473 13883 15531 13889
rect 17034 13880 17040 13892
rect 17092 13920 17098 13932
rect 20438 13920 20444 13932
rect 17092 13892 20444 13920
rect 17092 13880 17098 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16390 13512 16396 13524
rect 16163 13484 16396 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 7926 13308 7932 13320
rect 7887 13280 7932 13308
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15252 13280 16037 13308
rect 15252 13268 15258 13280
rect 16025 13277 16037 13280
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 6914 12968 6920 12980
rect 1627 12940 6920 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 13078 12832 13084 12844
rect 7975 12804 13084 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19058 12832 19064 12844
rect 18647 12804 19064 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12832 23719 12835
rect 23842 12832 23848 12844
rect 23707 12804 23848 12832
rect 23707 12801 23719 12804
rect 23661 12795 23719 12801
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 33318 12792 33324 12844
rect 33376 12832 33382 12844
rect 35529 12835 35587 12841
rect 35529 12832 35541 12835
rect 33376 12804 35541 12832
rect 33376 12792 33382 12804
rect 35529 12801 35541 12804
rect 35575 12801 35587 12835
rect 38010 12832 38016 12844
rect 37971 12804 38016 12832
rect 35529 12795 35587 12801
rect 38010 12792 38016 12804
rect 38068 12792 38074 12844
rect 5442 12588 5448 12640
rect 5500 12628 5506 12640
rect 8021 12631 8079 12637
rect 8021 12628 8033 12631
rect 5500 12600 8033 12628
rect 5500 12588 5506 12600
rect 8021 12597 8033 12600
rect 8067 12597 8079 12631
rect 18690 12628 18696 12640
rect 18651 12600 18696 12628
rect 8021 12591 8079 12597
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 23753 12631 23811 12637
rect 23753 12597 23765 12631
rect 23799 12628 23811 12631
rect 24670 12628 24676 12640
rect 23799 12600 24676 12628
rect 23799 12597 23811 12600
rect 23753 12591 23811 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 35342 12628 35348 12640
rect 35303 12600 35348 12628
rect 35342 12588 35348 12600
rect 35400 12588 35406 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 6454 12424 6460 12436
rect 6415 12396 6460 12424
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16632 12192 17141 12220
rect 16632 12180 16638 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 33413 12223 33471 12229
rect 33413 12189 33425 12223
rect 33459 12220 33471 12223
rect 38102 12220 38108 12232
rect 33459 12192 38108 12220
rect 33459 12189 33471 12192
rect 33413 12183 33471 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 18322 12084 18328 12096
rect 17267 12056 18328 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 33505 12087 33563 12093
rect 33505 12084 33517 12087
rect 21968 12056 33517 12084
rect 21968 12044 21974 12056
rect 33505 12053 33517 12056
rect 33551 12053 33563 12087
rect 33505 12047 33563 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 22370 11812 22376 11824
rect 13320 11784 22376 11812
rect 13320 11772 13326 11784
rect 22370 11772 22376 11784
rect 22428 11772 22434 11824
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 13446 11744 13452 11756
rect 5684 11716 13452 11744
rect 5684 11704 5690 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 37918 11744 37924 11756
rect 32355 11716 37924 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 37918 11704 37924 11716
rect 37976 11704 37982 11756
rect 24394 11500 24400 11552
rect 24452 11540 24458 11552
rect 32401 11543 32459 11549
rect 32401 11540 32413 11543
rect 24452 11512 32413 11540
rect 24452 11500 24458 11512
rect 32401 11509 32413 11512
rect 32447 11509 32459 11543
rect 32401 11503 32459 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 7558 11336 7564 11348
rect 1627 11308 7564 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 38194 11268 38200 11280
rect 38155 11240 38200 11268
rect 38194 11228 38200 11240
rect 38252 11228 38258 11280
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 20530 11132 20536 11144
rect 19475 11104 20536 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 38013 11135 38071 11141
rect 38013 11132 38025 11135
rect 37332 11104 38025 11132
rect 37332 11092 37338 11104
rect 38013 11101 38025 11104
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 19521 11067 19579 11073
rect 19521 11033 19533 11067
rect 19567 11064 19579 11067
rect 21174 11064 21180 11076
rect 19567 11036 21180 11064
rect 19567 11033 19579 11036
rect 19521 11027 19579 11033
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 22002 10684 22008 10736
rect 22060 10724 22066 10736
rect 22060 10696 26234 10724
rect 22060 10684 22066 10696
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11572 10628 11713 10656
rect 11572 10616 11578 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 11701 10619 11759 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17460 10628 18153 10656
rect 17460 10616 17466 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 23566 10656 23572 10668
rect 23527 10628 23572 10656
rect 18141 10619 18199 10625
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 26206 10656 26234 10696
rect 26421 10659 26479 10665
rect 26421 10656 26433 10659
rect 26206 10628 26433 10656
rect 26421 10625 26433 10628
rect 26467 10625 26479 10659
rect 26421 10619 26479 10625
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 11882 10452 11888 10464
rect 11839 10424 11888 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 15344 10424 16129 10452
rect 15344 10412 15350 10424
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16117 10415 16175 10421
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 20254 10452 20260 10464
rect 18279 10424 20260 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 23661 10455 23719 10461
rect 23661 10421 23673 10455
rect 23707 10452 23719 10455
rect 25590 10452 25596 10464
rect 23707 10424 25596 10452
rect 23707 10421 23719 10424
rect 23661 10415 23719 10421
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 26513 10455 26571 10461
rect 26513 10421 26525 10455
rect 26559 10452 26571 10455
rect 28350 10452 28356 10464
rect 26559 10424 28356 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 7926 10248 7932 10260
rect 1627 10220 7932 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 5442 10044 5448 10056
rect 4203 10016 5448 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 12066 10044 12072 10056
rect 10735 10016 12072 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 3970 9908 3976 9920
rect 3931 9880 3976 9908
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 9732 9880 10793 9908
rect 9732 9868 9738 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 13265 9163 13323 9169
rect 13265 9129 13277 9163
rect 13311 9160 13323 9163
rect 16942 9160 16948 9172
rect 13311 9132 16948 9160
rect 13311 9129 13323 9132
rect 13265 9123 13323 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 18233 9163 18291 9169
rect 18233 9129 18245 9163
rect 18279 9160 18291 9163
rect 21358 9160 21364 9172
rect 18279 9132 21364 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 13170 8956 13176 8968
rect 13131 8928 13176 8956
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 18138 8956 18144 8968
rect 18099 8928 18144 8956
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 35400 8928 38025 8956
rect 35400 8916 35406 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 11793 8619 11851 8625
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 12802 8616 12808 8628
rect 11839 8588 12808 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 22370 8616 22376 8628
rect 22331 8588 22376 8616
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 9585 8551 9643 8557
rect 9585 8517 9597 8551
rect 9631 8548 9643 8551
rect 12618 8548 12624 8560
rect 9631 8520 12624 8548
rect 9631 8517 9643 8520
rect 9585 8511 9643 8517
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 9490 8480 9496 8492
rect 9451 8452 9496 8480
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 22002 8480 22008 8492
rect 19291 8452 22008 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 11716 8412 11744 8443
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8480 22431 8483
rect 24854 8480 24860 8492
rect 22419 8452 24860 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 2372 8384 11744 8412
rect 2372 8372 2378 8384
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 6362 8072 6368 8084
rect 1627 8044 6368 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13630 8072 13636 8084
rect 13587 8044 13636 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 26973 8075 27031 8081
rect 26973 8072 26985 8075
rect 24176 8044 26985 8072
rect 24176 8032 24182 8044
rect 26973 8041 26985 8044
rect 27019 8041 27031 8075
rect 38102 8072 38108 8084
rect 38063 8044 38108 8072
rect 26973 8035 27031 8041
rect 38102 8032 38108 8044
rect 38160 8032 38166 8084
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8352 7840 9137 7868
rect 8352 7828 8358 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 14274 7868 14280 7880
rect 13495 7840 14280 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 26881 7871 26939 7877
rect 26881 7837 26893 7871
rect 26927 7868 26939 7871
rect 28626 7868 28632 7880
rect 26927 7840 28632 7868
rect 26927 7837 26939 7840
rect 26881 7831 26939 7837
rect 28626 7828 28632 7840
rect 28684 7828 28690 7880
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 35253 7871 35311 7877
rect 35253 7868 35265 7871
rect 34848 7840 35265 7868
rect 34848 7828 34854 7840
rect 35253 7837 35265 7840
rect 35299 7837 35311 7871
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 35253 7831 35311 7837
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 9217 7803 9275 7809
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 9263 7772 16574 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 16546 7732 16574 7772
rect 17126 7732 17132 7744
rect 16546 7704 17132 7732
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 35345 7735 35403 7741
rect 35345 7701 35357 7735
rect 35391 7732 35403 7735
rect 37090 7732 37096 7744
rect 35391 7704 37096 7732
rect 35391 7701 35403 7704
rect 35345 7695 35403 7701
rect 37090 7692 37096 7704
rect 37148 7692 37154 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 34241 7395 34299 7401
rect 34241 7361 34253 7395
rect 34287 7392 34299 7395
rect 35802 7392 35808 7404
rect 34287 7364 35808 7392
rect 34287 7361 34299 7364
rect 34241 7355 34299 7361
rect 35802 7352 35808 7364
rect 35860 7352 35866 7404
rect 22462 7148 22468 7200
rect 22520 7188 22526 7200
rect 34333 7191 34391 7197
rect 34333 7188 34345 7191
rect 22520 7160 34345 7188
rect 22520 7148 22526 7160
rect 34333 7157 34345 7160
rect 34379 7157 34391 7191
rect 34333 7151 34391 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 21450 6944 21456 6996
rect 21508 6984 21514 6996
rect 24765 6987 24823 6993
rect 24765 6984 24777 6987
rect 21508 6956 24777 6984
rect 21508 6944 21514 6956
rect 24765 6953 24777 6956
rect 24811 6953 24823 6987
rect 24765 6947 24823 6953
rect 24673 6783 24731 6789
rect 24673 6749 24685 6783
rect 24719 6780 24731 6783
rect 25406 6780 25412 6792
rect 24719 6752 25412 6780
rect 24719 6749 24731 6752
rect 24673 6743 24731 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 28902 6440 28908 6452
rect 28863 6412 28908 6440
rect 28902 6400 28908 6412
rect 28960 6400 28966 6452
rect 8757 6375 8815 6381
rect 8757 6341 8769 6375
rect 8803 6372 8815 6375
rect 12894 6372 12900 6384
rect 8803 6344 12900 6372
rect 8803 6341 8815 6344
rect 8757 6335 8815 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 3970 6304 3976 6316
rect 1627 6276 3976 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 4764 6276 8677 6304
rect 4764 6264 4770 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11204 6276 11713 6304
rect 11204 6264 11210 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 28813 6307 28871 6313
rect 28813 6273 28825 6307
rect 28859 6304 28871 6307
rect 30282 6304 30288 6316
rect 28859 6276 30288 6304
rect 28859 6273 28871 6276
rect 28813 6267 28871 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 38102 6304 38108 6316
rect 38063 6276 38108 6304
rect 38102 6264 38108 6276
rect 38160 6264 38166 6316
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 37274 6060 37280 6112
rect 37332 6100 37338 6112
rect 38197 6103 38255 6109
rect 38197 6100 38209 6103
rect 37332 6072 38209 6100
rect 37332 6060 37338 6072
rect 38197 6069 38209 6072
rect 38243 6069 38255 6103
rect 38197 6063 38255 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 9122 5896 9128 5908
rect 6503 5868 9128 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 15010 5760 15016 5772
rect 4724 5732 15016 5760
rect 4724 5701 4752 5732
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 32769 5763 32827 5769
rect 32769 5760 32781 5763
rect 17368 5732 32781 5760
rect 17368 5720 17374 5732
rect 32769 5729 32781 5732
rect 32815 5729 32827 5763
rect 32769 5723 32827 5729
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 6362 5692 6368 5704
rect 6323 5664 6368 5692
rect 4709 5655 4767 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 21174 5692 21180 5704
rect 21135 5664 21180 5692
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 23198 5652 23204 5704
rect 23256 5652 23262 5704
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24728 5664 24777 5692
rect 24728 5652 24734 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 30377 5695 30435 5701
rect 30377 5661 30389 5695
rect 30423 5692 30435 5695
rect 32582 5692 32588 5704
rect 30423 5664 32588 5692
rect 30423 5661 30435 5664
rect 30377 5655 30435 5661
rect 32582 5652 32588 5664
rect 32640 5652 32646 5704
rect 32677 5695 32735 5701
rect 32677 5661 32689 5695
rect 32723 5692 32735 5695
rect 34514 5692 34520 5704
rect 32723 5664 34520 5692
rect 32723 5661 32735 5664
rect 32677 5655 32735 5661
rect 34514 5652 34520 5664
rect 34572 5652 34578 5704
rect 37090 5692 37096 5704
rect 37051 5664 37096 5692
rect 37090 5652 37096 5664
rect 37148 5652 37154 5704
rect 23216 5624 23244 5652
rect 30469 5627 30527 5633
rect 30469 5624 30481 5627
rect 23216 5596 30481 5624
rect 30469 5593 30481 5596
rect 30515 5593 30527 5627
rect 30469 5587 30527 5593
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9180 5528 9505 5556
rect 9180 5516 9186 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 19426 5556 19432 5568
rect 18187 5528 19432 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 19426 5516 19432 5528
rect 19484 5516 19490 5568
rect 20993 5559 21051 5565
rect 20993 5525 21005 5559
rect 21039 5556 21051 5559
rect 23198 5556 23204 5568
rect 21039 5528 23204 5556
rect 21039 5525 21051 5528
rect 20993 5519 21051 5525
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 24581 5559 24639 5565
rect 24581 5525 24593 5559
rect 24627 5556 24639 5559
rect 25866 5556 25872 5568
rect 24627 5528 25872 5556
rect 24627 5525 24639 5528
rect 24581 5519 24639 5525
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 36909 5559 36967 5565
rect 36909 5525 36921 5559
rect 36955 5556 36967 5559
rect 37826 5556 37832 5568
rect 36955 5528 37832 5556
rect 36955 5525 36967 5528
rect 36909 5519 36967 5525
rect 37826 5516 37832 5528
rect 37884 5516 37890 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1854 5284 1860 5296
rect 1815 5256 1860 5284
rect 1854 5244 1860 5256
rect 1912 5244 1918 5296
rect 1670 5216 1676 5228
rect 1631 5188 1676 5216
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 11882 5216 11888 5228
rect 11843 5188 11888 5216
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 15286 5216 15292 5228
rect 15247 5188 15292 5216
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5216 17831 5219
rect 18690 5216 18696 5228
rect 17819 5188 18696 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 18690 5176 18696 5188
rect 18748 5176 18754 5228
rect 20254 5216 20260 5228
rect 20215 5188 20260 5216
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 25590 5176 25596 5228
rect 25648 5216 25654 5228
rect 27893 5219 27951 5225
rect 27893 5216 27905 5219
rect 25648 5188 27905 5216
rect 25648 5176 25654 5188
rect 27893 5185 27905 5188
rect 27939 5185 27951 5219
rect 27893 5179 27951 5185
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 4672 4984 5733 5012
rect 4672 4972 4678 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 5721 4975 5779 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14976 4984 15117 5012
rect 14976 4972 14982 4984
rect 15105 4981 15117 4984
rect 15151 4981 15163 5015
rect 15105 4975 15163 4981
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 16908 4984 17601 5012
rect 16908 4972 16914 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 17589 4975 17647 4981
rect 20073 5015 20131 5021
rect 20073 4981 20085 5015
rect 20119 5012 20131 5015
rect 22646 5012 22652 5024
rect 20119 4984 22652 5012
rect 20119 4981 20131 4984
rect 20073 4975 20131 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 27709 5015 27767 5021
rect 27709 4981 27721 5015
rect 27755 5012 27767 5015
rect 31662 5012 31668 5024
rect 27755 4984 31668 5012
rect 27755 4981 27767 4984
rect 27709 4975 27767 4981
rect 31662 4972 31668 4984
rect 31720 4972 31726 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 37918 4768 37924 4820
rect 37976 4808 37982 4820
rect 38105 4811 38163 4817
rect 38105 4808 38117 4811
rect 37976 4780 38117 4808
rect 37976 4768 37982 4780
rect 38105 4777 38117 4780
rect 38151 4777 38163 4811
rect 38105 4771 38163 4777
rect 28350 4564 28356 4616
rect 28408 4604 28414 4616
rect 31665 4607 31723 4613
rect 31665 4604 31677 4607
rect 28408 4576 31677 4604
rect 28408 4564 28414 4576
rect 31665 4573 31677 4576
rect 31711 4573 31723 4607
rect 38286 4604 38292 4616
rect 38247 4576 38292 4604
rect 31665 4567 31723 4573
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 31481 4471 31539 4477
rect 31481 4437 31493 4471
rect 31527 4468 31539 4471
rect 33962 4468 33968 4480
rect 31527 4440 33968 4468
rect 31527 4437 31539 4440
rect 31481 4431 31539 4437
rect 33962 4428 33968 4440
rect 34020 4428 34026 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 4798 4128 4804 4140
rect 3375 4100 4804 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 35805 4131 35863 4137
rect 35805 4128 35817 4131
rect 23164 4100 35817 4128
rect 23164 4088 23170 4100
rect 35805 4097 35817 4100
rect 35851 4097 35863 4131
rect 35805 4091 35863 4097
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 35897 3927 35955 3933
rect 35897 3893 35909 3927
rect 35943 3924 35955 3927
rect 37458 3924 37464 3936
rect 35943 3896 37464 3924
rect 35943 3893 35955 3896
rect 35897 3887 35955 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 8294 3720 8300 3732
rect 1627 3692 8300 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 34514 3680 34520 3732
rect 34572 3720 34578 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 34572 3692 38117 3720
rect 34572 3680 34578 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 37458 3516 37464 3528
rect 37419 3488 37464 3516
rect 37458 3476 37464 3488
rect 37516 3476 37522 3528
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 38289 3519 38347 3525
rect 38289 3516 38301 3519
rect 38160 3488 38301 3516
rect 38160 3476 38166 3488
rect 38289 3485 38301 3488
rect 38335 3485 38347 3519
rect 38289 3479 38347 3485
rect 37277 3383 37335 3389
rect 37277 3349 37289 3383
rect 37323 3380 37335 3383
rect 38010 3380 38016 3392
rect 37323 3352 38016 3380
rect 37323 3349 37335 3352
rect 37277 3343 37335 3349
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3145 3111 3179
rect 3053 3139 3111 3145
rect 3068 3108 3096 3139
rect 35802 3136 35808 3188
rect 35860 3176 35866 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 35860 3148 36737 3176
rect 35860 3136 35866 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 1596 3080 3096 3108
rect 1596 3049 1624 3080
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 4614 3040 4620 3052
rect 3283 3012 4620 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 2516 2972 2544 3003
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 37826 3000 37832 3052
rect 37884 3040 37890 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37884 3012 38025 3040
rect 37884 3000 37890 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 1360 2944 2544 2972
rect 1360 2932 1366 2944
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 72 2808 1777 2836
rect 72 2796 78 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 1765 2799 1823 2805
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 6362 2632 6368 2644
rect 2731 2604 6368 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 9490 2632 9496 2644
rect 7239 2604 9496 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 11146 2632 11152 2644
rect 10459 2604 11152 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 24912 2604 27169 2632
rect 24912 2592 24918 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 30377 2635 30435 2641
rect 30377 2632 30389 2635
rect 28684 2604 30389 2632
rect 28684 2592 28690 2604
rect 30377 2601 30389 2604
rect 30423 2601 30435 2635
rect 30377 2595 30435 2601
rect 32582 2592 32588 2644
rect 32640 2632 32646 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 32640 2604 34897 2632
rect 32640 2592 32646 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 4617 2567 4675 2573
rect 4617 2533 4629 2567
rect 4663 2564 4675 2567
rect 4706 2564 4712 2576
rect 4663 2536 4712 2564
rect 4663 2533 4675 2536
rect 4617 2527 4675 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 26206 2536 29745 2564
rect 3142 2496 3148 2508
rect 1596 2468 3148 2496
rect 1596 2437 1624 2468
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 25406 2456 25412 2508
rect 25464 2496 25470 2508
rect 26206 2496 26234 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 30282 2524 30288 2576
rect 30340 2564 30346 2576
rect 33597 2567 33655 2573
rect 33597 2564 33609 2567
rect 30340 2536 33609 2564
rect 30340 2524 30346 2536
rect 33597 2533 33609 2536
rect 33643 2533 33655 2567
rect 33597 2527 33655 2533
rect 25464 2468 26234 2496
rect 25464 2456 25470 2468
rect 33962 2456 33968 2508
rect 34020 2496 34026 2508
rect 34020 2468 35894 2496
rect 34020 2456 34026 2468
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2648 2400 2881 2428
rect 2648 2388 2654 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 5868 2400 6745 2428
rect 5868 2388 5874 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 7377 2391 7435 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 11698 2428 11704 2440
rect 11659 2400 11704 2428
rect 10597 2391 10655 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13596 2400 14473 2428
rect 13596 2388 13602 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 14461 2391 14519 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 18325 2391 18383 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 22189 2391 22247 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23256 2400 24593 2428
rect 23256 2388 23262 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 25866 2428 25872 2440
rect 25827 2400 25872 2428
rect 24581 2391 24639 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30340 2400 30573 2428
rect 30340 2388 30346 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 31662 2388 31668 2440
rect 31720 2428 31726 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31720 2400 32321 2428
rect 31720 2388 31726 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 33560 2400 33793 2428
rect 33560 2388 33566 2400
rect 33781 2397 33793 2400
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34848 2400 35081 2428
rect 34848 2388 34854 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35866 2428 35894 2468
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35866 2400 36185 2428
rect 35069 2391 35127 2397
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 38010 2428 38016 2440
rect 37971 2400 38016 2428
rect 36173 2391 36231 2397
rect 38010 2388 38016 2400
rect 38068 2388 38074 2440
rect 13170 2360 13176 2372
rect 6886 2332 13176 2360
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 6886 2292 6914 2332
rect 13170 2320 13176 2332
rect 13228 2320 13234 2372
rect 6595 2264 6914 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 23900 2264 24777 2292
rect 23900 2252 23906 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 31628 2264 32505 2292
rect 31628 2252 31634 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 38197 2295 38255 2301
rect 38197 2261 38209 2295
rect 38243 2292 38255 2295
rect 39298 2292 39304 2304
rect 38243 2264 39304 2292
rect 38243 2261 38255 2264
rect 38197 2255 38255 2261
rect 39298 2252 39304 2264
rect 39356 2252 39362 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 5908 37748 5960 37800
rect 11060 37748 11112 37800
rect 4528 37680 4580 37732
rect 6552 37680 6604 37732
rect 7012 37680 7064 37732
rect 13268 37680 13320 37732
rect 4068 37612 4120 37664
rect 19340 37612 19392 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5908 37408 5960 37460
rect 6000 37408 6052 37460
rect 11060 37451 11112 37460
rect 4712 37272 4764 37324
rect 7012 37315 7064 37324
rect 7012 37281 7021 37315
rect 7021 37281 7055 37315
rect 7055 37281 7064 37315
rect 7012 37272 7064 37281
rect 9956 37272 10008 37324
rect 11060 37417 11069 37451
rect 11069 37417 11103 37451
rect 11103 37417 11112 37451
rect 11060 37408 11112 37417
rect 13912 37408 13964 37460
rect 20 37204 72 37256
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 3976 37247 4028 37256
rect 3148 37136 3200 37188
rect 1584 37068 1636 37120
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 6736 37247 6788 37256
rect 6736 37213 6745 37247
rect 6745 37213 6779 37247
rect 6779 37213 6788 37247
rect 6736 37204 6788 37213
rect 9128 37204 9180 37256
rect 11060 37204 11112 37256
rect 15108 37204 15160 37256
rect 15752 37204 15804 37256
rect 16672 37204 16724 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18052 37204 18104 37256
rect 19248 37204 19300 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 21272 37204 21324 37256
rect 22560 37204 22612 37256
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25780 37204 25832 37256
rect 27712 37204 27764 37256
rect 29000 37204 29052 37256
rect 30380 37204 30432 37256
rect 32220 37204 32272 37256
rect 33508 37204 33560 37256
rect 34796 37204 34848 37256
rect 36728 37204 36780 37256
rect 37280 37204 37332 37256
rect 4804 37136 4856 37188
rect 3424 37068 3476 37120
rect 5724 37111 5776 37120
rect 5724 37077 5733 37111
rect 5733 37077 5767 37111
rect 5767 37077 5776 37111
rect 5724 37068 5776 37077
rect 8484 37111 8536 37120
rect 8484 37077 8493 37111
rect 8493 37077 8527 37111
rect 8527 37077 8536 37111
rect 8484 37068 8536 37077
rect 10600 37136 10652 37188
rect 12348 37068 12400 37120
rect 12624 37068 12676 37120
rect 15844 37136 15896 37188
rect 20628 37136 20680 37188
rect 13360 37068 13412 37120
rect 13544 37068 13596 37120
rect 15476 37068 15528 37120
rect 16764 37068 16816 37120
rect 18144 37111 18196 37120
rect 18144 37077 18153 37111
rect 18153 37077 18187 37111
rect 18187 37077 18196 37111
rect 18144 37068 18196 37077
rect 19432 37111 19484 37120
rect 19432 37077 19441 37111
rect 19441 37077 19475 37111
rect 19475 37077 19484 37111
rect 19432 37068 19484 37077
rect 19984 37068 20036 37120
rect 20352 37068 20404 37120
rect 23940 37136 23992 37188
rect 24492 37068 24544 37120
rect 31484 37136 31536 37188
rect 27804 37111 27856 37120
rect 27804 37077 27813 37111
rect 27813 37077 27847 37111
rect 27847 37077 27856 37111
rect 27804 37068 27856 37077
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 30380 37111 30432 37120
rect 30380 37077 30389 37111
rect 30389 37077 30423 37111
rect 30423 37077 30432 37111
rect 30380 37068 30432 37077
rect 30656 37068 30708 37120
rect 32404 37068 32456 37120
rect 34520 37068 34572 37120
rect 38200 37111 38252 37120
rect 38200 37077 38209 37111
rect 38209 37077 38243 37111
rect 38243 37077 38252 37111
rect 38200 37068 38252 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 7380 36864 7432 36916
rect 4436 36796 4488 36848
rect 12348 36864 12400 36916
rect 12532 36864 12584 36916
rect 16212 36864 16264 36916
rect 24676 36864 24728 36916
rect 27804 36864 27856 36916
rect 1584 36771 1636 36780
rect 1584 36737 1593 36771
rect 1593 36737 1627 36771
rect 1627 36737 1636 36771
rect 1584 36728 1636 36737
rect 3976 36728 4028 36780
rect 8668 36796 8720 36848
rect 9680 36796 9732 36848
rect 10048 36796 10100 36848
rect 3240 36660 3292 36712
rect 3608 36703 3660 36712
rect 3608 36669 3617 36703
rect 3617 36669 3651 36703
rect 3651 36669 3660 36703
rect 3608 36660 3660 36669
rect 6736 36660 6788 36712
rect 7288 36703 7340 36712
rect 7288 36669 7297 36703
rect 7297 36669 7331 36703
rect 7331 36669 7340 36703
rect 7288 36660 7340 36669
rect 7380 36660 7432 36712
rect 8024 36660 8076 36712
rect 6920 36592 6972 36644
rect 8760 36703 8812 36712
rect 8760 36669 8769 36703
rect 8769 36669 8803 36703
rect 8803 36669 8812 36703
rect 8760 36660 8812 36669
rect 9128 36660 9180 36712
rect 9588 36703 9640 36712
rect 8576 36592 8628 36644
rect 9588 36669 9597 36703
rect 9597 36669 9631 36703
rect 9631 36669 9640 36703
rect 9588 36660 9640 36669
rect 9680 36660 9732 36712
rect 12164 36796 12216 36848
rect 12624 36796 12676 36848
rect 13728 36796 13780 36848
rect 15568 36728 15620 36780
rect 15844 36728 15896 36780
rect 17500 36771 17552 36780
rect 17500 36737 17509 36771
rect 17509 36737 17543 36771
rect 17543 36737 17552 36771
rect 17500 36728 17552 36737
rect 19340 36728 19392 36780
rect 39304 36796 39356 36848
rect 38016 36728 38068 36780
rect 11060 36660 11112 36712
rect 11796 36592 11848 36644
rect 11152 36524 11204 36576
rect 13360 36660 13412 36712
rect 14188 36703 14240 36712
rect 14188 36669 14197 36703
rect 14197 36669 14231 36703
rect 14231 36669 14240 36703
rect 14188 36660 14240 36669
rect 15660 36660 15712 36712
rect 15476 36592 15528 36644
rect 35900 36592 35952 36644
rect 13636 36567 13688 36576
rect 13636 36533 13645 36567
rect 13645 36533 13679 36567
rect 13679 36533 13688 36567
rect 13636 36524 13688 36533
rect 14280 36524 14332 36576
rect 16764 36524 16816 36576
rect 17592 36567 17644 36576
rect 17592 36533 17601 36567
rect 17601 36533 17635 36567
rect 17635 36533 17644 36567
rect 17592 36524 17644 36533
rect 19340 36524 19392 36576
rect 35992 36524 36044 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1584 36227 1636 36236
rect 1584 36193 1593 36227
rect 1593 36193 1627 36227
rect 1627 36193 1636 36227
rect 1584 36184 1636 36193
rect 5724 36320 5776 36372
rect 8300 36320 8352 36372
rect 9128 36252 9180 36304
rect 10324 36320 10376 36372
rect 3976 36184 4028 36236
rect 6736 36227 6788 36236
rect 6736 36193 6745 36227
rect 6745 36193 6779 36227
rect 6779 36193 6788 36227
rect 6736 36184 6788 36193
rect 7012 36184 7064 36236
rect 7564 36184 7616 36236
rect 7748 36184 7800 36236
rect 8208 36184 8260 36236
rect 8300 36184 8352 36236
rect 8392 36116 8444 36168
rect 8852 36184 8904 36236
rect 11060 36184 11112 36236
rect 12072 36320 12124 36372
rect 15476 36320 15528 36372
rect 15752 36363 15804 36372
rect 15752 36329 15761 36363
rect 15761 36329 15795 36363
rect 15795 36329 15804 36363
rect 15752 36320 15804 36329
rect 16764 36320 16816 36372
rect 12164 36252 12216 36304
rect 14280 36252 14332 36304
rect 16856 36252 16908 36304
rect 17592 36184 17644 36236
rect 9864 36116 9916 36168
rect 3884 36048 3936 36100
rect 4620 36048 4672 36100
rect 4988 36048 5040 36100
rect 4896 35980 4948 36032
rect 7012 36091 7064 36100
rect 7012 36057 7021 36091
rect 7021 36057 7055 36091
rect 7055 36057 7064 36091
rect 7012 36048 7064 36057
rect 8300 36048 8352 36100
rect 9220 35980 9272 36032
rect 12440 36116 12492 36168
rect 10968 36091 11020 36100
rect 10968 36057 10977 36091
rect 10977 36057 11011 36091
rect 11011 36057 11020 36091
rect 10968 36048 11020 36057
rect 11428 36048 11480 36100
rect 12992 36048 13044 36100
rect 12440 36023 12492 36032
rect 12440 35989 12449 36023
rect 12449 35989 12483 36023
rect 12483 35989 12492 36023
rect 12440 35980 12492 35989
rect 12624 35980 12676 36032
rect 13636 36116 13688 36168
rect 14648 36159 14700 36168
rect 14648 36125 14657 36159
rect 14657 36125 14691 36159
rect 14691 36125 14700 36159
rect 14648 36116 14700 36125
rect 15844 36116 15896 36168
rect 16580 36159 16632 36168
rect 14740 36048 14792 36100
rect 16580 36125 16589 36159
rect 16589 36125 16623 36159
rect 16623 36125 16632 36159
rect 16580 36116 16632 36125
rect 17500 36159 17552 36168
rect 17500 36125 17509 36159
rect 17509 36125 17543 36159
rect 17543 36125 17552 36159
rect 17500 36116 17552 36125
rect 37188 36116 37240 36168
rect 17132 36091 17184 36100
rect 17132 36057 17141 36091
rect 17141 36057 17175 36091
rect 17175 36057 17184 36091
rect 17132 36048 17184 36057
rect 13544 35980 13596 36032
rect 15384 35980 15436 36032
rect 16304 35980 16356 36032
rect 17592 36023 17644 36032
rect 17592 35989 17601 36023
rect 17601 35989 17635 36023
rect 17635 35989 17644 36023
rect 17592 35980 17644 35989
rect 18420 35980 18472 36032
rect 36084 35980 36136 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5816 35776 5868 35828
rect 12256 35776 12308 35828
rect 1952 35640 2004 35692
rect 10692 35708 10744 35760
rect 14740 35776 14792 35828
rect 15108 35776 15160 35828
rect 15292 35776 15344 35828
rect 17132 35776 17184 35828
rect 2964 35572 3016 35624
rect 3332 35615 3384 35624
rect 1584 35504 1636 35556
rect 3332 35581 3341 35615
rect 3341 35581 3375 35615
rect 3375 35581 3384 35615
rect 3332 35572 3384 35581
rect 6736 35640 6788 35692
rect 5908 35572 5960 35624
rect 6184 35572 6236 35624
rect 7840 35572 7892 35624
rect 8576 35615 8628 35624
rect 8576 35581 8585 35615
rect 8585 35581 8619 35615
rect 8619 35581 8628 35615
rect 8576 35572 8628 35581
rect 9128 35615 9180 35624
rect 9128 35581 9137 35615
rect 9137 35581 9171 35615
rect 9171 35581 9180 35615
rect 9128 35572 9180 35581
rect 10416 35572 10468 35624
rect 3516 35436 3568 35488
rect 4712 35436 4764 35488
rect 5080 35436 5132 35488
rect 8392 35436 8444 35488
rect 17592 35708 17644 35760
rect 11060 35572 11112 35624
rect 10968 35504 11020 35556
rect 12072 35572 12124 35624
rect 14464 35640 14516 35692
rect 14924 35640 14976 35692
rect 15384 35683 15436 35692
rect 15384 35649 15393 35683
rect 15393 35649 15427 35683
rect 15427 35649 15436 35683
rect 15384 35640 15436 35649
rect 15476 35640 15528 35692
rect 16488 35640 16540 35692
rect 17500 35683 17552 35692
rect 17500 35649 17509 35683
rect 17509 35649 17543 35683
rect 17543 35649 17552 35683
rect 17500 35640 17552 35649
rect 18236 35572 18288 35624
rect 12992 35504 13044 35556
rect 10876 35479 10928 35488
rect 10876 35445 10885 35479
rect 10885 35445 10919 35479
rect 10919 35445 10928 35479
rect 10876 35436 10928 35445
rect 11152 35436 11204 35488
rect 16580 35504 16632 35556
rect 14556 35436 14608 35488
rect 15108 35436 15160 35488
rect 15936 35479 15988 35488
rect 15936 35445 15945 35479
rect 15945 35445 15979 35479
rect 15979 35445 15988 35479
rect 15936 35436 15988 35445
rect 16948 35479 17000 35488
rect 16948 35445 16957 35479
rect 16957 35445 16991 35479
rect 16991 35445 17000 35479
rect 16948 35436 17000 35445
rect 17592 35479 17644 35488
rect 17592 35445 17601 35479
rect 17601 35445 17635 35479
rect 17635 35445 17644 35479
rect 17592 35436 17644 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6368 35232 6420 35284
rect 6644 35232 6696 35284
rect 6184 35207 6236 35216
rect 6184 35173 6193 35207
rect 6193 35173 6227 35207
rect 6227 35173 6236 35207
rect 6184 35164 6236 35173
rect 1584 35139 1636 35148
rect 1584 35105 1593 35139
rect 1593 35105 1627 35139
rect 1627 35105 1636 35139
rect 1584 35096 1636 35105
rect 3240 35096 3292 35148
rect 3424 35096 3476 35148
rect 3976 35096 4028 35148
rect 9128 35139 9180 35148
rect 9128 35105 9137 35139
rect 9137 35105 9171 35139
rect 9171 35105 9180 35139
rect 9128 35096 9180 35105
rect 9404 35139 9456 35148
rect 9404 35105 9413 35139
rect 9413 35105 9447 35139
rect 9447 35105 9456 35139
rect 9404 35096 9456 35105
rect 11520 35232 11572 35284
rect 15936 35232 15988 35284
rect 24584 35232 24636 35284
rect 12808 35164 12860 35216
rect 14096 35096 14148 35148
rect 14188 35096 14240 35148
rect 20076 35164 20128 35216
rect 17868 35096 17920 35148
rect 8024 35028 8076 35080
rect 10508 35028 10560 35080
rect 11060 35028 11112 35080
rect 16120 35028 16172 35080
rect 16396 35028 16448 35080
rect 17684 35028 17736 35080
rect 22928 35071 22980 35080
rect 22928 35037 22937 35071
rect 22937 35037 22971 35071
rect 22971 35037 22980 35071
rect 22928 35028 22980 35037
rect 34244 35028 34296 35080
rect 3332 34935 3384 34944
rect 3332 34901 3341 34935
rect 3341 34901 3375 34935
rect 3375 34901 3384 34935
rect 3332 34892 3384 34901
rect 6092 34892 6144 34944
rect 6920 35003 6972 35012
rect 6920 34969 6929 35003
rect 6929 34969 6963 35003
rect 6963 34969 6972 35003
rect 6920 34960 6972 34969
rect 8392 34935 8444 34944
rect 8392 34901 8401 34935
rect 8401 34901 8435 34935
rect 8435 34901 8444 34935
rect 8392 34892 8444 34901
rect 10784 34892 10836 34944
rect 11152 34960 11204 35012
rect 12532 34960 12584 35012
rect 14556 35003 14608 35012
rect 14556 34969 14565 35003
rect 14565 34969 14599 35003
rect 14599 34969 14608 35003
rect 14556 34960 14608 34969
rect 13176 34892 13228 34944
rect 13268 34935 13320 34944
rect 13268 34901 13277 34935
rect 13277 34901 13311 34935
rect 13311 34901 13320 34935
rect 13268 34892 13320 34901
rect 13452 34892 13504 34944
rect 15936 34892 15988 34944
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2688 34688 2740 34740
rect 14004 34688 14056 34740
rect 14096 34688 14148 34740
rect 15016 34688 15068 34740
rect 17500 34688 17552 34740
rect 18236 34731 18288 34740
rect 18236 34697 18245 34731
rect 18245 34697 18279 34731
rect 18279 34697 18288 34731
rect 18236 34688 18288 34697
rect 4712 34620 4764 34672
rect 1952 34552 2004 34604
rect 2688 34552 2740 34604
rect 3976 34552 4028 34604
rect 5540 34552 5592 34604
rect 3056 34527 3108 34536
rect 3056 34493 3065 34527
rect 3065 34493 3099 34527
rect 3099 34493 3108 34527
rect 3056 34484 3108 34493
rect 7656 34620 7708 34672
rect 12072 34620 12124 34672
rect 16948 34620 17000 34672
rect 7196 34552 7248 34604
rect 6828 34484 6880 34536
rect 6552 34416 6604 34468
rect 4896 34348 4948 34400
rect 5172 34348 5224 34400
rect 6368 34348 6420 34400
rect 8116 34484 8168 34536
rect 9128 34484 9180 34536
rect 10508 34552 10560 34604
rect 11060 34552 11112 34604
rect 10876 34527 10928 34536
rect 10876 34493 10885 34527
rect 10885 34493 10919 34527
rect 10919 34493 10928 34527
rect 10876 34484 10928 34493
rect 11336 34484 11388 34536
rect 11980 34527 12032 34536
rect 11980 34493 11989 34527
rect 11989 34493 12023 34527
rect 12023 34493 12032 34527
rect 11980 34484 12032 34493
rect 12072 34484 12124 34536
rect 12440 34484 12492 34536
rect 12532 34484 12584 34536
rect 13728 34484 13780 34536
rect 14740 34595 14792 34604
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 15292 34552 15344 34604
rect 15476 34595 15528 34604
rect 15476 34561 15485 34595
rect 15485 34561 15519 34595
rect 15519 34561 15528 34595
rect 15476 34552 15528 34561
rect 16396 34552 16448 34604
rect 11244 34416 11296 34468
rect 16212 34484 16264 34536
rect 16948 34527 17000 34536
rect 16948 34493 16957 34527
rect 16957 34493 16991 34527
rect 16991 34493 17000 34527
rect 16948 34484 17000 34493
rect 16488 34416 16540 34468
rect 18604 34552 18656 34604
rect 9588 34391 9640 34400
rect 9588 34357 9597 34391
rect 9597 34357 9631 34391
rect 9631 34357 9640 34391
rect 10140 34391 10192 34400
rect 9588 34348 9640 34357
rect 10140 34357 10149 34391
rect 10149 34357 10183 34391
rect 10183 34357 10192 34391
rect 10140 34348 10192 34357
rect 12348 34348 12400 34400
rect 14096 34348 14148 34400
rect 14372 34348 14424 34400
rect 15108 34348 15160 34400
rect 16856 34348 16908 34400
rect 17592 34391 17644 34400
rect 17592 34357 17601 34391
rect 17601 34357 17635 34391
rect 17635 34357 17644 34391
rect 17592 34348 17644 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6736 34144 6788 34196
rect 10784 34144 10836 34196
rect 8116 34076 8168 34128
rect 3976 34051 4028 34060
rect 3976 34017 3985 34051
rect 3985 34017 4019 34051
rect 4019 34017 4028 34051
rect 3976 34008 4028 34017
rect 4712 34008 4764 34060
rect 6000 34051 6052 34060
rect 1952 33940 2004 33992
rect 3240 33940 3292 33992
rect 6000 34017 6009 34051
rect 6009 34017 6043 34051
rect 6043 34017 6052 34051
rect 6000 34008 6052 34017
rect 6368 34008 6420 34060
rect 11152 34076 11204 34128
rect 9772 34008 9824 34060
rect 10048 34008 10100 34060
rect 10968 34008 11020 34060
rect 11060 34008 11112 34060
rect 13268 34144 13320 34196
rect 13544 34144 13596 34196
rect 15108 34144 15160 34196
rect 12348 34008 12400 34060
rect 14372 34051 14424 34060
rect 14372 34017 14381 34051
rect 14381 34017 14415 34051
rect 14415 34017 14424 34051
rect 14372 34008 14424 34017
rect 15844 34076 15896 34128
rect 16488 34076 16540 34128
rect 17868 34144 17920 34196
rect 37280 34144 37332 34196
rect 19156 34076 19208 34128
rect 6552 33940 6604 33992
rect 6828 33983 6880 33992
rect 6828 33949 6837 33983
rect 6837 33949 6871 33983
rect 6871 33949 6880 33983
rect 6828 33940 6880 33949
rect 8208 33940 8260 33992
rect 10784 33940 10836 33992
rect 13176 33940 13228 33992
rect 1400 33872 1452 33924
rect 4160 33872 4212 33924
rect 6644 33872 6696 33924
rect 8484 33872 8536 33924
rect 9036 33872 9088 33924
rect 11888 33872 11940 33924
rect 13452 33872 13504 33924
rect 14004 33872 14056 33924
rect 12716 33804 12768 33856
rect 19248 34008 19300 34060
rect 16028 33940 16080 33992
rect 17316 33983 17368 33992
rect 17316 33949 17325 33983
rect 17325 33949 17359 33983
rect 17359 33949 17368 33983
rect 17316 33940 17368 33949
rect 18604 33983 18656 33992
rect 16212 33915 16264 33924
rect 16212 33881 16221 33915
rect 16221 33881 16255 33915
rect 16255 33881 16264 33915
rect 16212 33872 16264 33881
rect 16396 33872 16448 33924
rect 18604 33949 18613 33983
rect 18613 33949 18647 33983
rect 18647 33949 18656 33983
rect 18604 33940 18656 33949
rect 34520 33940 34572 33992
rect 17868 33804 17920 33856
rect 18696 33847 18748 33856
rect 18696 33813 18705 33847
rect 18705 33813 18739 33847
rect 18739 33813 18748 33847
rect 18696 33804 18748 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 2136 33600 2188 33652
rect 2320 33575 2372 33584
rect 2320 33541 2329 33575
rect 2329 33541 2363 33575
rect 2363 33541 2372 33575
rect 2320 33532 2372 33541
rect 5448 33600 5500 33652
rect 6920 33600 6972 33652
rect 7748 33600 7800 33652
rect 7840 33600 7892 33652
rect 9404 33600 9456 33652
rect 1584 33464 1636 33516
rect 3976 33464 4028 33516
rect 6552 33507 6604 33516
rect 4528 33439 4580 33448
rect 4528 33405 4537 33439
rect 4537 33405 4571 33439
rect 4571 33405 4580 33439
rect 4528 33396 4580 33405
rect 6552 33473 6561 33507
rect 6561 33473 6595 33507
rect 6595 33473 6604 33507
rect 6552 33464 6604 33473
rect 7104 33464 7156 33516
rect 7380 33464 7432 33516
rect 11520 33600 11572 33652
rect 12624 33600 12676 33652
rect 14004 33643 14056 33652
rect 10048 33532 10100 33584
rect 14004 33609 14013 33643
rect 14013 33609 14047 33643
rect 14047 33609 14056 33643
rect 14004 33600 14056 33609
rect 14096 33600 14148 33652
rect 15844 33600 15896 33652
rect 16028 33643 16080 33652
rect 16028 33609 16037 33643
rect 16037 33609 16071 33643
rect 16071 33609 16080 33643
rect 16028 33600 16080 33609
rect 16212 33600 16264 33652
rect 10416 33464 10468 33516
rect 10968 33507 11020 33516
rect 10968 33473 10977 33507
rect 10977 33473 11011 33507
rect 11011 33473 11020 33507
rect 10968 33464 11020 33473
rect 11060 33464 11112 33516
rect 13912 33507 13964 33516
rect 6828 33396 6880 33448
rect 9312 33396 9364 33448
rect 9404 33396 9456 33448
rect 11520 33396 11572 33448
rect 5540 33260 5592 33312
rect 6736 33260 6788 33312
rect 11152 33328 11204 33380
rect 12072 33396 12124 33448
rect 12716 33396 12768 33448
rect 12992 33396 13044 33448
rect 13912 33473 13921 33507
rect 13921 33473 13955 33507
rect 13955 33473 13964 33507
rect 13912 33464 13964 33473
rect 14004 33464 14056 33516
rect 14740 33464 14792 33516
rect 15200 33507 15252 33516
rect 15200 33473 15209 33507
rect 15209 33473 15243 33507
rect 15243 33473 15252 33507
rect 15200 33464 15252 33473
rect 17316 33532 17368 33584
rect 17868 33575 17920 33584
rect 17868 33541 17877 33575
rect 17877 33541 17911 33575
rect 17911 33541 17920 33575
rect 17868 33532 17920 33541
rect 20352 33464 20404 33516
rect 31484 33507 31536 33516
rect 31484 33473 31493 33507
rect 31493 33473 31527 33507
rect 31527 33473 31536 33507
rect 31484 33464 31536 33473
rect 37924 33464 37976 33516
rect 17592 33396 17644 33448
rect 19984 33396 20036 33448
rect 13544 33328 13596 33380
rect 15200 33328 15252 33380
rect 16212 33328 16264 33380
rect 16488 33328 16540 33380
rect 9772 33260 9824 33312
rect 10600 33260 10652 33312
rect 12072 33260 12124 33312
rect 14096 33260 14148 33312
rect 15844 33260 15896 33312
rect 21272 33328 21324 33380
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 20260 33303 20312 33312
rect 20260 33269 20269 33303
rect 20269 33269 20303 33303
rect 20303 33269 20312 33303
rect 20260 33260 20312 33269
rect 29000 33260 29052 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1768 33099 1820 33108
rect 1768 33065 1777 33099
rect 1777 33065 1811 33099
rect 1811 33065 1820 33099
rect 1768 33056 1820 33065
rect 3148 33056 3200 33108
rect 8944 33056 8996 33108
rect 13728 33056 13780 33108
rect 13820 33056 13872 33108
rect 18696 33056 18748 33108
rect 9588 32988 9640 33040
rect 9680 32988 9732 33040
rect 11152 32988 11204 33040
rect 2964 32920 3016 32972
rect 3332 32920 3384 32972
rect 1492 32852 1544 32904
rect 2320 32895 2372 32904
rect 2320 32861 2329 32895
rect 2329 32861 2363 32895
rect 2363 32861 2372 32895
rect 3148 32895 3200 32904
rect 2320 32852 2372 32861
rect 3148 32861 3157 32895
rect 3157 32861 3191 32895
rect 3191 32861 3200 32895
rect 3148 32852 3200 32861
rect 3240 32852 3292 32904
rect 4252 32852 4304 32904
rect 4988 32920 5040 32972
rect 4712 32852 4764 32904
rect 4896 32852 4948 32904
rect 5540 32920 5592 32972
rect 6552 32963 6604 32972
rect 6552 32929 6561 32963
rect 6561 32929 6595 32963
rect 6595 32929 6604 32963
rect 6552 32920 6604 32929
rect 6828 32920 6880 32972
rect 7380 32920 7432 32972
rect 6460 32784 6512 32836
rect 2412 32759 2464 32768
rect 2412 32725 2421 32759
rect 2421 32725 2455 32759
rect 2455 32725 2464 32759
rect 2412 32716 2464 32725
rect 3792 32716 3844 32768
rect 4712 32759 4764 32768
rect 4712 32725 4721 32759
rect 4721 32725 4755 32759
rect 4755 32725 4764 32759
rect 4712 32716 4764 32725
rect 5724 32716 5776 32768
rect 6092 32716 6144 32768
rect 8944 32852 8996 32904
rect 9220 32920 9272 32972
rect 9404 32852 9456 32904
rect 9956 32852 10008 32904
rect 10416 32895 10468 32904
rect 10416 32861 10425 32895
rect 10425 32861 10459 32895
rect 10459 32861 10468 32895
rect 10416 32852 10468 32861
rect 8484 32784 8536 32836
rect 7472 32716 7524 32768
rect 8116 32716 8168 32768
rect 11060 32920 11112 32972
rect 11520 32920 11572 32972
rect 15476 32988 15528 33040
rect 16672 32988 16724 33040
rect 21088 32988 21140 33040
rect 16948 32920 17000 32972
rect 14004 32852 14056 32904
rect 15016 32895 15068 32904
rect 9220 32759 9272 32768
rect 9220 32725 9229 32759
rect 9229 32725 9263 32759
rect 9263 32725 9272 32759
rect 9220 32716 9272 32725
rect 9404 32716 9456 32768
rect 10232 32716 10284 32768
rect 13268 32716 13320 32768
rect 13912 32784 13964 32836
rect 15016 32861 15025 32895
rect 15025 32861 15059 32895
rect 15059 32861 15068 32895
rect 15016 32852 15068 32861
rect 14832 32784 14884 32836
rect 15936 32784 15988 32836
rect 16488 32852 16540 32904
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 19248 32852 19300 32904
rect 18144 32784 18196 32836
rect 29736 32852 29788 32904
rect 35900 32852 35952 32904
rect 14372 32759 14424 32768
rect 14372 32725 14381 32759
rect 14381 32725 14415 32759
rect 14415 32725 14424 32759
rect 14372 32716 14424 32725
rect 14464 32716 14516 32768
rect 16028 32716 16080 32768
rect 16948 32759 17000 32768
rect 16948 32725 16957 32759
rect 16957 32725 16991 32759
rect 16991 32725 17000 32759
rect 16948 32716 17000 32725
rect 22192 32716 22244 32768
rect 22560 32716 22612 32768
rect 31760 32716 31812 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4252 32512 4304 32564
rect 2872 32444 2924 32496
rect 4804 32444 4856 32496
rect 4988 32419 5040 32428
rect 4988 32385 4997 32419
rect 4997 32385 5031 32419
rect 5031 32385 5040 32419
rect 4988 32376 5040 32385
rect 5816 32512 5868 32564
rect 6460 32512 6512 32564
rect 10600 32512 10652 32564
rect 10692 32512 10744 32564
rect 12164 32512 12216 32564
rect 7104 32444 7156 32496
rect 7656 32444 7708 32496
rect 11520 32444 11572 32496
rect 13820 32444 13872 32496
rect 6000 32376 6052 32428
rect 6828 32376 6880 32428
rect 9680 32376 9732 32428
rect 9956 32376 10008 32428
rect 10784 32376 10836 32428
rect 10968 32376 11020 32428
rect 11060 32376 11112 32428
rect 14004 32555 14056 32564
rect 14004 32521 14013 32555
rect 14013 32521 14047 32555
rect 14047 32521 14056 32555
rect 14004 32512 14056 32521
rect 14188 32512 14240 32564
rect 14464 32512 14516 32564
rect 14648 32512 14700 32564
rect 16212 32512 16264 32564
rect 16396 32512 16448 32564
rect 14372 32444 14424 32496
rect 1584 32308 1636 32360
rect 2688 32351 2740 32360
rect 2688 32317 2697 32351
rect 2697 32317 2731 32351
rect 2731 32317 2740 32351
rect 2688 32308 2740 32317
rect 5172 32240 5224 32292
rect 5632 32240 5684 32292
rect 5908 32240 5960 32292
rect 6644 32308 6696 32360
rect 8392 32308 8444 32360
rect 10600 32308 10652 32360
rect 15016 32376 15068 32428
rect 15384 32376 15436 32428
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 19524 32512 19576 32564
rect 20628 32512 20680 32564
rect 17776 32376 17828 32428
rect 22560 32419 22612 32428
rect 14372 32308 14424 32360
rect 6920 32240 6972 32292
rect 9036 32240 9088 32292
rect 9404 32240 9456 32292
rect 14188 32240 14240 32292
rect 18052 32308 18104 32360
rect 22560 32385 22569 32419
rect 22569 32385 22603 32419
rect 22603 32385 22612 32419
rect 22560 32376 22612 32385
rect 23940 32419 23992 32428
rect 23940 32385 23949 32419
rect 23949 32385 23983 32419
rect 23983 32385 23992 32419
rect 23940 32376 23992 32385
rect 2596 32172 2648 32224
rect 3516 32172 3568 32224
rect 9680 32172 9732 32224
rect 10232 32215 10284 32224
rect 10232 32181 10241 32215
rect 10241 32181 10275 32215
rect 10275 32181 10284 32215
rect 10232 32172 10284 32181
rect 10416 32172 10468 32224
rect 10784 32172 10836 32224
rect 11796 32172 11848 32224
rect 12532 32172 12584 32224
rect 12716 32172 12768 32224
rect 14556 32172 14608 32224
rect 14740 32172 14792 32224
rect 15200 32172 15252 32224
rect 15476 32240 15528 32292
rect 16488 32240 16540 32292
rect 18604 32240 18656 32292
rect 22744 32240 22796 32292
rect 26148 32240 26200 32292
rect 32220 32376 32272 32428
rect 34520 32444 34572 32496
rect 38292 32419 38344 32428
rect 38292 32385 38301 32419
rect 38301 32385 38335 32419
rect 38335 32385 38344 32419
rect 38292 32376 38344 32385
rect 35992 32308 36044 32360
rect 17500 32172 17552 32224
rect 18880 32172 18932 32224
rect 20352 32172 20404 32224
rect 22836 32215 22888 32224
rect 22836 32181 22845 32215
rect 22845 32181 22879 32215
rect 22879 32181 22888 32215
rect 22836 32172 22888 32181
rect 26332 32172 26384 32224
rect 32404 32215 32456 32224
rect 32404 32181 32413 32215
rect 32413 32181 32447 32215
rect 32447 32181 32456 32215
rect 32404 32172 32456 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3976 31968 4028 32020
rect 1584 31875 1636 31884
rect 1584 31841 1593 31875
rect 1593 31841 1627 31875
rect 1627 31841 1636 31875
rect 1584 31832 1636 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 5540 31968 5592 32020
rect 8116 31968 8168 32020
rect 15660 32011 15712 32020
rect 15660 31977 15669 32011
rect 15669 31977 15703 32011
rect 15703 31977 15712 32011
rect 15660 31968 15712 31977
rect 15936 31968 15988 32020
rect 16856 31968 16908 32020
rect 19984 31968 20036 32020
rect 22836 31968 22888 32020
rect 8576 31900 8628 31952
rect 9496 31900 9548 31952
rect 13636 31943 13688 31952
rect 13636 31909 13645 31943
rect 13645 31909 13679 31943
rect 13679 31909 13688 31943
rect 13636 31900 13688 31909
rect 20076 31900 20128 31952
rect 7288 31832 7340 31884
rect 7656 31832 7708 31884
rect 10692 31832 10744 31884
rect 11060 31832 11112 31884
rect 11704 31832 11756 31884
rect 14372 31875 14424 31884
rect 14372 31841 14381 31875
rect 14381 31841 14415 31875
rect 14415 31841 14424 31875
rect 14372 31832 14424 31841
rect 19340 31832 19392 31884
rect 21088 31900 21140 31952
rect 20536 31875 20588 31884
rect 3976 31807 4028 31816
rect 3976 31773 3985 31807
rect 3985 31773 4019 31807
rect 4019 31773 4028 31807
rect 3976 31764 4028 31773
rect 4804 31764 4856 31816
rect 6920 31807 6972 31816
rect 6920 31773 6929 31807
rect 6929 31773 6963 31807
rect 6963 31773 6972 31807
rect 6920 31764 6972 31773
rect 4620 31696 4672 31748
rect 6184 31696 6236 31748
rect 7380 31807 7432 31816
rect 7380 31773 7389 31807
rect 7389 31773 7423 31807
rect 7423 31773 7432 31807
rect 7380 31764 7432 31773
rect 8668 31764 8720 31816
rect 7472 31696 7524 31748
rect 7932 31696 7984 31748
rect 8852 31696 8904 31748
rect 9404 31696 9456 31748
rect 9864 31764 9916 31816
rect 10140 31764 10192 31816
rect 10416 31764 10468 31816
rect 13544 31807 13596 31816
rect 13544 31773 13553 31807
rect 13553 31773 13587 31807
rect 13587 31773 13596 31807
rect 13544 31764 13596 31773
rect 13820 31764 13872 31816
rect 14004 31764 14056 31816
rect 15016 31764 15068 31816
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 19524 31807 19576 31816
rect 19524 31773 19533 31807
rect 19533 31773 19567 31807
rect 19567 31773 19576 31807
rect 19524 31764 19576 31773
rect 10784 31696 10836 31748
rect 11612 31739 11664 31748
rect 11612 31705 11621 31739
rect 11621 31705 11655 31739
rect 11655 31705 11664 31739
rect 11612 31696 11664 31705
rect 12072 31696 12124 31748
rect 12992 31696 13044 31748
rect 20536 31841 20545 31875
rect 20545 31841 20579 31875
rect 20579 31841 20588 31875
rect 20536 31832 20588 31841
rect 22192 31875 22244 31884
rect 22192 31841 22201 31875
rect 22201 31841 22235 31875
rect 22235 31841 22244 31875
rect 22192 31832 22244 31841
rect 21824 31764 21876 31816
rect 32404 31832 32456 31884
rect 25136 31807 25188 31816
rect 25136 31773 25145 31807
rect 25145 31773 25179 31807
rect 25179 31773 25188 31807
rect 25136 31764 25188 31773
rect 25504 31764 25556 31816
rect 7104 31628 7156 31680
rect 10968 31628 11020 31680
rect 12624 31628 12676 31680
rect 20352 31739 20404 31748
rect 20352 31705 20361 31739
rect 20361 31705 20395 31739
rect 20395 31705 20404 31739
rect 20352 31696 20404 31705
rect 24860 31628 24912 31680
rect 25228 31671 25280 31680
rect 25228 31637 25237 31671
rect 25237 31637 25271 31671
rect 25271 31637 25280 31671
rect 25228 31628 25280 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1952 31467 2004 31476
rect 1952 31433 1961 31467
rect 1961 31433 1995 31467
rect 1995 31433 2004 31467
rect 1952 31424 2004 31433
rect 3056 31424 3108 31476
rect 4528 31356 4580 31408
rect 1860 31331 1912 31340
rect 1860 31297 1869 31331
rect 1869 31297 1903 31331
rect 1903 31297 1912 31331
rect 1860 31288 1912 31297
rect 2688 31331 2740 31340
rect 2688 31297 2697 31331
rect 2697 31297 2731 31331
rect 2731 31297 2740 31331
rect 2688 31288 2740 31297
rect 5632 31424 5684 31476
rect 6828 31424 6880 31476
rect 9128 31424 9180 31476
rect 9220 31424 9272 31476
rect 9404 31424 9456 31476
rect 10876 31424 10928 31476
rect 10968 31424 11020 31476
rect 13084 31424 13136 31476
rect 14280 31424 14332 31476
rect 17132 31424 17184 31476
rect 10784 31356 10836 31408
rect 19984 31424 20036 31476
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 5632 31331 5684 31340
rect 4988 31288 5040 31297
rect 5632 31297 5641 31331
rect 5641 31297 5675 31331
rect 5675 31297 5684 31331
rect 5632 31288 5684 31297
rect 5816 31288 5868 31340
rect 10968 31288 11020 31340
rect 11980 31288 12032 31340
rect 12532 31288 12584 31340
rect 5908 31220 5960 31272
rect 6552 31263 6604 31272
rect 6552 31229 6561 31263
rect 6561 31229 6595 31263
rect 6595 31229 6604 31263
rect 6552 31220 6604 31229
rect 6828 31263 6880 31272
rect 6828 31229 6837 31263
rect 6837 31229 6871 31263
rect 6871 31229 6880 31263
rect 6828 31220 6880 31229
rect 7196 31220 7248 31272
rect 4620 31084 4672 31136
rect 6920 31084 6972 31136
rect 8484 31084 8536 31136
rect 8760 31220 8812 31272
rect 9404 31263 9456 31272
rect 9404 31229 9413 31263
rect 9413 31229 9447 31263
rect 9447 31229 9456 31263
rect 9404 31220 9456 31229
rect 10600 31220 10652 31272
rect 12900 31220 12952 31272
rect 13452 31331 13504 31340
rect 13452 31297 13461 31331
rect 13461 31297 13495 31331
rect 13495 31297 13504 31331
rect 13452 31288 13504 31297
rect 13820 31220 13872 31272
rect 14280 31288 14332 31340
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 15384 31331 15436 31340
rect 15384 31297 15393 31331
rect 15393 31297 15427 31331
rect 15427 31297 15436 31331
rect 15384 31288 15436 31297
rect 16396 31288 16448 31340
rect 18604 31356 18656 31408
rect 20076 31399 20128 31408
rect 20076 31365 20085 31399
rect 20085 31365 20119 31399
rect 20119 31365 20128 31399
rect 20076 31356 20128 31365
rect 17960 31288 18012 31340
rect 18788 31263 18840 31272
rect 18788 31229 18797 31263
rect 18797 31229 18831 31263
rect 18831 31229 18840 31263
rect 18788 31220 18840 31229
rect 18972 31220 19024 31272
rect 12072 31152 12124 31204
rect 13636 31152 13688 31204
rect 19156 31152 19208 31204
rect 31760 31424 31812 31476
rect 25044 31331 25096 31340
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 25228 31288 25280 31340
rect 36084 31288 36136 31340
rect 29000 31220 29052 31272
rect 12900 31127 12952 31136
rect 12900 31093 12909 31127
rect 12909 31093 12943 31127
rect 12943 31093 12952 31127
rect 12900 31084 12952 31093
rect 13820 31084 13872 31136
rect 15292 31084 15344 31136
rect 19616 31084 19668 31136
rect 25320 31152 25372 31204
rect 20720 31084 20772 31136
rect 25596 31084 25648 31136
rect 32404 31127 32456 31136
rect 32404 31093 32413 31127
rect 32413 31093 32447 31127
rect 32447 31093 32456 31127
rect 32404 31084 32456 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4896 30880 4948 30932
rect 5356 30880 5408 30932
rect 5908 30880 5960 30932
rect 6276 30880 6328 30932
rect 6828 30880 6880 30932
rect 9588 30880 9640 30932
rect 11980 30923 12032 30932
rect 7380 30812 7432 30864
rect 11612 30812 11664 30864
rect 11980 30889 11989 30923
rect 11989 30889 12023 30923
rect 12023 30889 12032 30923
rect 11980 30880 12032 30889
rect 12440 30880 12492 30932
rect 13728 30880 13780 30932
rect 18788 30880 18840 30932
rect 21180 30880 21232 30932
rect 24860 30880 24912 30932
rect 26608 30880 26660 30932
rect 12992 30812 13044 30864
rect 15200 30812 15252 30864
rect 18236 30812 18288 30864
rect 2044 30744 2096 30796
rect 2320 30744 2372 30796
rect 4896 30744 4948 30796
rect 1860 30719 1912 30728
rect 1860 30685 1869 30719
rect 1869 30685 1903 30719
rect 1903 30685 1912 30719
rect 1860 30676 1912 30685
rect 2228 30676 2280 30728
rect 5632 30676 5684 30728
rect 6000 30719 6052 30728
rect 6000 30685 6009 30719
rect 6009 30685 6043 30719
rect 6043 30685 6052 30719
rect 6000 30676 6052 30685
rect 6644 30719 6696 30728
rect 6644 30685 6653 30719
rect 6653 30685 6687 30719
rect 6687 30685 6696 30719
rect 6644 30676 6696 30685
rect 6828 30676 6880 30728
rect 6092 30608 6144 30660
rect 2964 30540 3016 30592
rect 3884 30540 3936 30592
rect 4620 30540 4672 30592
rect 4988 30540 5040 30592
rect 7104 30540 7156 30592
rect 7196 30583 7248 30592
rect 7196 30549 7205 30583
rect 7205 30549 7239 30583
rect 7239 30549 7248 30583
rect 7196 30540 7248 30549
rect 9312 30719 9364 30728
rect 9312 30685 9321 30719
rect 9321 30685 9355 30719
rect 9355 30685 9364 30719
rect 9312 30676 9364 30685
rect 10232 30744 10284 30796
rect 11980 30744 12032 30796
rect 11060 30676 11112 30728
rect 11152 30676 11204 30728
rect 11888 30719 11940 30728
rect 11888 30685 11897 30719
rect 11897 30685 11931 30719
rect 11931 30685 11940 30719
rect 11888 30676 11940 30685
rect 19432 30744 19484 30796
rect 26148 30787 26200 30796
rect 26148 30753 26157 30787
rect 26157 30753 26191 30787
rect 26191 30753 26200 30787
rect 26148 30744 26200 30753
rect 12808 30676 12860 30728
rect 13084 30676 13136 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 14740 30676 14792 30728
rect 19616 30719 19668 30728
rect 10876 30608 10928 30660
rect 19616 30685 19625 30719
rect 19625 30685 19659 30719
rect 19659 30685 19668 30719
rect 19616 30676 19668 30685
rect 24676 30676 24728 30728
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26608 30676 26660 30685
rect 30656 30676 30708 30728
rect 18236 30651 18288 30660
rect 10416 30540 10468 30592
rect 10692 30540 10744 30592
rect 11520 30540 11572 30592
rect 12072 30540 12124 30592
rect 15384 30540 15436 30592
rect 18236 30617 18245 30651
rect 18245 30617 18279 30651
rect 18279 30617 18288 30651
rect 18236 30608 18288 30617
rect 18328 30651 18380 30660
rect 18328 30617 18337 30651
rect 18337 30617 18371 30651
rect 18371 30617 18380 30651
rect 18328 30608 18380 30617
rect 18972 30608 19024 30660
rect 25320 30608 25372 30660
rect 16304 30583 16356 30592
rect 16304 30549 16313 30583
rect 16313 30549 16347 30583
rect 16347 30549 16356 30583
rect 16304 30540 16356 30549
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6644 30336 6696 30388
rect 12348 30336 12400 30388
rect 13452 30311 13504 30320
rect 1584 30200 1636 30252
rect 3424 30132 3476 30184
rect 3976 30132 4028 30184
rect 5632 30200 5684 30252
rect 6276 30200 6328 30252
rect 5172 30132 5224 30184
rect 5908 30132 5960 30184
rect 6552 30132 6604 30184
rect 1952 29996 2004 30048
rect 5080 30039 5132 30048
rect 5080 30005 5089 30039
rect 5089 30005 5123 30039
rect 5123 30005 5132 30039
rect 5080 29996 5132 30005
rect 10232 30200 10284 30252
rect 8760 30132 8812 30184
rect 10784 30200 10836 30252
rect 10968 30200 11020 30252
rect 10508 30132 10560 30184
rect 12532 30200 12584 30252
rect 13452 30277 13461 30311
rect 13461 30277 13495 30311
rect 13495 30277 13504 30311
rect 13452 30268 13504 30277
rect 18328 30336 18380 30388
rect 17684 30311 17736 30320
rect 13820 30200 13872 30252
rect 14004 30200 14056 30252
rect 17684 30277 17693 30311
rect 17693 30277 17727 30311
rect 17727 30277 17736 30311
rect 17684 30268 17736 30277
rect 19432 30268 19484 30320
rect 25504 30311 25556 30320
rect 25504 30277 25513 30311
rect 25513 30277 25547 30311
rect 25547 30277 25556 30311
rect 25504 30268 25556 30277
rect 25596 30311 25648 30320
rect 25596 30277 25605 30311
rect 25605 30277 25639 30311
rect 25639 30277 25648 30311
rect 26148 30311 26200 30320
rect 25596 30268 25648 30277
rect 26148 30277 26157 30311
rect 26157 30277 26191 30311
rect 26191 30277 26200 30311
rect 26148 30268 26200 30277
rect 15384 30200 15436 30252
rect 17500 30200 17552 30252
rect 17868 30200 17920 30252
rect 24860 30243 24912 30252
rect 24860 30209 24869 30243
rect 24869 30209 24903 30243
rect 24903 30209 24912 30243
rect 24860 30200 24912 30209
rect 34612 30268 34664 30320
rect 34428 30243 34480 30252
rect 34428 30209 34437 30243
rect 34437 30209 34471 30243
rect 34471 30209 34480 30243
rect 34428 30200 34480 30209
rect 38292 30243 38344 30252
rect 38292 30209 38301 30243
rect 38301 30209 38335 30243
rect 38335 30209 38344 30243
rect 38292 30200 38344 30209
rect 8300 29996 8352 30048
rect 8668 29996 8720 30048
rect 10416 30064 10468 30116
rect 12440 30064 12492 30116
rect 17684 30132 17736 30184
rect 19432 30132 19484 30184
rect 15844 30107 15896 30116
rect 15844 30073 15853 30107
rect 15853 30073 15887 30107
rect 15887 30073 15896 30107
rect 15844 30064 15896 30073
rect 20444 30064 20496 30116
rect 25044 30064 25096 30116
rect 34244 30107 34296 30116
rect 34244 30073 34253 30107
rect 34253 30073 34287 30107
rect 34287 30073 34296 30107
rect 34244 30064 34296 30073
rect 10140 29996 10192 30048
rect 10324 29996 10376 30048
rect 12716 29996 12768 30048
rect 13728 29996 13780 30048
rect 13820 29996 13872 30048
rect 37004 29996 37056 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2228 29656 2280 29708
rect 3700 29656 3752 29708
rect 4068 29656 4120 29708
rect 1860 29631 1912 29640
rect 1860 29597 1869 29631
rect 1869 29597 1903 29631
rect 1903 29597 1912 29631
rect 5448 29792 5500 29844
rect 9864 29792 9916 29844
rect 10140 29792 10192 29844
rect 10876 29792 10928 29844
rect 11152 29792 11204 29844
rect 11336 29792 11388 29844
rect 12164 29792 12216 29844
rect 5908 29656 5960 29708
rect 1860 29588 1912 29597
rect 9128 29724 9180 29776
rect 23572 29792 23624 29844
rect 7104 29656 7156 29708
rect 12992 29724 13044 29776
rect 13084 29724 13136 29776
rect 13268 29724 13320 29776
rect 15108 29724 15160 29776
rect 15844 29724 15896 29776
rect 19616 29724 19668 29776
rect 7656 29588 7708 29640
rect 7932 29631 7984 29640
rect 7932 29597 7941 29631
rect 7941 29597 7975 29631
rect 7975 29597 7984 29631
rect 7932 29588 7984 29597
rect 4528 29520 4580 29572
rect 7012 29520 7064 29572
rect 7104 29520 7156 29572
rect 8208 29520 8260 29572
rect 3332 29452 3384 29504
rect 4068 29452 4120 29504
rect 8760 29588 8812 29640
rect 12716 29656 12768 29708
rect 14188 29656 14240 29708
rect 10876 29588 10928 29640
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 13728 29631 13780 29640
rect 8668 29520 8720 29572
rect 8944 29520 8996 29572
rect 8576 29495 8628 29504
rect 8576 29461 8585 29495
rect 8585 29461 8619 29495
rect 8619 29461 8628 29495
rect 11888 29520 11940 29572
rect 11980 29520 12032 29572
rect 12532 29520 12584 29572
rect 13728 29597 13737 29631
rect 13737 29597 13771 29631
rect 13771 29597 13780 29631
rect 13728 29588 13780 29597
rect 16304 29656 16356 29708
rect 15016 29588 15068 29640
rect 19524 29656 19576 29708
rect 18880 29631 18932 29640
rect 18880 29597 18889 29631
rect 18889 29597 18923 29631
rect 18923 29597 18932 29631
rect 18880 29588 18932 29597
rect 19156 29588 19208 29640
rect 10876 29495 10928 29504
rect 8576 29452 8628 29461
rect 10876 29461 10885 29495
rect 10885 29461 10919 29495
rect 10919 29461 10928 29495
rect 10876 29452 10928 29461
rect 12992 29452 13044 29504
rect 14464 29495 14516 29504
rect 14464 29461 14473 29495
rect 14473 29461 14507 29495
rect 14507 29461 14516 29495
rect 14464 29452 14516 29461
rect 17040 29452 17092 29504
rect 19248 29452 19300 29504
rect 19800 29588 19852 29640
rect 20352 29588 20404 29640
rect 25136 29588 25188 29640
rect 20812 29520 20864 29572
rect 19800 29452 19852 29504
rect 20168 29452 20220 29504
rect 21272 29452 21324 29504
rect 22192 29452 22244 29504
rect 24952 29452 25004 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1860 29248 1912 29300
rect 4068 29248 4120 29300
rect 5264 29180 5316 29232
rect 1584 29112 1636 29164
rect 4068 29112 4120 29164
rect 4896 29155 4948 29164
rect 4896 29121 4905 29155
rect 4905 29121 4939 29155
rect 4939 29121 4948 29155
rect 4896 29112 4948 29121
rect 8576 29248 8628 29300
rect 8668 29248 8720 29300
rect 10140 29248 10192 29300
rect 7196 29180 7248 29232
rect 7104 29155 7156 29164
rect 7104 29121 7113 29155
rect 7113 29121 7147 29155
rect 7147 29121 7156 29155
rect 7104 29112 7156 29121
rect 7380 29112 7432 29164
rect 7932 29112 7984 29164
rect 8760 29180 8812 29232
rect 14280 29248 14332 29300
rect 10600 29223 10652 29232
rect 10600 29189 10609 29223
rect 10609 29189 10643 29223
rect 10643 29189 10652 29223
rect 10600 29180 10652 29189
rect 10784 29180 10836 29232
rect 12256 29180 12308 29232
rect 14096 29180 14148 29232
rect 14464 29180 14516 29232
rect 11704 29155 11756 29164
rect 11704 29121 11713 29155
rect 11713 29121 11747 29155
rect 11747 29121 11756 29155
rect 11704 29112 11756 29121
rect 4896 28976 4948 29028
rect 9772 29044 9824 29096
rect 9956 29087 10008 29096
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10324 29044 10376 29096
rect 10508 29087 10560 29096
rect 10508 29053 10517 29087
rect 10517 29053 10551 29087
rect 10551 29053 10560 29087
rect 10508 29044 10560 29053
rect 11336 29044 11388 29096
rect 12440 29044 12492 29096
rect 12532 29044 12584 29096
rect 13912 29112 13964 29164
rect 14188 29155 14240 29164
rect 14188 29121 14197 29155
rect 14197 29121 14231 29155
rect 14231 29121 14240 29155
rect 14188 29112 14240 29121
rect 15016 29155 15068 29164
rect 15016 29121 15025 29155
rect 15025 29121 15059 29155
rect 15059 29121 15068 29155
rect 15016 29112 15068 29121
rect 19156 29248 19208 29300
rect 17040 29155 17092 29164
rect 17040 29121 17049 29155
rect 17049 29121 17083 29155
rect 17083 29121 17092 29155
rect 17040 29112 17092 29121
rect 19340 29180 19392 29232
rect 18052 29112 18104 29164
rect 20168 29155 20220 29164
rect 20168 29121 20177 29155
rect 20177 29121 20211 29155
rect 20211 29121 20220 29155
rect 20168 29112 20220 29121
rect 21364 29112 21416 29164
rect 22928 29248 22980 29300
rect 23572 29180 23624 29232
rect 23388 29155 23440 29164
rect 23388 29121 23397 29155
rect 23397 29121 23431 29155
rect 23431 29121 23440 29155
rect 23388 29112 23440 29121
rect 30380 29112 30432 29164
rect 18420 29087 18472 29096
rect 9588 28976 9640 29028
rect 10600 28976 10652 29028
rect 13176 28976 13228 29028
rect 14280 29019 14332 29028
rect 14280 28985 14289 29019
rect 14289 28985 14323 29019
rect 14323 28985 14332 29019
rect 14280 28976 14332 28985
rect 15200 28976 15252 29028
rect 16764 28976 16816 29028
rect 18420 29053 18429 29087
rect 18429 29053 18463 29087
rect 18463 29053 18472 29087
rect 18420 29044 18472 29053
rect 32404 29180 32456 29232
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 18236 28976 18288 29028
rect 20996 28976 21048 29028
rect 22008 29019 22060 29028
rect 22008 28985 22017 29019
rect 22017 28985 22051 29019
rect 22051 28985 22060 29019
rect 22008 28976 22060 28985
rect 23296 28976 23348 29028
rect 35440 28976 35492 29028
rect 2320 28908 2372 28960
rect 5816 28908 5868 28960
rect 8208 28908 8260 28960
rect 9864 28908 9916 28960
rect 9956 28908 10008 28960
rect 11244 28908 11296 28960
rect 11612 28908 11664 28960
rect 11980 28908 12032 28960
rect 22836 28951 22888 28960
rect 22836 28917 22845 28951
rect 22845 28917 22879 28951
rect 22879 28917 22888 28951
rect 22836 28908 22888 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2596 28704 2648 28756
rect 4528 28704 4580 28756
rect 7748 28704 7800 28756
rect 9588 28704 9640 28756
rect 1860 28611 1912 28620
rect 1860 28577 1869 28611
rect 1869 28577 1903 28611
rect 1903 28577 1912 28611
rect 1860 28568 1912 28577
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 7564 28636 7616 28688
rect 4988 28611 5040 28620
rect 4988 28577 4997 28611
rect 4997 28577 5031 28611
rect 5031 28577 5040 28611
rect 4988 28568 5040 28577
rect 5816 28568 5868 28620
rect 10692 28704 10744 28756
rect 10784 28704 10836 28756
rect 11428 28636 11480 28688
rect 14096 28636 14148 28688
rect 14648 28636 14700 28688
rect 18880 28704 18932 28756
rect 17868 28636 17920 28688
rect 10048 28611 10100 28620
rect 4436 28500 4488 28552
rect 5448 28500 5500 28552
rect 5908 28543 5960 28552
rect 5908 28509 5917 28543
rect 5917 28509 5951 28543
rect 5951 28509 5960 28543
rect 5908 28500 5960 28509
rect 3424 28432 3476 28484
rect 4988 28432 5040 28484
rect 10048 28577 10057 28611
rect 10057 28577 10091 28611
rect 10091 28577 10100 28611
rect 10048 28568 10100 28577
rect 10416 28568 10468 28620
rect 10876 28568 10928 28620
rect 9956 28500 10008 28552
rect 4252 28407 4304 28416
rect 4252 28373 4261 28407
rect 4261 28373 4295 28407
rect 4295 28373 4304 28407
rect 4252 28364 4304 28373
rect 4528 28364 4580 28416
rect 10600 28432 10652 28484
rect 10784 28432 10836 28484
rect 11980 28500 12032 28552
rect 12716 28543 12768 28552
rect 12716 28509 12725 28543
rect 12725 28509 12759 28543
rect 12759 28509 12768 28543
rect 12716 28500 12768 28509
rect 12348 28432 12400 28484
rect 17684 28568 17736 28620
rect 24032 28704 24084 28756
rect 24584 28636 24636 28688
rect 14372 28500 14424 28552
rect 15016 28500 15068 28552
rect 15476 28500 15528 28552
rect 16856 28543 16908 28552
rect 16856 28509 16865 28543
rect 16865 28509 16899 28543
rect 16899 28509 16908 28543
rect 16856 28500 16908 28509
rect 18052 28500 18104 28552
rect 19984 28611 20036 28620
rect 19984 28577 19993 28611
rect 19993 28577 20027 28611
rect 20027 28577 20036 28611
rect 19984 28568 20036 28577
rect 20260 28568 20312 28620
rect 20812 28611 20864 28620
rect 20812 28577 20821 28611
rect 20821 28577 20855 28611
rect 20855 28577 20864 28611
rect 20812 28568 20864 28577
rect 22744 28611 22796 28620
rect 22744 28577 22753 28611
rect 22753 28577 22787 28611
rect 22787 28577 22796 28611
rect 22744 28568 22796 28577
rect 22836 28568 22888 28620
rect 21916 28543 21968 28552
rect 21916 28509 21925 28543
rect 21925 28509 21959 28543
rect 21959 28509 21968 28543
rect 21916 28500 21968 28509
rect 17132 28432 17184 28484
rect 5448 28407 5500 28416
rect 5448 28373 5457 28407
rect 5457 28373 5491 28407
rect 5491 28373 5500 28407
rect 5448 28364 5500 28373
rect 6828 28364 6880 28416
rect 7932 28364 7984 28416
rect 11888 28364 11940 28416
rect 11980 28364 12032 28416
rect 12900 28364 12952 28416
rect 15660 28364 15712 28416
rect 15844 28407 15896 28416
rect 15844 28373 15853 28407
rect 15853 28373 15887 28407
rect 15887 28373 15896 28407
rect 15844 28364 15896 28373
rect 18604 28407 18656 28416
rect 18604 28373 18613 28407
rect 18613 28373 18647 28407
rect 18647 28373 18656 28407
rect 18604 28364 18656 28373
rect 21088 28364 21140 28416
rect 23664 28364 23716 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4252 28160 4304 28212
rect 8116 28160 8168 28212
rect 8208 28160 8260 28212
rect 10784 28160 10836 28212
rect 12716 28160 12768 28212
rect 12900 28160 12952 28212
rect 15016 28160 15068 28212
rect 18512 28160 18564 28212
rect 20720 28160 20772 28212
rect 1860 28135 1912 28144
rect 1860 28101 1869 28135
rect 1869 28101 1903 28135
rect 1903 28101 1912 28135
rect 1860 28092 1912 28101
rect 4344 28135 4396 28144
rect 4344 28101 4353 28135
rect 4353 28101 4387 28135
rect 4387 28101 4396 28135
rect 4344 28092 4396 28101
rect 4804 28092 4856 28144
rect 6920 28092 6972 28144
rect 9036 28135 9088 28144
rect 9036 28101 9045 28135
rect 9045 28101 9079 28135
rect 9079 28101 9088 28135
rect 9036 28092 9088 28101
rect 9680 28092 9732 28144
rect 10048 28092 10100 28144
rect 11980 28092 12032 28144
rect 13636 28092 13688 28144
rect 14648 28092 14700 28144
rect 2964 28024 3016 28076
rect 4068 28067 4120 28076
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 4068 28033 4077 28067
rect 4077 28033 4111 28067
rect 4111 28033 4120 28067
rect 4068 28024 4120 28033
rect 5908 28024 5960 28076
rect 6828 28024 6880 28076
rect 10692 28024 10744 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 14924 28024 14976 28076
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 16764 28024 16816 28076
rect 18052 28092 18104 28144
rect 21640 28160 21692 28212
rect 1584 27956 1636 27965
rect 3792 27956 3844 28008
rect 4436 27956 4488 28008
rect 4804 27956 4856 28008
rect 5816 27999 5868 28008
rect 5816 27965 5825 27999
rect 5825 27965 5859 27999
rect 5859 27965 5868 27999
rect 5816 27956 5868 27965
rect 7656 27956 7708 28008
rect 10508 27956 10560 28008
rect 12348 27956 12400 28008
rect 14464 27956 14516 28008
rect 16028 27956 16080 28008
rect 18512 27999 18564 28008
rect 8576 27888 8628 27940
rect 9312 27888 9364 27940
rect 10048 27888 10100 27940
rect 11704 27888 11756 27940
rect 13728 27888 13780 27940
rect 15476 27888 15528 27940
rect 18512 27965 18521 27999
rect 18521 27965 18555 27999
rect 18555 27965 18564 27999
rect 18512 27956 18564 27965
rect 21824 28024 21876 28076
rect 22192 28067 22244 28076
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 24952 28067 25004 28076
rect 20352 27956 20404 28008
rect 21732 27956 21784 28008
rect 20996 27888 21048 27940
rect 21916 27888 21968 27940
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 23480 27956 23532 28008
rect 5448 27820 5500 27872
rect 8668 27820 8720 27872
rect 9404 27820 9456 27872
rect 14372 27820 14424 27872
rect 14648 27820 14700 27872
rect 15752 27820 15804 27872
rect 16580 27820 16632 27872
rect 17500 27820 17552 27872
rect 19616 27820 19668 27872
rect 22192 27820 22244 27872
rect 24768 27863 24820 27872
rect 24768 27829 24777 27863
rect 24777 27829 24811 27863
rect 24811 27829 24820 27863
rect 24768 27820 24820 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1860 27659 1912 27668
rect 1860 27625 1890 27659
rect 1890 27625 1912 27659
rect 1860 27616 1912 27625
rect 8760 27616 8812 27668
rect 10968 27616 11020 27668
rect 11244 27616 11296 27668
rect 11704 27616 11756 27668
rect 13544 27616 13596 27668
rect 4068 27548 4120 27600
rect 4896 27548 4948 27600
rect 8668 27548 8720 27600
rect 15292 27616 15344 27668
rect 5908 27480 5960 27532
rect 6828 27480 6880 27532
rect 9128 27523 9180 27532
rect 9128 27489 9137 27523
rect 9137 27489 9171 27523
rect 9171 27489 9180 27523
rect 9128 27480 9180 27489
rect 9404 27523 9456 27532
rect 9404 27489 9413 27523
rect 9413 27489 9447 27523
rect 9447 27489 9456 27523
rect 9404 27480 9456 27489
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 3148 27412 3200 27464
rect 4896 27412 4948 27464
rect 7472 27412 7524 27464
rect 7656 27412 7708 27464
rect 7932 27455 7984 27464
rect 7932 27421 7941 27455
rect 7941 27421 7975 27455
rect 7975 27421 7984 27455
rect 7932 27412 7984 27421
rect 8116 27455 8168 27464
rect 8116 27421 8125 27455
rect 8125 27421 8159 27455
rect 8159 27421 8168 27455
rect 8116 27412 8168 27421
rect 8852 27412 8904 27464
rect 13912 27480 13964 27532
rect 18144 27548 18196 27600
rect 19984 27548 20036 27600
rect 21640 27591 21692 27600
rect 21640 27557 21649 27591
rect 21649 27557 21683 27591
rect 21683 27557 21692 27591
rect 21640 27548 21692 27557
rect 22744 27591 22796 27600
rect 22744 27557 22753 27591
rect 22753 27557 22787 27591
rect 22787 27557 22796 27591
rect 22744 27548 22796 27557
rect 23388 27548 23440 27600
rect 15660 27480 15712 27532
rect 18604 27480 18656 27532
rect 14464 27455 14516 27464
rect 4620 27344 4672 27396
rect 6736 27344 6788 27396
rect 7564 27344 7616 27396
rect 8944 27344 8996 27396
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 9312 27344 9364 27396
rect 11060 27344 11112 27396
rect 11704 27344 11756 27396
rect 12716 27344 12768 27396
rect 12992 27387 13044 27396
rect 12992 27353 13001 27387
rect 13001 27353 13035 27387
rect 13035 27353 13044 27387
rect 12992 27344 13044 27353
rect 15108 27387 15160 27396
rect 15108 27353 15117 27387
rect 15117 27353 15151 27387
rect 15151 27353 15160 27387
rect 15108 27344 15160 27353
rect 16212 27412 16264 27464
rect 17868 27412 17920 27464
rect 18788 27412 18840 27464
rect 19616 27455 19668 27464
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 21272 27455 21324 27464
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 22008 27480 22060 27532
rect 3424 27276 3476 27328
rect 5356 27276 5408 27328
rect 10324 27276 10376 27328
rect 13176 27276 13228 27328
rect 14832 27276 14884 27328
rect 18696 27344 18748 27396
rect 19248 27344 19300 27396
rect 16764 27319 16816 27328
rect 16764 27285 16773 27319
rect 16773 27285 16807 27319
rect 16807 27285 16816 27319
rect 16764 27276 16816 27285
rect 19064 27276 19116 27328
rect 23480 27412 23532 27464
rect 23572 27412 23624 27464
rect 24216 27412 24268 27464
rect 24308 27412 24360 27464
rect 35440 27412 35492 27464
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 23940 27344 23992 27396
rect 21548 27276 21600 27328
rect 23296 27276 23348 27328
rect 23480 27319 23532 27328
rect 23480 27285 23489 27319
rect 23489 27285 23523 27319
rect 23523 27285 23532 27319
rect 23480 27276 23532 27285
rect 23572 27276 23624 27328
rect 31760 27319 31812 27328
rect 31760 27285 31769 27319
rect 31769 27285 31803 27319
rect 31803 27285 31812 27319
rect 31760 27276 31812 27285
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1768 27115 1820 27124
rect 1768 27081 1777 27115
rect 1777 27081 1811 27115
rect 1811 27081 1820 27115
rect 1768 27072 1820 27081
rect 3148 27072 3200 27124
rect 9680 27072 9732 27124
rect 3608 27047 3660 27056
rect 3608 27013 3617 27047
rect 3617 27013 3651 27047
rect 3651 27013 3660 27047
rect 3608 27004 3660 27013
rect 5356 27047 5408 27056
rect 5356 27013 5365 27047
rect 5365 27013 5399 27047
rect 5399 27013 5408 27047
rect 5356 27004 5408 27013
rect 5724 27004 5776 27056
rect 8944 27004 8996 27056
rect 11704 27072 11756 27124
rect 11520 27004 11572 27056
rect 11888 27047 11940 27056
rect 11888 27013 11897 27047
rect 11897 27013 11931 27047
rect 11931 27013 11940 27047
rect 11888 27004 11940 27013
rect 1952 26936 2004 26988
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 4712 26936 4764 26988
rect 6092 26936 6144 26988
rect 6828 26936 6880 26988
rect 9128 26936 9180 26988
rect 14556 27004 14608 27056
rect 17500 27072 17552 27124
rect 18696 27115 18748 27124
rect 18696 27081 18705 27115
rect 18705 27081 18739 27115
rect 18739 27081 18748 27115
rect 18696 27072 18748 27081
rect 18788 27072 18840 27124
rect 21548 27072 21600 27124
rect 25320 27072 25372 27124
rect 34428 27072 34480 27124
rect 1676 26868 1728 26920
rect 8576 26868 8628 26920
rect 11244 26868 11296 26920
rect 12532 26868 12584 26920
rect 13728 26936 13780 26988
rect 14280 26936 14332 26988
rect 14556 26868 14608 26920
rect 15660 27004 15712 27056
rect 15752 27004 15804 27056
rect 16672 27004 16724 27056
rect 14832 26868 14884 26920
rect 15476 26868 15528 26920
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 21824 27004 21876 27056
rect 18328 26936 18380 26988
rect 19064 26936 19116 26988
rect 22836 27004 22888 27056
rect 24768 26936 24820 26988
rect 37004 26936 37056 26988
rect 18236 26911 18288 26920
rect 18236 26877 18245 26911
rect 18245 26877 18279 26911
rect 18279 26877 18288 26911
rect 18236 26868 18288 26877
rect 20260 26911 20312 26920
rect 20260 26877 20269 26911
rect 20269 26877 20303 26911
rect 20303 26877 20312 26911
rect 20260 26868 20312 26877
rect 20720 26868 20772 26920
rect 22192 26911 22244 26920
rect 7012 26800 7064 26852
rect 5724 26732 5776 26784
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 12164 26800 12216 26852
rect 12256 26800 12308 26852
rect 10968 26775 11020 26784
rect 10968 26741 10977 26775
rect 10977 26741 11011 26775
rect 11011 26741 11020 26775
rect 12900 26775 12952 26784
rect 10968 26732 11020 26741
rect 12900 26741 12909 26775
rect 12909 26741 12943 26775
rect 12943 26741 12952 26775
rect 12900 26732 12952 26741
rect 13636 26775 13688 26784
rect 13636 26741 13645 26775
rect 13645 26741 13679 26775
rect 13679 26741 13688 26775
rect 13636 26732 13688 26741
rect 14004 26800 14056 26852
rect 16764 26800 16816 26852
rect 17592 26800 17644 26852
rect 19984 26800 20036 26852
rect 22192 26877 22201 26911
rect 22201 26877 22235 26911
rect 22235 26877 22244 26911
rect 22192 26868 22244 26877
rect 23296 26911 23348 26920
rect 23296 26877 23305 26911
rect 23305 26877 23339 26911
rect 23339 26877 23348 26911
rect 23296 26868 23348 26877
rect 24492 26911 24544 26920
rect 24492 26877 24501 26911
rect 24501 26877 24535 26911
rect 24535 26877 24544 26911
rect 24492 26868 24544 26877
rect 17316 26732 17368 26784
rect 17500 26775 17552 26784
rect 17500 26741 17509 26775
rect 17509 26741 17543 26775
rect 17543 26741 17552 26775
rect 17500 26732 17552 26741
rect 20904 26732 20956 26784
rect 31760 26800 31812 26852
rect 24032 26732 24084 26784
rect 32588 26775 32640 26784
rect 32588 26741 32597 26775
rect 32597 26741 32631 26775
rect 32631 26741 32640 26775
rect 32588 26732 32640 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5724 26571 5776 26580
rect 5724 26537 5733 26571
rect 5733 26537 5767 26571
rect 5767 26537 5776 26571
rect 5724 26528 5776 26537
rect 10968 26528 11020 26580
rect 12532 26528 12584 26580
rect 18420 26528 18472 26580
rect 19524 26528 19576 26580
rect 23296 26528 23348 26580
rect 38016 26528 38068 26580
rect 3608 26460 3660 26512
rect 3976 26435 4028 26444
rect 3976 26401 3985 26435
rect 3985 26401 4019 26435
rect 4019 26401 4028 26435
rect 3976 26392 4028 26401
rect 5816 26392 5868 26444
rect 6828 26435 6880 26444
rect 6828 26401 6837 26435
rect 6837 26401 6871 26435
rect 6871 26401 6880 26435
rect 6828 26392 6880 26401
rect 9404 26460 9456 26512
rect 9588 26460 9640 26512
rect 11336 26460 11388 26512
rect 12256 26460 12308 26512
rect 16764 26503 16816 26512
rect 14372 26392 14424 26444
rect 14648 26435 14700 26444
rect 14648 26401 14657 26435
rect 14657 26401 14691 26435
rect 14691 26401 14700 26435
rect 14648 26392 14700 26401
rect 16764 26469 16773 26503
rect 16773 26469 16807 26503
rect 16807 26469 16816 26503
rect 16764 26460 16816 26469
rect 18696 26460 18748 26512
rect 21364 26460 21416 26512
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 2872 26256 2924 26308
rect 3884 26256 3936 26308
rect 5632 26256 5684 26308
rect 4528 26188 4580 26240
rect 7104 26188 7156 26240
rect 7748 26188 7800 26240
rect 9496 26256 9548 26308
rect 11244 26324 11296 26376
rect 12072 26324 12124 26376
rect 13176 26324 13228 26376
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 14280 26324 14332 26376
rect 15568 26324 15620 26376
rect 16212 26324 16264 26376
rect 16672 26324 16724 26376
rect 17316 26324 17368 26376
rect 18052 26324 18104 26376
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 20352 26324 20404 26376
rect 26332 26460 26384 26512
rect 23572 26435 23624 26444
rect 23572 26401 23581 26435
rect 23581 26401 23615 26435
rect 23615 26401 23624 26435
rect 23572 26392 23624 26401
rect 23756 26392 23808 26444
rect 23480 26324 23532 26376
rect 19524 26299 19576 26308
rect 13176 26188 13228 26240
rect 13544 26231 13596 26240
rect 13544 26197 13553 26231
rect 13553 26197 13587 26231
rect 13587 26197 13596 26231
rect 13544 26188 13596 26197
rect 14464 26188 14516 26240
rect 15660 26188 15712 26240
rect 17316 26188 17368 26240
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 21456 26256 21508 26308
rect 24952 26256 25004 26308
rect 34520 26324 34572 26376
rect 20628 26231 20680 26240
rect 20628 26197 20637 26231
rect 20637 26197 20671 26231
rect 20671 26197 20680 26231
rect 20628 26188 20680 26197
rect 20812 26188 20864 26240
rect 21916 26231 21968 26240
rect 21916 26197 21925 26231
rect 21925 26197 21959 26231
rect 21959 26197 21968 26231
rect 21916 26188 21968 26197
rect 22652 26231 22704 26240
rect 22652 26197 22661 26231
rect 22661 26197 22695 26231
rect 22695 26197 22704 26231
rect 22652 26188 22704 26197
rect 24124 26188 24176 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4528 25984 4580 26036
rect 4712 25984 4764 26036
rect 12164 25984 12216 26036
rect 15200 25984 15252 26036
rect 18328 25984 18380 26036
rect 20352 25984 20404 26036
rect 4620 25916 4672 25968
rect 5080 25916 5132 25968
rect 5908 25916 5960 25968
rect 8944 25916 8996 25968
rect 3976 25848 4028 25900
rect 6920 25848 6972 25900
rect 11704 25848 11756 25900
rect 12072 25891 12124 25900
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 12164 25848 12216 25900
rect 1584 25823 1636 25832
rect 1584 25789 1593 25823
rect 1593 25789 1627 25823
rect 1627 25789 1636 25823
rect 1584 25780 1636 25789
rect 3608 25823 3660 25832
rect 3608 25789 3617 25823
rect 3617 25789 3651 25823
rect 3651 25789 3660 25823
rect 3608 25780 3660 25789
rect 5816 25823 5868 25832
rect 5816 25789 5825 25823
rect 5825 25789 5859 25823
rect 5859 25789 5868 25823
rect 5816 25780 5868 25789
rect 7104 25823 7156 25832
rect 7104 25789 7113 25823
rect 7113 25789 7147 25823
rect 7147 25789 7156 25823
rect 7104 25780 7156 25789
rect 7472 25780 7524 25832
rect 1492 25644 1544 25696
rect 3976 25644 4028 25696
rect 5448 25712 5500 25764
rect 4712 25644 4764 25696
rect 10784 25712 10836 25764
rect 10876 25712 10928 25764
rect 12900 25848 12952 25900
rect 13636 25916 13688 25968
rect 14004 25848 14056 25900
rect 14096 25891 14148 25900
rect 14096 25857 14105 25891
rect 14105 25857 14139 25891
rect 14139 25857 14148 25891
rect 14096 25848 14148 25857
rect 15292 25848 15344 25900
rect 15476 25848 15528 25900
rect 17408 25848 17460 25900
rect 17592 25848 17644 25900
rect 19432 25916 19484 25968
rect 19156 25891 19208 25900
rect 17040 25780 17092 25832
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 20720 25984 20772 26036
rect 20812 25959 20864 25968
rect 20812 25925 20821 25959
rect 20821 25925 20855 25959
rect 20855 25925 20864 25959
rect 20812 25916 20864 25925
rect 20904 25959 20956 25968
rect 20904 25925 20913 25959
rect 20913 25925 20947 25959
rect 20947 25925 20956 25959
rect 21456 25959 21508 25968
rect 20904 25916 20956 25925
rect 21456 25925 21465 25959
rect 21465 25925 21499 25959
rect 21499 25925 21508 25959
rect 21456 25916 21508 25925
rect 23112 25916 23164 25968
rect 26608 25916 26660 25968
rect 23756 25891 23808 25900
rect 23756 25857 23765 25891
rect 23765 25857 23799 25891
rect 23799 25857 23808 25891
rect 23756 25848 23808 25857
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 9956 25687 10008 25696
rect 9956 25653 9965 25687
rect 9965 25653 9999 25687
rect 9999 25653 10008 25687
rect 9956 25644 10008 25653
rect 11244 25644 11296 25696
rect 12532 25644 12584 25696
rect 13268 25644 13320 25696
rect 14096 25644 14148 25696
rect 17224 25712 17276 25764
rect 21916 25780 21968 25832
rect 19984 25755 20036 25764
rect 19984 25721 19993 25755
rect 19993 25721 20027 25755
rect 20027 25721 20036 25755
rect 19984 25712 20036 25721
rect 21732 25712 21784 25764
rect 23112 25712 23164 25764
rect 16120 25644 16172 25696
rect 18236 25687 18288 25696
rect 18236 25653 18245 25687
rect 18245 25653 18279 25687
rect 18279 25653 18288 25687
rect 18236 25644 18288 25653
rect 21456 25644 21508 25696
rect 23848 25687 23900 25696
rect 23848 25653 23857 25687
rect 23857 25653 23891 25687
rect 23891 25653 23900 25687
rect 23848 25644 23900 25653
rect 38016 25644 38068 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3976 25483 4028 25492
rect 3976 25449 3985 25483
rect 3985 25449 4019 25483
rect 4019 25449 4028 25483
rect 3976 25440 4028 25449
rect 5540 25483 5592 25492
rect 5540 25449 5549 25483
rect 5549 25449 5583 25483
rect 5583 25449 5592 25483
rect 5540 25440 5592 25449
rect 7196 25440 7248 25492
rect 7472 25483 7524 25492
rect 7472 25449 7481 25483
rect 7481 25449 7515 25483
rect 7515 25449 7524 25483
rect 7472 25440 7524 25449
rect 3608 25372 3660 25424
rect 1584 25347 1636 25356
rect 1584 25313 1593 25347
rect 1593 25313 1627 25347
rect 1627 25313 1636 25347
rect 1584 25304 1636 25313
rect 2504 25304 2556 25356
rect 5172 25304 5224 25356
rect 11152 25372 11204 25424
rect 16580 25483 16632 25492
rect 3976 25168 4028 25220
rect 4344 25236 4396 25288
rect 5724 25279 5776 25288
rect 5724 25245 5733 25279
rect 5733 25245 5767 25279
rect 5767 25245 5776 25279
rect 5724 25236 5776 25245
rect 5908 25236 5960 25288
rect 7380 25279 7432 25288
rect 7380 25245 7389 25279
rect 7389 25245 7423 25279
rect 7423 25245 7432 25279
rect 7380 25236 7432 25245
rect 6644 25168 6696 25220
rect 2688 25100 2740 25152
rect 4988 25143 5040 25152
rect 4988 25109 4997 25143
rect 4997 25109 5031 25143
rect 5031 25109 5040 25143
rect 4988 25100 5040 25109
rect 9220 25236 9272 25288
rect 9588 25236 9640 25288
rect 9956 25168 10008 25220
rect 11060 25236 11112 25288
rect 11336 25236 11388 25288
rect 11796 25236 11848 25288
rect 13544 25304 13596 25356
rect 14372 25304 14424 25356
rect 15108 25304 15160 25356
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 16580 25449 16589 25483
rect 16589 25449 16623 25483
rect 16623 25449 16632 25483
rect 16580 25440 16632 25449
rect 17316 25440 17368 25492
rect 17592 25440 17644 25492
rect 18144 25440 18196 25492
rect 18880 25440 18932 25492
rect 20996 25440 21048 25492
rect 22744 25440 22796 25492
rect 23664 25440 23716 25492
rect 23756 25372 23808 25424
rect 24768 25372 24820 25424
rect 17224 25347 17276 25356
rect 17224 25313 17233 25347
rect 17233 25313 17267 25347
rect 17267 25313 17276 25347
rect 17224 25304 17276 25313
rect 17500 25304 17552 25356
rect 20260 25347 20312 25356
rect 20260 25313 20269 25347
rect 20269 25313 20303 25347
rect 20303 25313 20312 25347
rect 20260 25304 20312 25313
rect 20628 25304 20680 25356
rect 22652 25304 22704 25356
rect 24124 25304 24176 25356
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17868 25236 17920 25288
rect 19340 25236 19392 25288
rect 19432 25236 19484 25288
rect 21548 25236 21600 25288
rect 13084 25211 13136 25220
rect 9036 25100 9088 25152
rect 10048 25100 10100 25152
rect 10232 25100 10284 25152
rect 11612 25100 11664 25152
rect 11796 25143 11848 25152
rect 11796 25109 11805 25143
rect 11805 25109 11839 25143
rect 11839 25109 11848 25143
rect 11796 25100 11848 25109
rect 13084 25177 13093 25211
rect 13093 25177 13127 25211
rect 13127 25177 13136 25211
rect 13084 25168 13136 25177
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13728 25211 13780 25220
rect 13176 25168 13228 25177
rect 13728 25177 13737 25211
rect 13737 25177 13771 25211
rect 13771 25177 13780 25211
rect 13728 25168 13780 25177
rect 14004 25168 14056 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 14832 25168 14884 25220
rect 18972 25168 19024 25220
rect 21180 25168 21232 25220
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 25872 25236 25924 25288
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 15384 25100 15436 25152
rect 20812 25100 20864 25152
rect 24676 25143 24728 25152
rect 24676 25109 24685 25143
rect 24685 25109 24719 25143
rect 24719 25109 24728 25143
rect 24676 25100 24728 25109
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2412 24896 2464 24948
rect 12164 24896 12216 24948
rect 15936 24896 15988 24948
rect 3516 24828 3568 24880
rect 5816 24828 5868 24880
rect 12256 24828 12308 24880
rect 13084 24828 13136 24880
rect 14832 24828 14884 24880
rect 1768 24803 1820 24812
rect 1768 24769 1777 24803
rect 1777 24769 1811 24803
rect 1811 24769 1820 24803
rect 1768 24760 1820 24769
rect 2504 24803 2556 24812
rect 2504 24769 2513 24803
rect 2513 24769 2547 24803
rect 2547 24769 2556 24803
rect 2504 24760 2556 24769
rect 4068 24760 4120 24812
rect 5080 24803 5132 24812
rect 5080 24769 5089 24803
rect 5089 24769 5123 24803
rect 5123 24769 5132 24803
rect 5080 24760 5132 24769
rect 5540 24803 5592 24812
rect 5540 24769 5549 24803
rect 5549 24769 5583 24803
rect 5583 24769 5592 24803
rect 5540 24760 5592 24769
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 4712 24692 4764 24744
rect 7104 24692 7156 24744
rect 4344 24624 4396 24676
rect 4896 24667 4948 24676
rect 4896 24633 4905 24667
rect 4905 24633 4939 24667
rect 4939 24633 4948 24667
rect 4896 24624 4948 24633
rect 9220 24760 9272 24812
rect 9404 24803 9456 24812
rect 9404 24769 9413 24803
rect 9413 24769 9447 24803
rect 9447 24769 9456 24803
rect 9404 24760 9456 24769
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 10140 24760 10192 24812
rect 10600 24760 10652 24812
rect 24676 24828 24728 24880
rect 18512 24803 18564 24812
rect 14004 24735 14056 24744
rect 7748 24599 7800 24608
rect 7748 24565 7757 24599
rect 7757 24565 7791 24599
rect 7791 24565 7800 24599
rect 7748 24556 7800 24565
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 9588 24624 9640 24676
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 15200 24735 15252 24744
rect 15200 24701 15209 24735
rect 15209 24701 15243 24735
rect 15243 24701 15252 24735
rect 15200 24692 15252 24701
rect 16396 24692 16448 24744
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 18696 24803 18748 24812
rect 18696 24769 18705 24803
rect 18705 24769 18739 24803
rect 18739 24769 18748 24803
rect 18696 24760 18748 24769
rect 19432 24760 19484 24812
rect 20812 24760 20864 24812
rect 17684 24667 17736 24676
rect 11888 24556 11940 24608
rect 13912 24556 13964 24608
rect 17684 24633 17693 24667
rect 17693 24633 17727 24667
rect 17727 24633 17736 24667
rect 17684 24624 17736 24633
rect 18880 24667 18932 24676
rect 18880 24633 18889 24667
rect 18889 24633 18923 24667
rect 18923 24633 18932 24667
rect 18880 24624 18932 24633
rect 20168 24692 20220 24744
rect 21364 24624 21416 24676
rect 16028 24556 16080 24608
rect 20536 24556 20588 24608
rect 20996 24599 21048 24608
rect 20996 24565 21005 24599
rect 21005 24565 21039 24599
rect 21039 24565 21048 24599
rect 20996 24556 21048 24565
rect 22284 24599 22336 24608
rect 22284 24565 22293 24599
rect 22293 24565 22327 24599
rect 22327 24565 22336 24599
rect 22284 24556 22336 24565
rect 24400 24760 24452 24812
rect 26332 24760 26384 24812
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 34520 24760 34572 24812
rect 23664 24692 23716 24744
rect 23756 24667 23808 24676
rect 23756 24633 23765 24667
rect 23765 24633 23799 24667
rect 23799 24633 23808 24667
rect 23756 24624 23808 24633
rect 24400 24556 24452 24608
rect 25596 24599 25648 24608
rect 25596 24565 25605 24599
rect 25605 24565 25639 24599
rect 25639 24565 25648 24599
rect 25596 24556 25648 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2412 24395 2464 24404
rect 2412 24361 2421 24395
rect 2421 24361 2455 24395
rect 2455 24361 2464 24395
rect 2412 24352 2464 24361
rect 3056 24395 3108 24404
rect 3056 24361 3065 24395
rect 3065 24361 3099 24395
rect 3099 24361 3108 24395
rect 3056 24352 3108 24361
rect 4068 24395 4120 24404
rect 4068 24361 4077 24395
rect 4077 24361 4111 24395
rect 4111 24361 4120 24395
rect 4068 24352 4120 24361
rect 5080 24352 5132 24404
rect 6000 24352 6052 24404
rect 8484 24352 8536 24404
rect 9680 24352 9732 24404
rect 9956 24395 10008 24404
rect 9956 24361 9965 24395
rect 9965 24361 9999 24395
rect 9999 24361 10008 24395
rect 9956 24352 10008 24361
rect 12348 24352 12400 24404
rect 1400 24284 1452 24336
rect 3332 24216 3384 24268
rect 3240 24148 3292 24200
rect 3700 24148 3752 24200
rect 9404 24284 9456 24336
rect 4804 24216 4856 24268
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 8852 24216 8904 24268
rect 10692 24216 10744 24268
rect 7564 24191 7616 24200
rect 7564 24157 7573 24191
rect 7573 24157 7607 24191
rect 7607 24157 7616 24191
rect 7564 24148 7616 24157
rect 10416 24148 10468 24200
rect 11152 24259 11204 24268
rect 11152 24225 11161 24259
rect 11161 24225 11195 24259
rect 11195 24225 11204 24259
rect 11152 24216 11204 24225
rect 11336 24216 11388 24268
rect 11704 24216 11756 24268
rect 11980 24216 12032 24268
rect 12256 24191 12308 24200
rect 10048 24080 10100 24132
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 12348 24148 12400 24200
rect 14188 24352 14240 24404
rect 17500 24352 17552 24404
rect 13360 24284 13412 24336
rect 16304 24284 16356 24336
rect 16396 24284 16448 24336
rect 17132 24284 17184 24336
rect 19708 24352 19760 24404
rect 23940 24352 23992 24404
rect 24952 24395 25004 24404
rect 24952 24361 24961 24395
rect 24961 24361 24995 24395
rect 24995 24361 25004 24395
rect 24952 24352 25004 24361
rect 26332 24395 26384 24404
rect 26332 24361 26341 24395
rect 26341 24361 26375 24395
rect 26375 24361 26384 24395
rect 26332 24352 26384 24361
rect 19432 24284 19484 24336
rect 24308 24284 24360 24336
rect 13452 24216 13504 24268
rect 11980 24080 12032 24132
rect 12072 24080 12124 24132
rect 14096 24148 14148 24200
rect 16856 24148 16908 24200
rect 19708 24191 19760 24200
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 11520 24012 11572 24064
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 14188 24012 14240 24064
rect 15292 24055 15344 24064
rect 15292 24021 15301 24055
rect 15301 24021 15335 24055
rect 15335 24021 15344 24055
rect 15292 24012 15344 24021
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 16672 24080 16724 24132
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 20536 24191 20588 24200
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24148 20588 24157
rect 23848 24216 23900 24268
rect 24492 24216 24544 24268
rect 25596 24216 25648 24268
rect 25872 24191 25924 24200
rect 25872 24157 25881 24191
rect 25881 24157 25915 24191
rect 25915 24157 25924 24191
rect 25872 24148 25924 24157
rect 26608 24148 26660 24200
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 18144 24080 18196 24132
rect 27528 24080 27580 24132
rect 16580 24012 16632 24064
rect 17776 24012 17828 24064
rect 18512 24055 18564 24064
rect 18512 24021 18521 24055
rect 18521 24021 18555 24055
rect 18555 24021 18564 24055
rect 18512 24012 18564 24021
rect 19984 24012 20036 24064
rect 20352 24055 20404 24064
rect 20352 24021 20361 24055
rect 20361 24021 20395 24055
rect 20395 24021 20404 24055
rect 20352 24012 20404 24021
rect 21456 24012 21508 24064
rect 22744 24012 22796 24064
rect 25688 24055 25740 24064
rect 25688 24021 25697 24055
rect 25697 24021 25731 24055
rect 25731 24021 25740 24055
rect 25688 24012 25740 24021
rect 30196 24012 30248 24064
rect 38108 24055 38160 24064
rect 38108 24021 38117 24055
rect 38117 24021 38151 24055
rect 38151 24021 38160 24055
rect 38108 24012 38160 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2136 23808 2188 23860
rect 5632 23808 5684 23860
rect 3608 23783 3660 23792
rect 3608 23749 3617 23783
rect 3617 23749 3651 23783
rect 3651 23749 3660 23783
rect 3608 23740 3660 23749
rect 1952 23672 2004 23724
rect 2780 23672 2832 23724
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 7012 23672 7064 23724
rect 8576 23672 8628 23724
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 11152 23715 11204 23724
rect 11152 23681 11161 23715
rect 11161 23681 11195 23715
rect 11195 23681 11204 23715
rect 11152 23672 11204 23681
rect 11336 23672 11388 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 11980 23808 12032 23860
rect 13820 23808 13872 23860
rect 15292 23808 15344 23860
rect 18052 23808 18104 23860
rect 18512 23808 18564 23860
rect 21088 23808 21140 23860
rect 12348 23740 12400 23792
rect 15016 23740 15068 23792
rect 20444 23740 20496 23792
rect 24400 23808 24452 23860
rect 22836 23783 22888 23792
rect 22836 23749 22845 23783
rect 22845 23749 22879 23783
rect 22879 23749 22888 23783
rect 22836 23740 22888 23749
rect 11980 23672 12032 23724
rect 13360 23672 13412 23724
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 17132 23672 17184 23724
rect 17776 23715 17828 23724
rect 17776 23681 17785 23715
rect 17785 23681 17819 23715
rect 17819 23681 17828 23715
rect 17776 23672 17828 23681
rect 18236 23672 18288 23724
rect 8300 23536 8352 23588
rect 8760 23536 8812 23588
rect 12716 23604 12768 23656
rect 13268 23604 13320 23656
rect 15016 23604 15068 23656
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 16580 23604 16632 23656
rect 20996 23672 21048 23724
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 24584 23715 24636 23724
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 11520 23536 11572 23588
rect 8668 23468 8720 23520
rect 11336 23468 11388 23520
rect 15476 23536 15528 23588
rect 17224 23536 17276 23588
rect 20260 23604 20312 23656
rect 22376 23604 22428 23656
rect 13360 23511 13412 23520
rect 13360 23477 13369 23511
rect 13369 23477 13403 23511
rect 13403 23477 13412 23511
rect 13360 23468 13412 23477
rect 17040 23468 17092 23520
rect 17868 23468 17920 23520
rect 20904 23468 20956 23520
rect 32588 23468 32640 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2596 23264 2648 23316
rect 6092 23264 6144 23316
rect 11060 23264 11112 23316
rect 11520 23307 11572 23316
rect 11520 23273 11529 23307
rect 11529 23273 11563 23307
rect 11563 23273 11572 23307
rect 11520 23264 11572 23273
rect 12164 23264 12216 23316
rect 6368 23196 6420 23248
rect 4988 23128 5040 23180
rect 9496 23128 9548 23180
rect 1676 23060 1728 23112
rect 1952 23060 2004 23112
rect 5264 23060 5316 23112
rect 9956 23196 10008 23248
rect 14924 23196 14976 23248
rect 9864 23128 9916 23180
rect 10876 23171 10928 23180
rect 10876 23137 10885 23171
rect 10885 23137 10919 23171
rect 10919 23137 10928 23171
rect 10876 23128 10928 23137
rect 11796 23128 11848 23180
rect 13360 23128 13412 23180
rect 16580 23264 16632 23316
rect 24584 23307 24636 23316
rect 24584 23273 24593 23307
rect 24593 23273 24627 23307
rect 24627 23273 24636 23307
rect 24584 23264 24636 23273
rect 16672 23196 16724 23248
rect 16856 23196 16908 23248
rect 2320 23035 2372 23044
rect 2320 23001 2329 23035
rect 2329 23001 2363 23035
rect 2363 23001 2372 23035
rect 2320 22992 2372 23001
rect 8116 22992 8168 23044
rect 10048 23060 10100 23112
rect 10692 23060 10744 23112
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 12072 23060 12124 23112
rect 12348 23060 12400 23112
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15568 23103 15620 23112
rect 15568 23069 15577 23103
rect 15577 23069 15611 23103
rect 15611 23069 15620 23103
rect 15568 23060 15620 23069
rect 18144 23128 18196 23180
rect 20812 23196 20864 23248
rect 21180 23196 21232 23248
rect 20352 23128 20404 23180
rect 22836 23171 22888 23180
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 24952 23196 25004 23248
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 16672 23060 16724 23112
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 20168 23060 20220 23112
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 10324 22992 10376 23044
rect 13544 22992 13596 23044
rect 16948 23035 17000 23044
rect 16948 23001 16957 23035
rect 16957 23001 16991 23035
rect 16991 23001 17000 23035
rect 16948 22992 17000 23001
rect 17040 23035 17092 23044
rect 17040 23001 17049 23035
rect 17049 23001 17083 23035
rect 17083 23001 17092 23035
rect 17040 22992 17092 23001
rect 21272 22992 21324 23044
rect 22284 23035 22336 23044
rect 22284 23001 22293 23035
rect 22293 23001 22327 23035
rect 22327 23001 22336 23035
rect 22284 22992 22336 23001
rect 7748 22967 7800 22976
rect 7748 22933 7757 22967
rect 7757 22933 7791 22967
rect 7791 22933 7800 22967
rect 7748 22924 7800 22933
rect 12348 22924 12400 22976
rect 12808 22924 12860 22976
rect 16856 22924 16908 22976
rect 17132 22924 17184 22976
rect 19432 22924 19484 22976
rect 21640 22967 21692 22976
rect 21640 22933 21649 22967
rect 21649 22933 21683 22967
rect 21683 22933 21692 22967
rect 21640 22924 21692 22933
rect 22744 22924 22796 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 6736 22720 6788 22772
rect 11060 22720 11112 22772
rect 11612 22720 11664 22772
rect 7748 22652 7800 22704
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 7288 22584 7340 22636
rect 7840 22584 7892 22636
rect 9496 22516 9548 22568
rect 10048 22584 10100 22636
rect 11060 22584 11112 22636
rect 11336 22584 11388 22636
rect 11428 22516 11480 22568
rect 16212 22720 16264 22772
rect 12164 22584 12216 22636
rect 15384 22652 15436 22704
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 18420 22652 18472 22704
rect 21088 22720 21140 22772
rect 21180 22720 21232 22772
rect 24032 22720 24084 22772
rect 19984 22652 20036 22704
rect 20904 22695 20956 22704
rect 20904 22661 20913 22695
rect 20913 22661 20947 22695
rect 20947 22661 20956 22695
rect 20904 22652 20956 22661
rect 23848 22652 23900 22704
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17868 22627 17920 22636
rect 17868 22593 17877 22627
rect 17877 22593 17911 22627
rect 17911 22593 17920 22627
rect 17868 22584 17920 22593
rect 25688 22652 25740 22704
rect 12256 22516 12308 22568
rect 14188 22516 14240 22568
rect 10140 22448 10192 22500
rect 10324 22491 10376 22500
rect 10324 22457 10333 22491
rect 10333 22457 10367 22491
rect 10367 22457 10376 22491
rect 10324 22448 10376 22457
rect 10416 22448 10468 22500
rect 16856 22448 16908 22500
rect 6000 22380 6052 22432
rect 8576 22380 8628 22432
rect 11060 22380 11112 22432
rect 12256 22380 12308 22432
rect 17316 22380 17368 22432
rect 18512 22516 18564 22568
rect 20812 22559 20864 22568
rect 19064 22448 19116 22500
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 20168 22448 20220 22500
rect 24768 22584 24820 22636
rect 38108 22652 38160 22704
rect 22100 22516 22152 22568
rect 23388 22516 23440 22568
rect 30196 22516 30248 22568
rect 20260 22380 20312 22432
rect 23480 22380 23532 22432
rect 28264 22380 28316 22432
rect 38016 22380 38068 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3792 22176 3844 22228
rect 11060 22176 11112 22228
rect 11428 22176 11480 22228
rect 12072 22176 12124 22228
rect 12256 22176 12308 22228
rect 17040 22176 17092 22228
rect 18144 22176 18196 22228
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 9220 22040 9272 22092
rect 9496 22108 9548 22160
rect 10324 22108 10376 22160
rect 12348 22151 12400 22160
rect 10140 22040 10192 22092
rect 12348 22117 12357 22151
rect 12357 22117 12391 22151
rect 12391 22117 12400 22151
rect 12348 22108 12400 22117
rect 15108 22108 15160 22160
rect 11060 22040 11112 22092
rect 12072 22040 12124 22092
rect 1584 21972 1636 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 8024 21972 8076 22024
rect 10324 21972 10376 22024
rect 10692 21972 10744 22024
rect 9404 21904 9456 21956
rect 10508 21904 10560 21956
rect 11612 21972 11664 22024
rect 12808 22040 12860 22092
rect 14924 22083 14976 22092
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 17592 22108 17644 22160
rect 18236 22040 18288 22092
rect 20260 22108 20312 22160
rect 6736 21879 6788 21888
rect 6736 21845 6745 21879
rect 6745 21845 6779 21879
rect 6779 21845 6788 21879
rect 6736 21836 6788 21845
rect 10600 21836 10652 21888
rect 15568 21947 15620 21956
rect 15568 21913 15577 21947
rect 15577 21913 15611 21947
rect 15611 21913 15620 21947
rect 15568 21904 15620 21913
rect 12624 21836 12676 21888
rect 13360 21836 13412 21888
rect 15200 21836 15252 21888
rect 16856 21947 16908 21956
rect 16856 21913 16865 21947
rect 16865 21913 16899 21947
rect 16899 21913 16908 21947
rect 17960 21947 18012 21956
rect 16856 21904 16908 21913
rect 17960 21913 17969 21947
rect 17969 21913 18003 21947
rect 18003 21913 18012 21947
rect 17960 21904 18012 21913
rect 18052 21947 18104 21956
rect 18052 21913 18061 21947
rect 18061 21913 18095 21947
rect 18095 21913 18104 21947
rect 18052 21904 18104 21913
rect 16028 21879 16080 21888
rect 16028 21845 16037 21879
rect 16037 21845 16071 21879
rect 16071 21845 16080 21879
rect 16028 21836 16080 21845
rect 17132 21836 17184 21888
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 38292 22015 38344 22024
rect 21456 21904 21508 21956
rect 22652 21904 22704 21956
rect 23480 21904 23532 21956
rect 23756 21904 23808 21956
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 9404 21632 9456 21684
rect 10416 21632 10468 21684
rect 10508 21632 10560 21684
rect 11152 21632 11204 21684
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 17960 21632 18012 21684
rect 21640 21632 21692 21684
rect 22652 21675 22704 21684
rect 22652 21641 22661 21675
rect 22661 21641 22695 21675
rect 22695 21641 22704 21675
rect 22652 21632 22704 21641
rect 6736 21564 6788 21616
rect 8484 21496 8536 21548
rect 8668 21496 8720 21548
rect 10508 21539 10560 21548
rect 10508 21505 10517 21539
rect 10517 21505 10551 21539
rect 10551 21505 10560 21539
rect 10508 21496 10560 21505
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 12348 21564 12400 21616
rect 14556 21607 14608 21616
rect 12072 21496 12124 21548
rect 13360 21496 13412 21548
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 5540 21360 5592 21412
rect 9220 21471 9272 21480
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 13176 21471 13228 21480
rect 12900 21360 12952 21412
rect 13176 21437 13185 21471
rect 13185 21437 13219 21471
rect 13219 21437 13228 21471
rect 13176 21428 13228 21437
rect 13084 21360 13136 21412
rect 14556 21573 14565 21607
rect 14565 21573 14599 21607
rect 14599 21573 14608 21607
rect 14556 21564 14608 21573
rect 16488 21564 16540 21616
rect 18696 21564 18748 21616
rect 16028 21496 16080 21548
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 20720 21564 20772 21616
rect 13452 21360 13504 21412
rect 13636 21360 13688 21412
rect 14004 21360 14056 21412
rect 19432 21496 19484 21548
rect 22100 21496 22152 21548
rect 24216 21564 24268 21616
rect 19248 21428 19300 21480
rect 19340 21428 19392 21480
rect 20812 21471 20864 21480
rect 20812 21437 20821 21471
rect 20821 21437 20855 21471
rect 20855 21437 20864 21471
rect 20812 21428 20864 21437
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 8484 21292 8536 21344
rect 9588 21292 9640 21344
rect 9680 21292 9732 21344
rect 10968 21292 11020 21344
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 12348 21335 12400 21344
rect 11060 21292 11112 21301
rect 12348 21301 12357 21335
rect 12357 21301 12391 21335
rect 12391 21301 12400 21335
rect 12348 21292 12400 21301
rect 22836 21360 22888 21412
rect 15568 21292 15620 21344
rect 19524 21292 19576 21344
rect 20260 21292 20312 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 9220 21088 9272 21140
rect 10784 21131 10836 21140
rect 10784 21097 10793 21131
rect 10793 21097 10827 21131
rect 10827 21097 10836 21131
rect 10784 21088 10836 21097
rect 11704 21131 11756 21140
rect 11704 21097 11713 21131
rect 11713 21097 11747 21131
rect 11747 21097 11756 21131
rect 11704 21088 11756 21097
rect 12348 21088 12400 21140
rect 16948 21088 17000 21140
rect 17960 21088 18012 21140
rect 20996 21088 21048 21140
rect 23020 21088 23072 21140
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 8024 21020 8076 21072
rect 8300 21020 8352 21072
rect 7104 20952 7156 21004
rect 7380 20884 7432 20936
rect 7840 20884 7892 20936
rect 8576 20927 8628 20936
rect 8576 20893 8585 20927
rect 8585 20893 8619 20927
rect 8619 20893 8628 20927
rect 8576 20884 8628 20893
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 13084 21020 13136 21072
rect 11336 20952 11388 21004
rect 13176 20952 13228 21004
rect 13452 20995 13504 21004
rect 13452 20961 13461 20995
rect 13461 20961 13495 20995
rect 13495 20961 13504 20995
rect 13452 20952 13504 20961
rect 13728 20952 13780 21004
rect 10692 20884 10744 20936
rect 15568 20952 15620 21004
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 21272 20952 21324 21004
rect 21640 20952 21692 21004
rect 10508 20816 10560 20868
rect 13084 20859 13136 20868
rect 13084 20825 13093 20859
rect 13093 20825 13127 20859
rect 13127 20825 13136 20859
rect 13084 20816 13136 20825
rect 7656 20748 7708 20800
rect 9404 20748 9456 20800
rect 10416 20748 10468 20800
rect 12164 20748 12216 20800
rect 12900 20748 12952 20800
rect 13360 20748 13412 20800
rect 15200 20884 15252 20936
rect 15476 20884 15528 20936
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 19432 20884 19484 20936
rect 20168 20884 20220 20936
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 22560 20884 22612 20936
rect 25044 20884 25096 20936
rect 38016 20927 38068 20936
rect 38016 20893 38025 20927
rect 38025 20893 38059 20927
rect 38059 20893 38068 20927
rect 38016 20884 38068 20893
rect 16764 20748 16816 20800
rect 19524 20748 19576 20800
rect 20168 20748 20220 20800
rect 24032 20748 24084 20800
rect 38200 20791 38252 20800
rect 38200 20757 38209 20791
rect 38209 20757 38243 20791
rect 38243 20757 38252 20791
rect 38200 20748 38252 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5540 20544 5592 20596
rect 8300 20544 8352 20596
rect 13084 20544 13136 20596
rect 13176 20544 13228 20596
rect 1584 20408 1636 20460
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 7656 20408 7708 20460
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 10324 20408 10376 20460
rect 9036 20340 9088 20392
rect 9404 20340 9456 20392
rect 11336 20408 11388 20460
rect 11520 20476 11572 20528
rect 11888 20519 11940 20528
rect 11888 20485 11897 20519
rect 11897 20485 11931 20519
rect 11931 20485 11940 20519
rect 11888 20476 11940 20485
rect 12992 20476 13044 20528
rect 16120 20476 16172 20528
rect 18880 20476 18932 20528
rect 20812 20544 20864 20596
rect 25044 20587 25096 20596
rect 25044 20553 25053 20587
rect 25053 20553 25087 20587
rect 25087 20553 25096 20587
rect 25044 20544 25096 20553
rect 20352 20519 20404 20528
rect 20352 20485 20361 20519
rect 20361 20485 20395 20519
rect 20395 20485 20404 20519
rect 20352 20476 20404 20485
rect 22836 20519 22888 20528
rect 22836 20485 22845 20519
rect 22845 20485 22879 20519
rect 22879 20485 22888 20519
rect 22836 20476 22888 20485
rect 24032 20519 24084 20528
rect 24032 20485 24041 20519
rect 24041 20485 24075 20519
rect 24075 20485 24084 20519
rect 24032 20476 24084 20485
rect 7104 20204 7156 20256
rect 10876 20204 10928 20256
rect 11888 20340 11940 20392
rect 15476 20408 15528 20460
rect 16764 20408 16816 20460
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 24584 20408 24636 20460
rect 11152 20272 11204 20324
rect 13360 20383 13412 20392
rect 12900 20272 12952 20324
rect 12992 20272 13044 20324
rect 13360 20349 13369 20383
rect 13369 20349 13403 20383
rect 13403 20349 13412 20383
rect 13360 20340 13412 20349
rect 13636 20340 13688 20392
rect 13728 20340 13780 20392
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 17224 20340 17276 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 22744 20383 22796 20392
rect 22744 20349 22753 20383
rect 22753 20349 22787 20383
rect 22787 20349 22796 20383
rect 22744 20340 22796 20349
rect 23940 20383 23992 20392
rect 23940 20349 23949 20383
rect 23949 20349 23983 20383
rect 23983 20349 23992 20383
rect 23940 20340 23992 20349
rect 17592 20272 17644 20324
rect 19340 20272 19392 20324
rect 13636 20204 13688 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 18236 20204 18288 20256
rect 22560 20272 22612 20324
rect 24492 20315 24544 20324
rect 24492 20281 24501 20315
rect 24501 20281 24535 20315
rect 24535 20281 24544 20315
rect 24492 20272 24544 20281
rect 26332 20204 26384 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7932 20000 7984 20052
rect 6460 19932 6512 19984
rect 7104 19864 7156 19916
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 7196 19796 7248 19848
rect 9220 19864 9272 19916
rect 10324 19864 10376 19916
rect 10784 19932 10836 19984
rect 10968 20000 11020 20052
rect 13360 20000 13412 20052
rect 13820 20000 13872 20052
rect 17224 20000 17276 20052
rect 20352 20000 20404 20052
rect 21272 20000 21324 20052
rect 21548 20043 21600 20052
rect 21548 20009 21557 20043
rect 21557 20009 21591 20043
rect 21591 20009 21600 20043
rect 21548 20000 21600 20009
rect 22836 20000 22888 20052
rect 13176 19932 13228 19984
rect 13268 19932 13320 19984
rect 10876 19864 10928 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 20260 19932 20312 19984
rect 17592 19864 17644 19916
rect 21364 19864 21416 19916
rect 8300 19796 8352 19848
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 11244 19796 11296 19848
rect 11520 19728 11572 19780
rect 12256 19796 12308 19848
rect 12716 19796 12768 19848
rect 13544 19796 13596 19848
rect 14832 19796 14884 19848
rect 9680 19660 9732 19712
rect 11060 19660 11112 19712
rect 12440 19660 12492 19712
rect 13636 19728 13688 19780
rect 17132 19796 17184 19848
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 18880 19796 18932 19848
rect 20904 19796 20956 19848
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 22744 19932 22796 19984
rect 22468 19864 22520 19916
rect 22284 19839 22336 19848
rect 13544 19660 13596 19712
rect 17868 19728 17920 19780
rect 18420 19728 18472 19780
rect 19984 19728 20036 19780
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 23204 19839 23256 19848
rect 23204 19805 23213 19839
rect 23213 19805 23247 19839
rect 23247 19805 23256 19839
rect 23204 19796 23256 19805
rect 23480 19796 23532 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 23296 19728 23348 19780
rect 16948 19660 17000 19712
rect 17684 19660 17736 19712
rect 22100 19660 22152 19712
rect 28264 19660 28316 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 8576 19456 8628 19508
rect 10968 19456 11020 19508
rect 11060 19456 11112 19508
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 8300 19320 8352 19372
rect 9128 19320 9180 19372
rect 9864 19320 9916 19372
rect 9864 19184 9916 19236
rect 11704 19388 11756 19440
rect 10416 19320 10468 19372
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 12808 19456 12860 19508
rect 13084 19456 13136 19508
rect 15568 19456 15620 19508
rect 10600 19252 10652 19304
rect 11980 19295 12032 19304
rect 11980 19261 11989 19295
rect 11989 19261 12023 19295
rect 12023 19261 12032 19295
rect 11980 19252 12032 19261
rect 12072 19252 12124 19304
rect 12440 19252 12492 19304
rect 14832 19388 14884 19440
rect 18328 19456 18380 19508
rect 13176 19252 13228 19304
rect 15200 19320 15252 19372
rect 16488 19320 16540 19372
rect 19340 19388 19392 19440
rect 20536 19456 20588 19508
rect 21180 19456 21232 19508
rect 22744 19499 22796 19508
rect 22744 19465 22753 19499
rect 22753 19465 22787 19499
rect 22787 19465 22796 19499
rect 22744 19456 22796 19465
rect 23664 19456 23716 19508
rect 23940 19456 23992 19508
rect 18420 19363 18472 19372
rect 11152 19184 11204 19236
rect 15016 19184 15068 19236
rect 15292 19252 15344 19304
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19432 19320 19484 19372
rect 20076 19320 20128 19372
rect 20812 19320 20864 19372
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 23296 19320 23348 19372
rect 24492 19320 24544 19372
rect 30288 19320 30340 19372
rect 16120 19184 16172 19236
rect 22928 19252 22980 19304
rect 19984 19184 20036 19236
rect 20444 19184 20496 19236
rect 22192 19184 22244 19236
rect 8576 19116 8628 19168
rect 10048 19116 10100 19168
rect 11704 19116 11756 19168
rect 13176 19116 13228 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 13728 19116 13780 19168
rect 17316 19116 17368 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10048 18912 10100 18964
rect 9680 18844 9732 18896
rect 7196 18776 7248 18828
rect 10600 18844 10652 18896
rect 11796 18844 11848 18896
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 9864 18708 9916 18760
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10784 18776 10836 18828
rect 14372 18819 14424 18828
rect 14372 18785 14381 18819
rect 14381 18785 14415 18819
rect 14415 18785 14424 18819
rect 14372 18776 14424 18785
rect 11244 18683 11296 18692
rect 8116 18572 8168 18624
rect 10048 18572 10100 18624
rect 11244 18649 11253 18683
rect 11253 18649 11287 18683
rect 11287 18649 11296 18683
rect 11244 18640 11296 18649
rect 11520 18640 11572 18692
rect 14188 18708 14240 18760
rect 13728 18640 13780 18692
rect 15292 18708 15344 18760
rect 18144 18844 18196 18896
rect 20720 18912 20772 18964
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 23480 18955 23532 18964
rect 23480 18921 23489 18955
rect 23489 18921 23523 18955
rect 23523 18921 23532 18955
rect 23480 18912 23532 18921
rect 18328 18844 18380 18896
rect 19616 18844 19668 18896
rect 22284 18844 22336 18896
rect 17408 18683 17460 18692
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 13820 18572 13872 18624
rect 14556 18572 14608 18624
rect 16304 18572 16356 18624
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 19340 18776 19392 18828
rect 20812 18708 20864 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 23296 18708 23348 18760
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 23756 18708 23808 18760
rect 30288 18708 30340 18760
rect 18604 18640 18656 18692
rect 19616 18683 19668 18692
rect 19616 18649 19625 18683
rect 19625 18649 19659 18683
rect 19659 18649 19668 18683
rect 20168 18683 20220 18692
rect 19616 18640 19668 18649
rect 20168 18649 20177 18683
rect 20177 18649 20211 18683
rect 20211 18649 20220 18683
rect 20168 18640 20220 18649
rect 34796 18640 34848 18692
rect 20904 18572 20956 18624
rect 33048 18572 33100 18624
rect 38016 18572 38068 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 5816 18368 5868 18420
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 7380 18232 7432 18284
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 10784 18368 10836 18420
rect 10968 18368 11020 18420
rect 11796 18343 11848 18352
rect 11796 18309 11805 18343
rect 11805 18309 11839 18343
rect 11839 18309 11848 18343
rect 11796 18300 11848 18309
rect 12532 18368 12584 18420
rect 16304 18411 16356 18420
rect 16304 18377 16313 18411
rect 16313 18377 16347 18411
rect 16347 18377 16356 18411
rect 16304 18368 16356 18377
rect 18604 18411 18656 18420
rect 18604 18377 18613 18411
rect 18613 18377 18647 18411
rect 18647 18377 18656 18411
rect 18604 18368 18656 18377
rect 26240 18368 26292 18420
rect 20168 18300 20220 18352
rect 20996 18300 21048 18352
rect 22192 18343 22244 18352
rect 22192 18309 22201 18343
rect 22201 18309 22235 18343
rect 22235 18309 22244 18343
rect 22192 18300 22244 18309
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 13636 18232 13688 18284
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 18880 18232 18932 18284
rect 8392 18164 8444 18216
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 12072 18207 12124 18216
rect 12072 18173 12081 18207
rect 12081 18173 12115 18207
rect 12115 18173 12124 18207
rect 12072 18164 12124 18173
rect 12808 18164 12860 18216
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 13176 18164 13228 18216
rect 16764 18164 16816 18216
rect 19432 18207 19484 18216
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 11244 18028 11296 18080
rect 14004 18096 14056 18148
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 19432 18164 19484 18173
rect 20260 18164 20312 18216
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 23112 18207 23164 18216
rect 22100 18164 22152 18173
rect 23112 18173 23121 18207
rect 23121 18173 23155 18207
rect 23155 18173 23164 18207
rect 23112 18164 23164 18173
rect 12900 18028 12952 18080
rect 13176 18028 13228 18080
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 15752 18028 15804 18080
rect 23388 18028 23440 18080
rect 24124 18028 24176 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1860 17824 1912 17876
rect 9220 17756 9272 17808
rect 10508 17756 10560 17808
rect 11796 17756 11848 17808
rect 12532 17756 12584 17808
rect 14648 17756 14700 17808
rect 19432 17824 19484 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 22192 17824 22244 17876
rect 20812 17756 20864 17808
rect 22376 17756 22428 17808
rect 9680 17688 9732 17740
rect 7288 17620 7340 17672
rect 8392 17663 8444 17672
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 9220 17620 9272 17672
rect 8024 17552 8076 17604
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11152 17620 11204 17672
rect 16488 17731 16540 17740
rect 16488 17697 16497 17731
rect 16497 17697 16531 17731
rect 16531 17697 16540 17731
rect 16488 17688 16540 17697
rect 21916 17688 21968 17740
rect 22100 17688 22152 17740
rect 18236 17663 18288 17672
rect 8484 17484 8536 17536
rect 8944 17484 8996 17536
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 20536 17620 20588 17672
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 26332 17620 26384 17672
rect 12532 17484 12584 17536
rect 12808 17595 12860 17604
rect 12808 17561 12817 17595
rect 12817 17561 12851 17595
rect 12851 17561 12860 17595
rect 12808 17552 12860 17561
rect 13176 17552 13228 17604
rect 13452 17552 13504 17604
rect 14832 17595 14884 17604
rect 14832 17561 14841 17595
rect 14841 17561 14875 17595
rect 14875 17561 14884 17595
rect 14832 17552 14884 17561
rect 15108 17484 15160 17536
rect 15476 17552 15528 17604
rect 17224 17552 17276 17604
rect 18052 17484 18104 17536
rect 34520 17484 34572 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7932 17280 7984 17332
rect 7380 17212 7432 17264
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 8944 17144 8996 17153
rect 10324 17187 10376 17196
rect 7012 17076 7064 17128
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 13084 17280 13136 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 17408 17280 17460 17332
rect 16488 17212 16540 17264
rect 16764 17212 16816 17264
rect 11060 17144 11112 17196
rect 10876 17076 10928 17128
rect 11796 17076 11848 17128
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 14280 17076 14332 17128
rect 14924 17119 14976 17128
rect 10508 16940 10560 16992
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 17868 17076 17920 17128
rect 18972 17076 19024 17128
rect 18696 17008 18748 17060
rect 21088 17280 21140 17332
rect 22836 17280 22888 17332
rect 20996 17212 21048 17264
rect 19616 17144 19668 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 20812 17144 20864 17196
rect 38016 17187 38068 17196
rect 38016 17153 38025 17187
rect 38025 17153 38059 17187
rect 38059 17153 38068 17187
rect 38016 17144 38068 17153
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 15108 16940 15160 16992
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 18052 16940 18104 16992
rect 19892 17008 19944 17060
rect 22376 17008 22428 17060
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 22008 16940 22060 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 10324 16736 10376 16788
rect 15200 16736 15252 16788
rect 17408 16736 17460 16788
rect 18236 16736 18288 16788
rect 19524 16736 19576 16788
rect 9312 16532 9364 16584
rect 10416 16532 10468 16584
rect 11336 16668 11388 16720
rect 13544 16668 13596 16720
rect 12532 16600 12584 16652
rect 12992 16600 13044 16652
rect 14464 16643 14516 16652
rect 14464 16609 14473 16643
rect 14473 16609 14507 16643
rect 14507 16609 14516 16643
rect 14464 16600 14516 16609
rect 15108 16600 15160 16652
rect 17224 16600 17276 16652
rect 19248 16668 19300 16720
rect 11060 16532 11112 16584
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 12440 16532 12492 16584
rect 12716 16532 12768 16584
rect 15292 16532 15344 16584
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 23572 16600 23624 16652
rect 26240 16600 26292 16652
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 19616 16575 19668 16584
rect 19616 16541 19625 16575
rect 19625 16541 19659 16575
rect 19659 16541 19668 16575
rect 19616 16532 19668 16541
rect 10968 16464 11020 16516
rect 9956 16396 10008 16448
rect 10324 16396 10376 16448
rect 12808 16396 12860 16448
rect 15108 16439 15160 16448
rect 15108 16405 15117 16439
rect 15117 16405 15151 16439
rect 15151 16405 15160 16439
rect 15108 16396 15160 16405
rect 15384 16464 15436 16516
rect 20352 16532 20404 16584
rect 35808 16600 35860 16652
rect 16304 16396 16356 16448
rect 19892 16396 19944 16448
rect 33508 16396 33560 16448
rect 33692 16439 33744 16448
rect 33692 16405 33701 16439
rect 33701 16405 33735 16439
rect 33735 16405 33744 16439
rect 33692 16396 33744 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 9220 16192 9272 16244
rect 10600 16192 10652 16244
rect 10876 16192 10928 16244
rect 12808 16192 12860 16244
rect 15108 16192 15160 16244
rect 18328 16235 18380 16244
rect 14188 16167 14240 16176
rect 14188 16133 14197 16167
rect 14197 16133 14231 16167
rect 14231 16133 14240 16167
rect 15568 16167 15620 16176
rect 14188 16124 14240 16133
rect 15568 16133 15577 16167
rect 15577 16133 15611 16167
rect 15611 16133 15620 16167
rect 15568 16124 15620 16133
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 18972 16235 19024 16244
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 20536 16192 20588 16244
rect 33692 16192 33744 16244
rect 35808 16192 35860 16244
rect 5724 16056 5776 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9312 16056 9364 16108
rect 9864 16056 9916 16108
rect 11336 16056 11388 16108
rect 12348 16056 12400 16108
rect 16672 16056 16724 16108
rect 17316 16056 17368 16108
rect 18696 16124 18748 16176
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 22560 16056 22612 16108
rect 33508 16056 33560 16108
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 11704 15920 11756 15972
rect 13176 15988 13228 16040
rect 13268 15920 13320 15972
rect 14188 15920 14240 15972
rect 17408 15988 17460 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 9312 15852 9364 15904
rect 13912 15852 13964 15904
rect 18236 15852 18288 15904
rect 19616 15852 19668 15904
rect 33324 15852 33376 15904
rect 35348 15852 35400 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 10324 15648 10376 15700
rect 11428 15648 11480 15700
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 13544 15648 13596 15700
rect 13820 15648 13872 15700
rect 15476 15648 15528 15700
rect 18144 15648 18196 15700
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 9312 15512 9364 15521
rect 13176 15512 13228 15564
rect 15936 15512 15988 15564
rect 16764 15512 16816 15564
rect 16948 15512 17000 15564
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9956 15444 10008 15496
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 12624 15444 12676 15496
rect 14372 15444 14424 15496
rect 15292 15487 15344 15496
rect 12716 15376 12768 15428
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 16396 15487 16448 15496
rect 15660 15376 15712 15428
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 18236 15444 18288 15496
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 33048 15444 33100 15496
rect 17960 15419 18012 15428
rect 17960 15385 17969 15419
rect 17969 15385 18003 15419
rect 18003 15385 18012 15419
rect 17960 15376 18012 15385
rect 16028 15308 16080 15360
rect 38016 15308 38068 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 11152 15104 11204 15156
rect 12440 15104 12492 15156
rect 13268 15036 13320 15088
rect 14924 15104 14976 15156
rect 16120 15147 16172 15156
rect 16120 15113 16129 15147
rect 16129 15113 16163 15147
rect 16163 15113 16172 15147
rect 16120 15104 16172 15113
rect 17960 15147 18012 15156
rect 17960 15113 17969 15147
rect 17969 15113 18003 15147
rect 18003 15113 18012 15147
rect 17960 15104 18012 15113
rect 15568 15036 15620 15088
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 12716 14968 12768 15020
rect 13544 14968 13596 15020
rect 15476 14968 15528 15020
rect 16304 15011 16356 15020
rect 14740 14900 14792 14952
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 17500 14943 17552 14952
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 13728 14832 13780 14884
rect 15384 14832 15436 14884
rect 20352 14832 20404 14884
rect 18052 14764 18104 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 8852 14560 8904 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 14832 14560 14884 14612
rect 15476 14603 15528 14612
rect 15476 14569 15485 14603
rect 15485 14569 15519 14603
rect 15519 14569 15528 14603
rect 15476 14560 15528 14569
rect 15844 14560 15896 14612
rect 17684 14560 17736 14612
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 10232 14424 10284 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14740 14356 14792 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16672 14356 16724 14408
rect 18604 14424 18656 14476
rect 19248 14424 19300 14476
rect 28908 14424 28960 14476
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 34520 14356 34572 14408
rect 35348 14356 35400 14408
rect 37280 14220 37332 14272
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 14464 14016 14516 14068
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 17500 14016 17552 14068
rect 13912 13880 13964 13932
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 20444 13880 20496 13932
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 16396 13472 16448 13524
rect 7932 13311 7984 13320
rect 7932 13277 7941 13311
rect 7941 13277 7975 13311
rect 7975 13277 7984 13311
rect 7932 13268 7984 13277
rect 15200 13268 15252 13320
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 6920 12928 6972 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 13084 12792 13136 12844
rect 19064 12792 19116 12844
rect 23848 12792 23900 12844
rect 33324 12792 33376 12844
rect 38016 12835 38068 12844
rect 38016 12801 38025 12835
rect 38025 12801 38059 12835
rect 38059 12801 38068 12835
rect 38016 12792 38068 12801
rect 5448 12588 5500 12640
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 24676 12588 24728 12640
rect 35348 12631 35400 12640
rect 35348 12597 35357 12631
rect 35357 12597 35391 12631
rect 35391 12597 35400 12631
rect 35348 12588 35400 12597
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 16580 12180 16632 12232
rect 38108 12180 38160 12232
rect 18328 12044 18380 12096
rect 21916 12044 21968 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 13268 11772 13320 11824
rect 22376 11772 22428 11824
rect 5632 11704 5684 11756
rect 13452 11704 13504 11756
rect 37924 11704 37976 11756
rect 24400 11500 24452 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7564 11296 7616 11348
rect 38200 11271 38252 11280
rect 38200 11237 38209 11271
rect 38209 11237 38243 11271
rect 38243 11237 38252 11271
rect 38200 11228 38252 11237
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 20536 11092 20588 11144
rect 37280 11092 37332 11144
rect 21180 11024 21232 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 22008 10684 22060 10736
rect 11520 10616 11572 10668
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 17408 10616 17460 10668
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 11888 10412 11940 10464
rect 15292 10412 15344 10464
rect 20260 10412 20312 10464
rect 25596 10412 25648 10464
rect 28356 10412 28408 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 7932 10208 7984 10260
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 5448 10004 5500 10056
rect 12072 10004 12124 10056
rect 3976 9911 4028 9920
rect 3976 9877 3985 9911
rect 3985 9877 4019 9911
rect 4019 9877 4028 9911
rect 3976 9868 4028 9877
rect 9680 9868 9732 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 16948 9120 17000 9172
rect 21364 9120 21416 9172
rect 13176 8959 13228 8968
rect 13176 8925 13185 8959
rect 13185 8925 13219 8959
rect 13219 8925 13228 8959
rect 13176 8916 13228 8925
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 35348 8916 35400 8968
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 12808 8576 12860 8628
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 22376 8619 22428 8628
rect 22376 8585 22385 8619
rect 22385 8585 22419 8619
rect 22419 8585 22428 8619
rect 22376 8576 22428 8585
rect 12624 8508 12676 8560
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 2320 8372 2372 8424
rect 22008 8440 22060 8492
rect 24860 8440 24912 8492
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 6368 8032 6420 8084
rect 13636 8032 13688 8084
rect 24124 8032 24176 8084
rect 38108 8075 38160 8084
rect 38108 8041 38117 8075
rect 38117 8041 38151 8075
rect 38151 8041 38160 8075
rect 38108 8032 38160 8041
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 8300 7828 8352 7880
rect 14280 7828 14332 7880
rect 28632 7828 28684 7880
rect 34796 7828 34848 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 17132 7692 17184 7744
rect 37096 7692 37148 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 35808 7352 35860 7404
rect 22468 7148 22520 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 21456 6944 21508 6996
rect 25412 6740 25464 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 28908 6443 28960 6452
rect 28908 6409 28917 6443
rect 28917 6409 28951 6443
rect 28951 6409 28960 6443
rect 28908 6400 28960 6409
rect 12900 6332 12952 6384
rect 3976 6264 4028 6316
rect 4712 6264 4764 6316
rect 11152 6264 11204 6316
rect 30288 6264 30340 6316
rect 38108 6307 38160 6316
rect 38108 6273 38117 6307
rect 38117 6273 38151 6307
rect 38151 6273 38160 6307
rect 38108 6264 38160 6273
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 37280 6060 37332 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 9128 5856 9180 5908
rect 15016 5720 15068 5772
rect 17316 5720 17368 5772
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 21180 5695 21232 5704
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 23204 5652 23256 5704
rect 24676 5652 24728 5704
rect 32588 5652 32640 5704
rect 34520 5652 34572 5704
rect 37096 5695 37148 5704
rect 37096 5661 37105 5695
rect 37105 5661 37139 5695
rect 37139 5661 37148 5695
rect 37096 5652 37148 5661
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 9128 5516 9180 5568
rect 19432 5516 19484 5568
rect 23204 5516 23256 5568
rect 25872 5516 25924 5568
rect 37832 5516 37884 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1860 5287 1912 5296
rect 1860 5253 1869 5287
rect 1869 5253 1903 5287
rect 1903 5253 1912 5287
rect 1860 5244 1912 5253
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 18696 5176 18748 5228
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 25596 5176 25648 5228
rect 4620 4972 4672 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 14924 4972 14976 5024
rect 16856 4972 16908 5024
rect 22652 4972 22704 5024
rect 31668 4972 31720 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37924 4768 37976 4820
rect 28356 4564 28408 4616
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 33968 4428 34020 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4804 4088 4856 4140
rect 23112 4088 23164 4140
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 37464 3884 37516 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8300 3680 8352 3732
rect 34520 3680 34572 3732
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 38108 3476 38160 3528
rect 38016 3340 38068 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 35808 3136 35860 3188
rect 1308 2932 1360 2984
rect 4620 3000 4672 3052
rect 36912 3043 36964 3052
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 37832 3000 37884 3052
rect 20 2796 72 2848
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6368 2592 6420 2644
rect 9496 2592 9548 2644
rect 11152 2592 11204 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 24860 2592 24912 2644
rect 28632 2592 28684 2644
rect 32588 2592 32640 2644
rect 4712 2524 4764 2576
rect 3148 2456 3200 2508
rect 25412 2456 25464 2508
rect 30288 2524 30340 2576
rect 33968 2456 34020 2508
rect 2596 2388 2648 2440
rect 4528 2388 4580 2440
rect 5816 2388 5868 2440
rect 7104 2388 7156 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 10324 2388 10376 2440
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 13544 2388 13596 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 18052 2388 18104 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 21272 2388 21324 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 23204 2388 23256 2440
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 27068 2388 27120 2440
rect 29000 2388 29052 2440
rect 30288 2388 30340 2440
rect 31668 2388 31720 2440
rect 33508 2388 33560 2440
rect 34796 2388 34848 2440
rect 38016 2431 38068 2440
rect 38016 2397 38025 2431
rect 38025 2397 38059 2431
rect 38059 2397 38068 2431
rect 38016 2388 38068 2397
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 13176 2320 13228 2372
rect 9036 2252 9088 2304
rect 11612 2252 11664 2304
rect 14832 2252 14884 2304
rect 16764 2252 16816 2304
rect 19340 2252 19392 2304
rect 22560 2252 22612 2304
rect 23848 2252 23900 2304
rect 25780 2252 25832 2304
rect 31576 2252 31628 2304
rect 36084 2252 36136 2304
rect 39304 2252 39356 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 3344 39222 3556 39250
rect 32 37262 60 39200
rect 20 37256 72 37262
rect 20 37198 72 37204
rect 1320 35873 1348 39200
rect 3252 39114 3280 39200
rect 3344 39114 3372 39222
rect 3252 39086 3372 39114
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1596 37126 1624 37198
rect 3148 37188 3200 37194
rect 3148 37130 3200 37136
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 1596 36786 1624 37062
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1596 36242 1624 36722
rect 1584 36236 1636 36242
rect 1584 36178 1636 36184
rect 1306 35864 1362 35873
rect 1306 35799 1362 35808
rect 1596 35562 1624 36178
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1584 35556 1636 35562
rect 1584 35498 1636 35504
rect 1596 35154 1624 35498
rect 1584 35148 1636 35154
rect 1584 35090 1636 35096
rect 1400 33924 1452 33930
rect 1400 33866 1452 33872
rect 1412 24342 1440 33866
rect 1596 33522 1624 35090
rect 1964 34610 1992 35634
rect 2964 35624 3016 35630
rect 2964 35566 3016 35572
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 2700 34610 2728 34682
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 2688 34604 2740 34610
rect 2688 34546 2740 34552
rect 1964 33998 1992 34546
rect 1952 33992 2004 33998
rect 1952 33934 2004 33940
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1504 25702 1532 32846
rect 1596 32366 1624 33458
rect 1766 33416 1822 33425
rect 1766 33351 1822 33360
rect 1780 33114 1808 33351
rect 1768 33108 1820 33114
rect 1768 33050 1820 33056
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1596 31890 1624 32302
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1596 30258 1624 31826
rect 1872 31793 1900 31826
rect 1858 31784 1914 31793
rect 1858 31719 1914 31728
rect 1964 31482 1992 33934
rect 2136 33652 2188 33658
rect 2136 33594 2188 33600
rect 1952 31476 2004 31482
rect 1952 31418 2004 31424
rect 1860 31340 1912 31346
rect 1860 31282 1912 31288
rect 1872 30734 1900 31282
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 1860 30728 1912 30734
rect 1674 30696 1730 30705
rect 1860 30670 1912 30676
rect 1674 30631 1730 30640
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 29170 1624 30194
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1596 28014 1624 28494
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 27470 1624 27950
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 26908 1624 27406
rect 1688 27010 1716 30631
rect 1872 29646 1900 30670
rect 1952 30048 2004 30054
rect 1952 29990 2004 29996
rect 1860 29640 1912 29646
rect 1858 29608 1860 29617
rect 1912 29608 1914 29617
rect 1858 29543 1914 29552
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 1872 28626 1900 29242
rect 1860 28620 1912 28626
rect 1860 28562 1912 28568
rect 1860 28144 1912 28150
rect 1858 28112 1860 28121
rect 1912 28112 1914 28121
rect 1858 28047 1914 28056
rect 1858 27704 1914 27713
rect 1858 27639 1860 27648
rect 1912 27639 1914 27648
rect 1860 27610 1912 27616
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1780 27130 1808 27231
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1688 26982 1808 27010
rect 1676 26920 1728 26926
rect 1596 26880 1676 26908
rect 1596 26382 1624 26880
rect 1676 26862 1728 26868
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 25838 1624 26318
rect 1780 26234 1808 26982
rect 1688 26206 1808 26234
rect 1584 25832 1636 25838
rect 1584 25774 1636 25780
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1596 25362 1624 25774
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1688 23118 1716 26206
rect 1766 25256 1822 25265
rect 1766 25191 1822 25200
rect 1780 24818 1808 25191
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1676 23112 1728 23118
rect 1676 23054 1728 23060
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21146 1624 21966
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 1766 20496 1822 20505
rect 1584 20460 1636 20466
rect 1766 20431 1822 20440
rect 1584 20402 1636 20408
rect 1596 19514 1624 20402
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 19145 1808 19314
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 1872 17882 1900 27610
rect 1964 26994 1992 29990
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 2056 26234 2084 30738
rect 1964 26206 2084 26234
rect 1964 23730 1992 26206
rect 2148 23866 2176 33594
rect 2320 33584 2372 33590
rect 2318 33552 2320 33561
rect 2372 33552 2374 33561
rect 2318 33487 2374 33496
rect 2976 32978 3004 35566
rect 3056 34536 3108 34542
rect 3056 34478 3108 34484
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 2332 30802 2360 32846
rect 2412 32768 2464 32774
rect 2412 32710 2464 32716
rect 2320 30796 2372 30802
rect 2320 30738 2372 30744
rect 2228 30728 2280 30734
rect 2228 30670 2280 30676
rect 2240 29714 2268 30670
rect 2228 29708 2280 29714
rect 2228 29650 2280 29656
rect 2320 28960 2372 28966
rect 2318 28928 2320 28937
rect 2372 28928 2374 28937
rect 2318 28863 2374 28872
rect 2424 27985 2452 32710
rect 2872 32496 2924 32502
rect 2872 32438 2924 32444
rect 2688 32360 2740 32366
rect 2884 32337 2912 32438
rect 2688 32302 2740 32308
rect 2870 32328 2926 32337
rect 2596 32224 2648 32230
rect 2596 32166 2648 32172
rect 2608 28762 2636 32166
rect 2700 31346 2728 32302
rect 2870 32263 2926 32272
rect 3068 31482 3096 34478
rect 3160 33114 3188 37130
rect 3424 37120 3476 37126
rect 3424 37062 3476 37068
rect 3240 36712 3292 36718
rect 3240 36654 3292 36660
rect 3252 35442 3280 36654
rect 3332 35624 3384 35630
rect 3330 35592 3332 35601
rect 3384 35592 3386 35601
rect 3330 35527 3386 35536
rect 3252 35414 3372 35442
rect 3240 35148 3292 35154
rect 3240 35090 3292 35096
rect 3252 35057 3280 35090
rect 3238 35048 3294 35057
rect 3238 34983 3294 34992
rect 3344 34950 3372 35414
rect 3436 35154 3464 37062
rect 3528 35494 3556 39222
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 4066 38176 4122 38185
rect 4066 38111 4122 38120
rect 4080 37670 4108 38111
rect 4540 37738 4568 39200
rect 4528 37732 4580 37738
rect 4528 37674 4580 37680
rect 4068 37664 4120 37670
rect 4068 37606 4120 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4712 37324 4764 37330
rect 4712 37266 4764 37272
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3988 36786 4016 37198
rect 4436 36848 4488 36854
rect 4434 36816 4436 36825
rect 4488 36816 4490 36825
rect 3976 36780 4028 36786
rect 4434 36751 4490 36760
rect 3976 36722 4028 36728
rect 3608 36712 3660 36718
rect 3608 36654 3660 36660
rect 3620 36281 3648 36654
rect 3606 36272 3662 36281
rect 3606 36207 3662 36216
rect 3882 36272 3938 36281
rect 3988 36242 4016 36722
rect 4618 36544 4674 36553
rect 4214 36476 4522 36485
rect 4618 36479 4674 36488
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3882 36207 3938 36216
rect 3976 36236 4028 36242
rect 3896 36106 3924 36207
rect 3976 36178 4028 36184
rect 3884 36100 3936 36106
rect 3884 36042 3936 36048
rect 3516 35488 3568 35494
rect 3516 35430 3568 35436
rect 3988 35154 4016 36178
rect 4632 36106 4660 36479
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4724 35494 4752 37266
rect 4804 37188 4856 37194
rect 4804 37130 4856 37136
rect 4816 36009 4844 37130
rect 5724 37120 5776 37126
rect 5722 37088 5724 37097
rect 5776 37088 5778 37097
rect 5722 37023 5778 37032
rect 5736 36378 5764 37023
rect 5724 36372 5776 36378
rect 5724 36314 5776 36320
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 4896 36032 4948 36038
rect 4802 36000 4858 36009
rect 4896 35974 4948 35980
rect 4802 35935 4858 35944
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3424 35148 3476 35154
rect 3424 35090 3476 35096
rect 3976 35148 4028 35154
rect 3976 35090 4028 35096
rect 3332 34944 3384 34950
rect 3330 34912 3332 34921
rect 3384 34912 3386 34921
rect 3330 34847 3386 34856
rect 3988 34610 4016 35090
rect 4712 34672 4764 34678
rect 4712 34614 4764 34620
rect 3976 34604 4028 34610
rect 3976 34546 4028 34552
rect 3988 34066 4016 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4724 34066 4752 34614
rect 4908 34406 4936 35974
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 3976 34060 4028 34066
rect 3976 34002 4028 34008
rect 4712 34060 4764 34066
rect 4712 34002 4764 34008
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3252 32910 3280 33934
rect 3988 33522 4016 34002
rect 4160 33924 4212 33930
rect 4160 33866 4212 33872
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 4172 33402 4200 33866
rect 4528 33448 4580 33454
rect 4080 33374 4200 33402
rect 4526 33416 4528 33425
rect 4580 33416 4582 33425
rect 3332 32972 3384 32978
rect 3332 32914 3384 32920
rect 3148 32904 3200 32910
rect 3148 32846 3200 32852
rect 3240 32904 3292 32910
rect 3240 32846 3292 32852
rect 3056 31476 3108 31482
rect 2884 31436 3056 31464
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2884 28994 2912 31436
rect 3056 31418 3108 31424
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2792 28966 2912 28994
rect 2596 28756 2648 28762
rect 2596 28698 2648 28704
rect 2686 28112 2742 28121
rect 2686 28047 2742 28056
rect 2410 27976 2466 27985
rect 2410 27911 2466 27920
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2412 24948 2464 24954
rect 2412 24890 2464 24896
rect 2424 24410 2452 24890
rect 2516 24818 2544 25298
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2412 24404 2464 24410
rect 2412 24346 2464 24352
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1964 23118 1992 23666
rect 2608 23322 2636 26930
rect 2700 25158 2728 28047
rect 2688 25152 2740 25158
rect 2688 25094 2740 25100
rect 2792 23730 2820 28966
rect 2976 28370 3004 30534
rect 3160 28665 3188 32846
rect 3344 31754 3372 32914
rect 3792 32768 3844 32774
rect 3792 32710 3844 32716
rect 3516 32224 3568 32230
rect 3516 32166 3568 32172
rect 3252 31726 3372 31754
rect 3146 28656 3202 28665
rect 3146 28591 3202 28600
rect 2884 28342 3004 28370
rect 2884 26314 2912 28342
rect 2964 28076 3016 28082
rect 2964 28018 3016 28024
rect 2976 27554 3004 28018
rect 2976 27526 3096 27554
rect 2872 26308 2924 26314
rect 2872 26250 2924 26256
rect 3068 24410 3096 27526
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3160 27130 3188 27406
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3252 24206 3280 31726
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3332 29504 3384 29510
rect 3332 29446 3384 29452
rect 3344 24274 3372 29446
rect 3436 28490 3464 30126
rect 3424 28484 3476 28490
rect 3424 28426 3476 28432
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 3436 27033 3464 27270
rect 3422 27024 3478 27033
rect 3422 26959 3478 26968
rect 3528 24886 3556 32166
rect 3700 29708 3752 29714
rect 3700 29650 3752 29656
rect 3606 27568 3662 27577
rect 3606 27503 3662 27512
rect 3620 27062 3648 27503
rect 3608 27056 3660 27062
rect 3608 26998 3660 27004
rect 3606 26888 3662 26897
rect 3606 26823 3662 26832
rect 3620 26518 3648 26823
rect 3608 26512 3660 26518
rect 3608 26454 3660 26460
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3620 25430 3648 25774
rect 3608 25424 3660 25430
rect 3608 25366 3660 25372
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 3712 24206 3740 29650
rect 3804 29073 3832 32710
rect 4080 32586 4108 33374
rect 4526 33351 4582 33360
rect 4618 33280 4674 33289
rect 4214 33212 4522 33221
rect 4618 33215 4674 33224
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4252 32904 4304 32910
rect 4252 32846 4304 32852
rect 3988 32558 4108 32586
rect 4264 32570 4292 32846
rect 4252 32564 4304 32570
rect 3988 32026 4016 32558
rect 4252 32506 4304 32512
rect 4066 32328 4122 32337
rect 4066 32263 4122 32272
rect 3976 32020 4028 32026
rect 3976 31962 4028 31968
rect 3988 31929 4016 31962
rect 3974 31920 4030 31929
rect 3974 31855 4030 31864
rect 3976 31816 4028 31822
rect 4080 31804 4108 32263
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4526 31920 4582 31929
rect 4526 31855 4582 31864
rect 4028 31776 4108 31804
rect 3976 31758 4028 31764
rect 3884 30592 3936 30598
rect 3884 30534 3936 30540
rect 3790 29064 3846 29073
rect 3790 28999 3846 29008
rect 3790 28248 3846 28257
rect 3790 28183 3846 28192
rect 3804 28014 3832 28183
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3606 23896 3662 23905
rect 3606 23831 3662 23840
rect 3620 23798 3648 23831
rect 3608 23792 3660 23798
rect 3608 23734 3660 23740
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 2318 23080 2374 23089
rect 2318 23015 2320 23024
rect 2372 23015 2374 23024
rect 2320 22986 2372 22992
rect 3804 22234 3832 27950
rect 3896 26314 3924 30534
rect 3976 30184 4028 30190
rect 3976 30126 4028 30132
rect 3988 28257 4016 30126
rect 4080 29714 4108 31776
rect 4540 31414 4568 31855
rect 4632 31754 4660 33215
rect 4724 32910 4752 34002
rect 5000 33425 5028 36042
rect 5828 35834 5856 39200
rect 5908 37800 5960 37806
rect 5908 37742 5960 37748
rect 5920 37466 5948 37742
rect 6552 37732 6604 37738
rect 6552 37674 6604 37680
rect 7012 37732 7064 37738
rect 7012 37674 7064 37680
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 6000 37460 6052 37466
rect 6000 37402 6052 37408
rect 5816 35828 5868 35834
rect 5816 35770 5868 35776
rect 5908 35624 5960 35630
rect 5908 35566 5960 35572
rect 5080 35488 5132 35494
rect 5080 35430 5132 35436
rect 4986 33416 5042 33425
rect 4986 33351 5042 33360
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4712 32768 4764 32774
rect 4712 32710 4764 32716
rect 4620 31748 4672 31754
rect 4620 31690 4672 31696
rect 4528 31408 4580 31414
rect 4528 31350 4580 31356
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30920 4660 31078
rect 4540 30892 4660 30920
rect 4540 30433 4568 30892
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4526 30424 4582 30433
rect 4526 30359 4582 30368
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 4526 29608 4582 29617
rect 4526 29543 4528 29552
rect 4580 29543 4582 29552
rect 4528 29514 4580 29520
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 29306 4108 29446
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4080 29170 4108 29242
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4528 28756 4580 28762
rect 4528 28698 4580 28704
rect 4434 28656 4490 28665
rect 4434 28591 4490 28600
rect 4448 28558 4476 28591
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4342 28384 4398 28393
rect 3974 28248 4030 28257
rect 4264 28218 4292 28358
rect 4342 28319 4398 28328
rect 3974 28183 4030 28192
rect 4252 28212 4304 28218
rect 3988 27316 4016 28183
rect 4252 28154 4304 28160
rect 4356 28150 4384 28319
rect 4344 28144 4396 28150
rect 4344 28086 4396 28092
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 4080 27606 4108 28018
rect 4448 28014 4476 28494
rect 4540 28422 4568 28698
rect 4528 28416 4580 28422
rect 4528 28358 4580 28364
rect 4436 28008 4488 28014
rect 4436 27950 4488 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4632 27402 4660 30534
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 3988 27288 4108 27316
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 3884 26308 3936 26314
rect 3884 26250 3936 26256
rect 3988 25906 4016 26386
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3988 25498 4016 25638
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3974 25392 4030 25401
rect 3974 25327 4030 25336
rect 3988 25226 4016 25327
rect 3976 25220 4028 25226
rect 3976 25162 4028 25168
rect 4080 24818 4108 27288
rect 4618 27024 4674 27033
rect 4724 26994 4752 32710
rect 4804 32496 4856 32502
rect 4804 32438 4856 32444
rect 4816 32065 4844 32438
rect 4802 32056 4858 32065
rect 4802 31991 4858 32000
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4816 28150 4844 31758
rect 4908 30938 4936 32846
rect 5000 32434 5028 32914
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5000 31249 5028 31282
rect 4986 31240 5042 31249
rect 4986 31175 5042 31184
rect 4896 30932 4948 30938
rect 4896 30874 4948 30880
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 4908 29170 4936 30738
rect 4988 30592 5040 30598
rect 4988 30534 5040 30540
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4804 28008 4856 28014
rect 4804 27950 4856 27956
rect 4618 26959 4674 26968
rect 4712 26988 4764 26994
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4528 26240 4580 26246
rect 4528 26182 4580 26188
rect 4540 26042 4568 26182
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4632 25974 4660 26959
rect 4712 26930 4764 26936
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 4724 25702 4752 25978
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4066 24712 4122 24721
rect 4356 24682 4384 25230
rect 4724 24750 4752 25638
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4066 24647 4122 24656
rect 4344 24676 4396 24682
rect 4080 24410 4108 24647
rect 4344 24618 4396 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4816 24274 4844 27950
rect 4908 27606 4936 28970
rect 5000 28626 5028 30534
rect 5092 30161 5120 35430
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5552 34513 5580 34546
rect 5538 34504 5594 34513
rect 5538 34439 5594 34448
rect 5172 34400 5224 34406
rect 5172 34342 5224 34348
rect 5184 34082 5212 34342
rect 5184 34054 5396 34082
rect 5262 32736 5318 32745
rect 5262 32671 5318 32680
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5184 30705 5212 32234
rect 5170 30696 5226 30705
rect 5170 30631 5226 30640
rect 5172 30184 5224 30190
rect 5078 30152 5134 30161
rect 5172 30126 5224 30132
rect 5078 30087 5134 30096
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 4988 28484 5040 28490
rect 4988 28426 5040 28432
rect 4896 27600 4948 27606
rect 4896 27542 4948 27548
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 4908 24682 4936 27406
rect 5000 25786 5028 28426
rect 5092 25974 5120 29990
rect 5080 25968 5132 25974
rect 5080 25910 5132 25916
rect 5000 25758 5120 25786
rect 4988 25152 5040 25158
rect 5092 25129 5120 25758
rect 5184 25362 5212 30126
rect 5276 29238 5304 32671
rect 5368 31090 5396 34054
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5460 31226 5488 33594
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5552 32978 5580 33254
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5552 32026 5580 32914
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5632 32292 5684 32298
rect 5632 32234 5684 32240
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5644 31482 5672 32234
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5460 31198 5580 31226
rect 5368 31062 5488 31090
rect 5356 30932 5408 30938
rect 5356 30874 5408 30880
rect 5264 29232 5316 29238
rect 5264 29174 5316 29180
rect 5368 29084 5396 30874
rect 5460 30297 5488 31062
rect 5446 30288 5502 30297
rect 5446 30223 5502 30232
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 5276 29056 5396 29084
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 4988 25094 5040 25100
rect 5078 25120 5134 25129
rect 4896 24676 4948 24682
rect 4896 24618 4948 24624
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5000 23186 5028 25094
rect 5078 25055 5134 25064
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5092 24410 5120 24754
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5276 23118 5304 29056
rect 5460 28642 5488 29786
rect 5368 28614 5488 28642
rect 5552 28642 5580 31198
rect 5644 30734 5672 31282
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5644 30258 5672 30670
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5552 28614 5672 28642
rect 5368 27418 5396 28614
rect 5448 28552 5500 28558
rect 5500 28512 5580 28540
rect 5448 28494 5500 28500
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 27878 5488 28358
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5368 27390 5488 27418
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5368 27062 5396 27270
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 5460 25770 5488 27390
rect 5448 25764 5500 25770
rect 5448 25706 5500 25712
rect 5552 25498 5580 28512
rect 5644 26874 5672 28614
rect 5736 27062 5764 32710
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5828 31346 5856 32506
rect 5920 32298 5948 35566
rect 6012 34066 6040 37402
rect 6184 35624 6236 35630
rect 6184 35566 6236 35572
rect 6196 35222 6224 35566
rect 6368 35284 6420 35290
rect 6368 35226 6420 35232
rect 6184 35216 6236 35222
rect 6184 35158 6236 35164
rect 6092 34944 6144 34950
rect 6092 34886 6144 34892
rect 6000 34060 6052 34066
rect 6000 34002 6052 34008
rect 6104 32858 6132 34886
rect 6380 34406 6408 35226
rect 6564 34474 6592 37674
rect 7024 37330 7052 37674
rect 7012 37324 7064 37330
rect 7012 37266 7064 37272
rect 6736 37256 6788 37262
rect 6736 37198 6788 37204
rect 6748 36718 6776 37198
rect 7380 36916 7432 36922
rect 7380 36858 7432 36864
rect 7392 36718 7420 36858
rect 6736 36712 6788 36718
rect 6736 36654 6788 36660
rect 7288 36712 7340 36718
rect 7288 36654 7340 36660
rect 7380 36712 7432 36718
rect 7380 36654 7432 36660
rect 6748 36242 6776 36654
rect 6920 36644 6972 36650
rect 6920 36586 6972 36592
rect 6932 36258 6960 36586
rect 6932 36242 7052 36258
rect 6736 36236 6788 36242
rect 6932 36236 7064 36242
rect 6932 36230 7012 36236
rect 6736 36178 6788 36184
rect 7012 36178 7064 36184
rect 6748 35698 6776 36178
rect 7012 36100 7064 36106
rect 7012 36042 7064 36048
rect 7024 35737 7052 36042
rect 7300 36009 7328 36654
rect 7378 36408 7434 36417
rect 7378 36343 7434 36352
rect 7286 36000 7342 36009
rect 7286 35935 7342 35944
rect 7010 35728 7066 35737
rect 6736 35692 6788 35698
rect 7010 35663 7066 35672
rect 6736 35634 6788 35640
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6552 34468 6604 34474
rect 6552 34410 6604 34416
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6368 34060 6420 34066
rect 6368 34002 6420 34008
rect 6012 32830 6132 32858
rect 6012 32434 6040 32830
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 5908 32292 5960 32298
rect 5908 32234 5960 32240
rect 5816 31340 5868 31346
rect 5816 31282 5868 31288
rect 5908 31272 5960 31278
rect 5908 31214 5960 31220
rect 5920 30938 5948 31214
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 6104 30818 6132 32710
rect 6184 31748 6236 31754
rect 6184 31690 6236 31696
rect 5828 30790 6132 30818
rect 5828 28966 5856 30790
rect 6000 30728 6052 30734
rect 6000 30670 6052 30676
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5920 29714 5948 30126
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 5828 28014 5856 28562
rect 5920 28558 5948 29650
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5920 28082 5948 28494
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 5816 28008 5868 28014
rect 5816 27950 5868 27956
rect 5920 27538 5948 28018
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 5724 27056 5776 27062
rect 5724 26998 5776 27004
rect 5644 26846 5948 26874
rect 5724 26784 5776 26790
rect 5724 26726 5776 26732
rect 5736 26586 5764 26726
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5538 24848 5594 24857
rect 5538 24783 5540 24792
rect 5592 24783 5594 24792
rect 5540 24754 5592 24760
rect 5644 23866 5672 26250
rect 5828 25838 5856 26386
rect 5920 25974 5948 26846
rect 5908 25968 5960 25974
rect 5908 25910 5960 25916
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 5722 25528 5778 25537
rect 5722 25463 5778 25472
rect 5736 25294 5764 25463
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5828 24886 5856 25774
rect 5920 25294 5948 25910
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5816 24880 5868 24886
rect 5816 24822 5868 24828
rect 5920 24206 5948 25230
rect 6012 24410 6040 30670
rect 6092 30660 6144 30666
rect 6092 30602 6144 30608
rect 6104 26994 6132 30602
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 6196 26568 6224 31690
rect 6276 30932 6328 30938
rect 6276 30874 6328 30880
rect 6288 30258 6316 30874
rect 6276 30252 6328 30258
rect 6276 30194 6328 30200
rect 6104 26540 6224 26568
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 6104 23322 6132 26540
rect 6182 26480 6238 26489
rect 6182 26415 6238 26424
rect 6196 26382 6224 26415
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 6380 23254 6408 34002
rect 6552 33992 6604 33998
rect 6552 33934 6604 33940
rect 6564 33522 6592 33934
rect 6656 33930 6684 35226
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6734 34232 6790 34241
rect 6734 34167 6736 34176
rect 6788 34167 6790 34176
rect 6736 34138 6788 34144
rect 6840 33998 6868 34478
rect 6828 33992 6880 33998
rect 6828 33934 6880 33940
rect 6644 33924 6696 33930
rect 6644 33866 6696 33872
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 6564 33289 6592 33458
rect 6840 33454 6868 33934
rect 6932 33658 6960 34954
rect 7196 34604 7248 34610
rect 7196 34546 7248 34552
rect 6920 33652 6972 33658
rect 6920 33594 6972 33600
rect 7104 33516 7156 33522
rect 7104 33458 7156 33464
rect 6828 33448 6880 33454
rect 6828 33390 6880 33396
rect 6736 33312 6788 33318
rect 6550 33280 6606 33289
rect 6736 33254 6788 33260
rect 6550 33215 6606 33224
rect 6552 32972 6604 32978
rect 6552 32914 6604 32920
rect 6460 32836 6512 32842
rect 6460 32778 6512 32784
rect 6472 32570 6500 32778
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 6564 32348 6592 32914
rect 6644 32360 6696 32366
rect 6564 32320 6644 32348
rect 6564 31278 6592 32320
rect 6644 32302 6696 32308
rect 6552 31272 6604 31278
rect 6552 31214 6604 31220
rect 6564 30190 6592 31214
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 6656 30394 6684 30670
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6552 30184 6604 30190
rect 6552 30126 6604 30132
rect 6748 27402 6776 33254
rect 6840 32978 6868 33390
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 7116 32502 7144 33458
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 6840 32337 6868 32370
rect 6826 32328 6882 32337
rect 6826 32263 6882 32272
rect 6920 32292 6972 32298
rect 6920 32234 6972 32240
rect 6932 31822 6960 32234
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7116 31686 7144 32438
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6840 31278 6868 31418
rect 7208 31278 7236 34546
rect 7392 33522 7420 36343
rect 7760 36242 7788 39200
rect 8484 37120 8536 37126
rect 8482 37088 8484 37097
rect 8536 37088 8538 37097
rect 8482 37023 8538 37032
rect 8850 37088 8906 37097
rect 8850 37023 8906 37032
rect 8666 36952 8722 36961
rect 8666 36887 8722 36896
rect 8680 36854 8708 36887
rect 8668 36848 8720 36854
rect 7944 36774 8616 36802
rect 8668 36790 8720 36796
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7748 36236 7800 36242
rect 7748 36178 7800 36184
rect 7380 33516 7432 33522
rect 7380 33458 7432 33464
rect 7380 32972 7432 32978
rect 7380 32914 7432 32920
rect 7392 32756 7420 32914
rect 7472 32768 7524 32774
rect 7392 32728 7472 32756
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 7196 31272 7248 31278
rect 7196 31214 7248 31220
rect 6920 31136 6972 31142
rect 6920 31078 6972 31084
rect 6828 30932 6880 30938
rect 6828 30874 6880 30880
rect 6840 30734 6868 30874
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28082 6868 28358
rect 6932 28150 6960 31078
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7196 30592 7248 30598
rect 7196 30534 7248 30540
rect 7116 29714 7144 30534
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 7104 29572 7156 29578
rect 7104 29514 7156 29520
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6840 27538 6868 28018
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6840 26994 6868 27474
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6550 26616 6606 26625
rect 6550 26551 6606 26560
rect 6564 24818 6592 26551
rect 6840 26450 6868 26930
rect 7024 26858 7052 29514
rect 7116 29170 7144 29514
rect 7208 29238 7236 30534
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7300 29050 7328 31826
rect 7392 31822 7420 32728
rect 7472 32710 7524 32716
rect 7380 31816 7432 31822
rect 7380 31758 7432 31764
rect 7472 31748 7524 31754
rect 7472 31690 7524 31696
rect 7380 30864 7432 30870
rect 7380 30806 7432 30812
rect 7392 29628 7420 30806
rect 7484 29753 7512 31690
rect 7470 29744 7526 29753
rect 7470 29679 7526 29688
rect 7392 29600 7512 29628
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7116 29022 7328 29050
rect 7012 26852 7064 26858
rect 7012 26794 7064 26800
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6840 26330 6868 26386
rect 6840 26302 6960 26330
rect 6932 25906 6960 26302
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6644 25220 6696 25226
rect 6644 25162 6696 25168
rect 6656 24818 6684 25162
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 7024 23730 7052 26794
rect 7116 26246 7144 29022
rect 7104 26240 7156 26246
rect 7104 26182 7156 26188
rect 7104 25832 7156 25838
rect 7392 25786 7420 29106
rect 7484 27470 7512 29600
rect 7576 28694 7604 36178
rect 7840 35624 7892 35630
rect 7840 35566 7892 35572
rect 7656 34672 7708 34678
rect 7656 34614 7708 34620
rect 7668 32502 7696 34614
rect 7852 33658 7880 35566
rect 7748 33652 7800 33658
rect 7748 33594 7800 33600
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7656 32496 7708 32502
rect 7656 32438 7708 32444
rect 7668 31890 7696 32438
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 7656 29640 7708 29646
rect 7760 29628 7788 33594
rect 7944 33538 7972 36774
rect 8024 36712 8076 36718
rect 8076 36660 8524 36666
rect 8024 36654 8524 36660
rect 8036 36638 8524 36654
rect 8588 36650 8616 36774
rect 8760 36712 8812 36718
rect 8758 36680 8760 36689
rect 8812 36680 8814 36689
rect 8300 36372 8352 36378
rect 8300 36314 8352 36320
rect 8312 36242 8340 36314
rect 8208 36236 8260 36242
rect 8208 36178 8260 36184
rect 8300 36236 8352 36242
rect 8300 36178 8352 36184
rect 8220 36122 8248 36178
rect 8392 36168 8444 36174
rect 8220 36106 8340 36122
rect 8392 36110 8444 36116
rect 8220 36100 8352 36106
rect 8220 36094 8300 36100
rect 8300 36042 8352 36048
rect 8404 35986 8432 36110
rect 8312 35958 8432 35986
rect 8024 35080 8076 35086
rect 8024 35022 8076 35028
rect 7708 29600 7788 29628
rect 7852 33510 7972 33538
rect 7656 29582 7708 29588
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 7668 28642 7696 29582
rect 7746 29200 7802 29209
rect 7746 29135 7802 29144
rect 7760 28762 7788 29135
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7576 27402 7604 28630
rect 7668 28614 7788 28642
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7668 27713 7696 27950
rect 7654 27704 7710 27713
rect 7654 27639 7710 27648
rect 7656 27464 7708 27470
rect 7656 27406 7708 27412
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 7104 25774 7156 25780
rect 7116 24750 7144 25774
rect 7208 25758 7420 25786
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7208 25498 7236 25758
rect 7286 25664 7342 25673
rect 7286 25599 7342 25608
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7300 23882 7328 25599
rect 7484 25498 7512 25774
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7208 23854 7328 23882
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 6748 22778 6776 23666
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 5552 20602 5580 21354
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6012 20466 6040 22374
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21622 6776 21830
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7116 21010 7144 21422
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 5828 18426 5856 19790
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 5736 16114 5764 18022
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1766 15736 1822 15745
rect 4214 15739 4522 15748
rect 1766 15671 1822 15680
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 1820 14376 1822 14385
rect 1766 14311 1822 14320
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1780 12345 1808 12786
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 5460 10062 5488 12582
rect 6472 12442 6500 19926
rect 7116 19922 7144 20198
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7208 19854 7236 23854
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7300 22030 7328 22578
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7392 20942 7420 25230
rect 7562 24712 7618 24721
rect 7562 24647 7618 24656
rect 7576 24206 7604 24647
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7668 22273 7696 27406
rect 7760 26246 7788 28614
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7748 24608 7800 24614
rect 7746 24576 7748 24585
rect 7800 24576 7802 24585
rect 7746 24511 7802 24520
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22710 7788 22918
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7852 22642 7880 33510
rect 8036 32756 8064 35022
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 8128 34134 8156 34478
rect 8116 34128 8168 34134
rect 8312 34105 8340 35958
rect 8392 35488 8444 35494
rect 8392 35430 8444 35436
rect 8404 35329 8432 35430
rect 8390 35320 8446 35329
rect 8390 35255 8446 35264
rect 8392 34944 8444 34950
rect 8392 34886 8444 34892
rect 8116 34070 8168 34076
rect 8298 34096 8354 34105
rect 8298 34031 8354 34040
rect 8208 33992 8260 33998
rect 8206 33960 8208 33969
rect 8260 33960 8262 33969
rect 8206 33895 8262 33904
rect 8404 33153 8432 34886
rect 8496 33930 8524 36638
rect 8576 36644 8628 36650
rect 8758 36615 8814 36624
rect 8576 36586 8628 36592
rect 8864 36242 8892 37023
rect 8942 36272 8998 36281
rect 8852 36236 8904 36242
rect 8942 36207 8998 36216
rect 8852 36178 8904 36184
rect 8956 36009 8984 36207
rect 8942 36000 8998 36009
rect 8942 35935 8998 35944
rect 8574 35728 8630 35737
rect 8574 35663 8630 35672
rect 8588 35630 8616 35663
rect 8576 35624 8628 35630
rect 8576 35566 8628 35572
rect 9048 34524 9076 39200
rect 9956 37324 10008 37330
rect 9956 37266 10008 37272
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9140 36718 9168 37198
rect 9586 36952 9642 36961
rect 9586 36887 9642 36896
rect 9600 36718 9628 36887
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9692 36718 9720 36790
rect 9128 36712 9180 36718
rect 9588 36712 9640 36718
rect 9128 36654 9180 36660
rect 9402 36680 9458 36689
rect 9140 36310 9168 36654
rect 9588 36654 9640 36660
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9402 36615 9458 36624
rect 9128 36304 9180 36310
rect 9128 36246 9180 36252
rect 9218 36272 9274 36281
rect 9140 35630 9168 36246
rect 9218 36207 9274 36216
rect 9232 36038 9260 36207
rect 9220 36032 9272 36038
rect 9220 35974 9272 35980
rect 9128 35624 9180 35630
rect 9128 35566 9180 35572
rect 9140 35154 9168 35566
rect 9416 35154 9444 36615
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9586 35728 9642 35737
rect 9586 35663 9642 35672
rect 9128 35148 9180 35154
rect 9128 35090 9180 35096
rect 9404 35148 9456 35154
rect 9404 35090 9456 35096
rect 9494 34912 9550 34921
rect 9494 34847 9550 34856
rect 9128 34536 9180 34542
rect 9048 34496 9128 34524
rect 9128 34478 9180 34484
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 9036 33924 9088 33930
rect 9036 33866 9088 33872
rect 8390 33144 8446 33153
rect 8390 33079 8446 33088
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8956 32910 8984 33050
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 8116 32768 8168 32774
rect 8036 32728 8116 32756
rect 8116 32710 8168 32716
rect 8392 32360 8444 32366
rect 8220 32320 8392 32348
rect 8114 32056 8170 32065
rect 8114 31991 8116 32000
rect 8168 31991 8170 32000
rect 8116 31962 8168 31968
rect 8220 31754 8248 32320
rect 8392 32302 8444 32308
rect 8496 31906 8524 32778
rect 8666 32328 8722 32337
rect 9048 32298 9076 33866
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 9416 33454 9444 33594
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 9404 33448 9456 33454
rect 9404 33390 9456 33396
rect 9220 32972 9272 32978
rect 9220 32914 9272 32920
rect 9232 32858 9260 32914
rect 9140 32830 9260 32858
rect 8666 32263 8722 32272
rect 9036 32292 9088 32298
rect 7932 31748 7984 31754
rect 7932 31690 7984 31696
rect 8036 31726 8248 31754
rect 8312 31878 8524 31906
rect 8576 31952 8628 31958
rect 8576 31894 8628 31900
rect 7944 29646 7972 31690
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 7944 28422 7972 29106
rect 7932 28416 7984 28422
rect 7932 28358 7984 28364
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7944 26353 7972 27406
rect 7930 26344 7986 26353
rect 7930 26279 7986 26288
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7654 22264 7710 22273
rect 7654 22199 7710 22208
rect 8036 22030 8064 31726
rect 8312 30054 8340 31878
rect 8588 31754 8616 31894
rect 8680 31822 8708 32263
rect 9036 32234 9088 32240
rect 8668 31816 8720 31822
rect 8668 31758 8720 31764
rect 9140 31754 9168 32830
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 9232 32337 9260 32710
rect 9218 32328 9274 32337
rect 9218 32263 9274 32272
rect 8496 31726 8616 31754
rect 8852 31748 8904 31754
rect 8496 31142 8524 31726
rect 8852 31690 8904 31696
rect 9048 31726 9168 31754
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8300 30048 8352 30054
rect 8206 30016 8262 30025
rect 8300 29990 8352 29996
rect 8206 29951 8262 29960
rect 8220 29578 8248 29951
rect 8208 29572 8260 29578
rect 8208 29514 8260 29520
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8220 28218 8248 28902
rect 8116 28212 8168 28218
rect 8116 28154 8168 28160
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8128 27470 8156 28154
rect 8312 27962 8340 29990
rect 8312 27934 8432 27962
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8298 24984 8354 24993
rect 8298 24919 8354 24928
rect 8312 23594 8340 24919
rect 8300 23588 8352 23594
rect 8300 23530 8352 23536
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8128 22098 8156 22986
rect 8116 22092 8168 22098
rect 8404 22094 8432 27934
rect 8496 24410 8524 31078
rect 8772 30190 8800 31214
rect 8760 30184 8812 30190
rect 8760 30126 8812 30132
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8680 29578 8708 29990
rect 8772 29646 8800 30126
rect 8760 29640 8812 29646
rect 8760 29582 8812 29588
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8588 29306 8616 29446
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8576 27940 8628 27946
rect 8576 27882 8628 27888
rect 8588 26926 8616 27882
rect 8680 27878 8708 29242
rect 8772 29238 8800 29582
rect 8760 29232 8812 29238
rect 8760 29174 8812 29180
rect 8758 29064 8814 29073
rect 8758 28999 8814 29008
rect 8668 27872 8720 27878
rect 8668 27814 8720 27820
rect 8680 27606 8708 27814
rect 8772 27674 8800 28999
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 8668 27600 8720 27606
rect 8668 27542 8720 27548
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8772 26790 8800 27610
rect 8864 27470 8892 31690
rect 8944 29572 8996 29578
rect 8944 29514 8996 29520
rect 8956 27985 8984 29514
rect 9048 28150 9076 31726
rect 9128 31476 9180 31482
rect 9128 31418 9180 31424
rect 9220 31476 9272 31482
rect 9220 31418 9272 31424
rect 9140 31385 9168 31418
rect 9126 31376 9182 31385
rect 9126 31311 9182 31320
rect 9128 29776 9180 29782
rect 9128 29718 9180 29724
rect 9140 29617 9168 29718
rect 9126 29608 9182 29617
rect 9126 29543 9182 29552
rect 9036 28144 9088 28150
rect 9036 28086 9088 28092
rect 8942 27976 8998 27985
rect 8942 27911 8998 27920
rect 8852 27464 8904 27470
rect 8852 27406 8904 27412
rect 8944 27396 8996 27402
rect 8944 27338 8996 27344
rect 8956 27062 8984 27338
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8850 26888 8906 26897
rect 8850 26823 8906 26832
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8864 24970 8892 26823
rect 8942 26208 8998 26217
rect 8942 26143 8998 26152
rect 8956 25974 8984 26143
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 9048 25158 9076 28086
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 9140 26994 9168 27474
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9126 25936 9182 25945
rect 9126 25871 9182 25880
rect 9036 25152 9088 25158
rect 9036 25094 9088 25100
rect 8864 24942 9076 24970
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8758 24440 8814 24449
rect 8484 24404 8536 24410
rect 8758 24375 8814 24384
rect 8484 24346 8536 24352
rect 8772 23730 8800 24375
rect 8864 24274 8892 24550
rect 8852 24268 8904 24274
rect 8852 24210 8904 24216
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8588 23610 8616 23666
rect 8588 23594 8800 23610
rect 8588 23588 8812 23594
rect 8588 23582 8760 23588
rect 8760 23530 8812 23536
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8404 22066 8524 22094
rect 8116 22034 8168 22040
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 20466 7696 20742
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7852 19938 7880 20878
rect 7944 20058 7972 21966
rect 8036 21078 8064 21966
rect 8496 21554 8524 22066
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8496 21350 8524 21490
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 8312 20602 8340 21014
rect 8588 20942 8616 22374
rect 8680 21554 8708 23462
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7852 19910 7972 19938
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7208 18834 7236 19790
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7944 18766 7972 19910
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8312 19378 8340 19790
rect 8588 19514 8616 20402
rect 9048 20398 9076 24942
rect 9140 21026 9168 25871
rect 9232 25294 9260 31418
rect 9324 30818 9352 33390
rect 9404 32904 9456 32910
rect 9402 32872 9404 32881
rect 9508 32892 9536 34847
rect 9600 34490 9628 35663
rect 9876 34490 9904 36110
rect 9968 35465 9996 37266
rect 10048 36848 10100 36854
rect 10048 36790 10100 36796
rect 10060 36145 10088 36790
rect 10336 36378 10364 39200
rect 11060 37800 11112 37806
rect 11060 37742 11112 37748
rect 11072 37466 11100 37742
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 12268 37346 12296 39200
rect 13268 37732 13320 37738
rect 13268 37674 13320 37680
rect 12268 37318 12572 37346
rect 11060 37256 11112 37262
rect 11060 37198 11112 37204
rect 12346 37224 12402 37233
rect 10600 37188 10652 37194
rect 10600 37130 10652 37136
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10046 36136 10102 36145
rect 10046 36071 10102 36080
rect 10416 35624 10468 35630
rect 10416 35566 10468 35572
rect 9954 35456 10010 35465
rect 9954 35391 10010 35400
rect 9600 34462 9720 34490
rect 9876 34462 10272 34490
rect 9588 34400 9640 34406
rect 9588 34342 9640 34348
rect 9692 34354 9720 34462
rect 10140 34400 10192 34406
rect 9600 33046 9628 34342
rect 9692 34326 9904 34354
rect 10140 34342 10192 34348
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9784 33697 9812 34002
rect 9770 33688 9826 33697
rect 9770 33623 9826 33632
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9588 33040 9640 33046
rect 9586 33008 9588 33017
rect 9680 33040 9732 33046
rect 9640 33008 9642 33017
rect 9680 32982 9732 32988
rect 9586 32943 9642 32952
rect 9456 32872 9458 32881
rect 9508 32864 9628 32892
rect 9402 32807 9458 32816
rect 9404 32768 9456 32774
rect 9402 32736 9404 32745
rect 9456 32736 9458 32745
rect 9402 32671 9458 32680
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9416 31754 9444 32234
rect 9496 31952 9548 31958
rect 9496 31894 9548 31900
rect 9404 31748 9456 31754
rect 9404 31690 9456 31696
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 9416 31278 9444 31418
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9324 30790 9444 30818
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 9324 27946 9352 30670
rect 9416 29345 9444 30790
rect 9402 29336 9458 29345
rect 9402 29271 9458 29280
rect 9312 27940 9364 27946
rect 9312 27882 9364 27888
rect 9404 27872 9456 27878
rect 9404 27814 9456 27820
rect 9416 27538 9444 27814
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9324 26194 9352 27338
rect 9416 26518 9444 27474
rect 9508 27010 9536 31894
rect 9600 30938 9628 32864
rect 9692 32434 9720 32982
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9692 31793 9720 32166
rect 9678 31784 9734 31793
rect 9678 31719 9734 31728
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 9600 30274 9628 30874
rect 9600 30246 9720 30274
rect 9588 29028 9640 29034
rect 9588 28970 9640 28976
rect 9692 28994 9720 30246
rect 9784 29617 9812 33254
rect 9876 32065 9904 34326
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 10060 33590 10088 34002
rect 10048 33584 10100 33590
rect 10048 33526 10100 33532
rect 9954 33280 10010 33289
rect 9954 33215 10010 33224
rect 9968 32910 9996 33215
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9956 32428 10008 32434
rect 9956 32370 10008 32376
rect 9862 32056 9918 32065
rect 9862 31991 9918 32000
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9876 29850 9904 31758
rect 9864 29844 9916 29850
rect 9864 29786 9916 29792
rect 9770 29608 9826 29617
rect 9770 29543 9826 29552
rect 9968 29458 9996 32370
rect 9784 29430 9996 29458
rect 9784 29102 9812 29430
rect 9954 29336 10010 29345
rect 9954 29271 10010 29280
rect 9968 29102 9996 29271
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 10060 28994 10088 33526
rect 10152 31822 10180 34342
rect 10244 32774 10272 34462
rect 10428 33674 10456 35566
rect 10506 35184 10562 35193
rect 10506 35119 10562 35128
rect 10520 35086 10548 35119
rect 10508 35080 10560 35086
rect 10612 35057 10640 37130
rect 11072 36718 11100 37198
rect 12346 37159 12402 37168
rect 12360 37126 12388 37159
rect 12348 37120 12400 37126
rect 12254 37088 12310 37097
rect 12544 37108 12572 37318
rect 12624 37120 12676 37126
rect 12544 37080 12624 37108
rect 12348 37062 12400 37068
rect 12624 37062 12676 37068
rect 12254 37023 12310 37032
rect 12164 36848 12216 36854
rect 11610 36816 11666 36825
rect 12164 36790 12216 36796
rect 11610 36751 11666 36760
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 10966 36544 11022 36553
rect 10966 36479 11022 36488
rect 10980 36106 11008 36479
rect 11072 36242 11100 36654
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11060 36236 11112 36242
rect 11060 36178 11112 36184
rect 10968 36100 11020 36106
rect 10968 36042 11020 36048
rect 10692 35760 10744 35766
rect 10692 35702 10744 35708
rect 10508 35022 10560 35028
rect 10598 35048 10654 35057
rect 10598 34983 10654 34992
rect 10508 34604 10560 34610
rect 10508 34546 10560 34552
rect 10336 33646 10456 33674
rect 10232 32768 10284 32774
rect 10232 32710 10284 32716
rect 10232 32224 10284 32230
rect 10232 32166 10284 32172
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10244 30802 10272 32166
rect 10232 30796 10284 30802
rect 10232 30738 10284 30744
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10138 30152 10194 30161
rect 10138 30087 10194 30096
rect 10152 30054 10180 30087
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10140 29844 10192 29850
rect 10140 29786 10192 29792
rect 10152 29306 10180 29786
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 9600 28762 9628 28970
rect 9692 28966 9812 28994
rect 10060 28966 10180 28994
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9692 27130 9720 28086
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9508 26982 9628 27010
rect 9600 26772 9628 26982
rect 9508 26744 9628 26772
rect 9404 26512 9456 26518
rect 9404 26454 9456 26460
rect 9508 26314 9536 26744
rect 9586 26616 9642 26625
rect 9586 26551 9642 26560
rect 9600 26518 9628 26551
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9324 26166 9628 26194
rect 9600 25294 9628 26166
rect 9784 25684 9812 28966
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9956 28960 10008 28966
rect 9956 28902 10008 28908
rect 9876 28801 9904 28902
rect 9862 28792 9918 28801
rect 9862 28727 9918 28736
rect 9968 28558 9996 28902
rect 10048 28620 10100 28626
rect 10048 28562 10100 28568
rect 9956 28552 10008 28558
rect 10060 28529 10088 28562
rect 9956 28494 10008 28500
rect 10046 28520 10102 28529
rect 10046 28455 10102 28464
rect 10048 28144 10100 28150
rect 10048 28086 10100 28092
rect 10060 27946 10088 28086
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 9956 25696 10008 25702
rect 9784 25656 9956 25684
rect 9956 25638 10008 25644
rect 9220 25288 9272 25294
rect 9588 25288 9640 25294
rect 9220 25230 9272 25236
rect 9310 25256 9366 25265
rect 9232 24818 9260 25230
rect 9588 25230 9640 25236
rect 9310 25191 9366 25200
rect 9956 25220 10008 25226
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 9232 22001 9260 22034
rect 9218 21992 9274 22001
rect 9218 21927 9274 21936
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9232 21146 9260 21422
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9140 20998 9260 21026
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9232 19922 9260 20998
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 9126 19408 9182 19417
rect 8300 19372 8352 19378
rect 9126 19343 9128 19352
rect 8300 19314 8352 19320
rect 9180 19343 9182 19352
rect 9128 19314 9180 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18766 8616 19110
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17678 7328 18022
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7392 17270 7420 18226
rect 7944 17338 7972 18702
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8128 18290 8156 18566
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8404 18057 8432 18158
rect 8390 18048 8446 18057
rect 8390 17983 8446 17992
rect 8404 17678 8432 17983
rect 9220 17808 9272 17814
rect 9220 17750 9272 17756
rect 9232 17678 9260 17750
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7024 15162 7052 17070
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 6932 12986 6960 14962
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 1780 9625 1808 9998
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7585 1808 7822
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 1858 5400 1914 5409
rect 1858 5335 1914 5344
rect 1872 5302 1900 5335
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 4865 1716 5170
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1320 800 1348 2926
rect 1780 2825 1808 3470
rect 2332 3194 2360 8366
rect 3988 6322 4016 9862
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1766 2816 1822 2825
rect 1766 2751 1822 2760
rect 3160 2514 3188 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3058 4660 4966
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2582 4752 6258
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 4146 4844 5510
rect 5644 5234 5672 11698
rect 6380 8090 6408 12174
rect 7576 11354 7604 14962
rect 8036 13530 8064 17546
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8496 17202 8524 17478
rect 8956 17202 8984 17478
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9232 16250 9260 17614
rect 9324 16590 9352 25191
rect 9956 25162 10008 25168
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9416 24342 9444 24754
rect 9404 24336 9456 24342
rect 9404 24278 9456 24284
rect 9508 23186 9536 24754
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9600 24449 9628 24618
rect 9862 24576 9918 24585
rect 9862 24511 9918 24520
rect 9586 24440 9642 24449
rect 9586 24375 9642 24384
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9508 22166 9536 22510
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9416 21690 9444 21898
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9692 21350 9720 24346
rect 9876 23186 9904 24511
rect 9968 24410 9996 25162
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10060 24138 10088 25094
rect 10152 24818 10180 28966
rect 10244 25158 10272 30194
rect 10336 30054 10364 33646
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10428 33289 10456 33458
rect 10414 33280 10470 33289
rect 10520 33266 10548 34546
rect 10598 33688 10654 33697
rect 10598 33623 10654 33632
rect 10612 33318 10640 33623
rect 10470 33238 10548 33266
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10414 33215 10470 33224
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 10428 32230 10456 32846
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10428 30841 10456 31758
rect 10520 31521 10548 33238
rect 10704 32570 10732 35702
rect 11072 35630 11100 36178
rect 11164 36145 11192 36518
rect 11150 36136 11206 36145
rect 11150 36071 11206 36080
rect 11428 36100 11480 36106
rect 11428 36042 11480 36048
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 10968 35556 11020 35562
rect 10968 35498 11020 35504
rect 10876 35488 10928 35494
rect 10874 35456 10876 35465
rect 10928 35456 10930 35465
rect 10874 35391 10930 35400
rect 10784 34944 10836 34950
rect 10784 34886 10836 34892
rect 10796 34202 10824 34886
rect 10876 34536 10928 34542
rect 10876 34478 10928 34484
rect 10784 34196 10836 34202
rect 10784 34138 10836 34144
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 32609 10824 33934
rect 10782 32600 10838 32609
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10692 32564 10744 32570
rect 10782 32535 10838 32544
rect 10692 32506 10744 32512
rect 10612 32366 10640 32506
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10600 32360 10652 32366
rect 10600 32302 10652 32308
rect 10796 32230 10824 32370
rect 10784 32224 10836 32230
rect 10784 32166 10836 32172
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10506 31512 10562 31521
rect 10506 31447 10562 31456
rect 10598 31376 10654 31385
rect 10598 31311 10654 31320
rect 10612 31278 10640 31311
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 10414 30832 10470 30841
rect 10414 30767 10470 30776
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10428 30122 10456 30534
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10520 29102 10548 30126
rect 10612 29345 10640 31214
rect 10704 30841 10732 31826
rect 10796 31754 10824 32166
rect 10784 31748 10836 31754
rect 10784 31690 10836 31696
rect 10796 31414 10824 31690
rect 10888 31482 10916 34478
rect 10980 34066 11008 35498
rect 11072 35086 11100 35566
rect 11152 35488 11204 35494
rect 11152 35430 11204 35436
rect 11164 35329 11192 35430
rect 11150 35320 11206 35329
rect 11150 35255 11206 35264
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 11072 34610 11100 35022
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 11164 34921 11192 34954
rect 11150 34912 11206 34921
rect 11150 34847 11206 34856
rect 11150 34776 11206 34785
rect 11150 34711 11206 34720
rect 11060 34604 11112 34610
rect 11060 34546 11112 34552
rect 11072 34066 11100 34546
rect 11164 34134 11192 34711
rect 11336 34536 11388 34542
rect 11336 34478 11388 34484
rect 11244 34468 11296 34474
rect 11244 34410 11296 34416
rect 11256 34377 11284 34410
rect 11242 34368 11298 34377
rect 11242 34303 11298 34312
rect 11152 34128 11204 34134
rect 11204 34088 11284 34116
rect 11152 34070 11204 34076
rect 10968 34060 11020 34066
rect 10968 34002 11020 34008
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 11072 33522 11100 34002
rect 10968 33516 11020 33522
rect 10968 33458 11020 33464
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10980 32434 11008 33458
rect 11072 32978 11100 33458
rect 11152 33380 11204 33386
rect 11152 33322 11204 33328
rect 11164 33046 11192 33322
rect 11152 33040 11204 33046
rect 11152 32982 11204 32988
rect 11060 32972 11112 32978
rect 11060 32914 11112 32920
rect 11072 32434 11100 32914
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 11072 31890 11100 32370
rect 11256 31906 11284 34088
rect 11060 31884 11112 31890
rect 11060 31826 11112 31832
rect 11164 31878 11284 31906
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10980 31482 11008 31622
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 10784 31408 10836 31414
rect 10784 31350 10836 31356
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10690 30832 10746 30841
rect 10690 30767 10746 30776
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 10692 30592 10744 30598
rect 10692 30534 10744 30540
rect 10598 29336 10654 29345
rect 10598 29271 10654 29280
rect 10600 29232 10652 29238
rect 10600 29174 10652 29180
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10508 29096 10560 29102
rect 10508 29038 10560 29044
rect 10336 28393 10364 29038
rect 10612 29034 10640 29174
rect 10600 29028 10652 29034
rect 10600 28970 10652 28976
rect 10704 28762 10732 30534
rect 10888 30433 10916 30602
rect 10874 30424 10930 30433
rect 10874 30359 10930 30368
rect 10980 30258 11008 31282
rect 11164 30734 11192 31878
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 10796 29238 10824 30194
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 10888 29646 10916 29786
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10784 29232 10836 29238
rect 10784 29174 10836 29180
rect 10796 28937 10824 29174
rect 10782 28928 10838 28937
rect 10782 28863 10838 28872
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10796 28642 10824 28698
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 10704 28614 10824 28642
rect 10888 28626 10916 29446
rect 10966 28792 11022 28801
rect 10966 28727 11022 28736
rect 10876 28620 10928 28626
rect 10322 28384 10378 28393
rect 10322 28319 10378 28328
rect 10428 28064 10456 28562
rect 10704 28506 10732 28614
rect 10876 28562 10928 28568
rect 10612 28490 10732 28506
rect 10600 28484 10732 28490
rect 10652 28478 10732 28484
rect 10784 28484 10836 28490
rect 10600 28426 10652 28432
rect 10784 28426 10836 28432
rect 10598 28384 10654 28393
rect 10598 28319 10654 28328
rect 10336 28036 10456 28064
rect 10336 27334 10364 28036
rect 10508 28008 10560 28014
rect 10508 27950 10560 27956
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10336 26081 10364 27270
rect 10322 26072 10378 26081
rect 10322 26007 10378 26016
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10140 24812 10192 24818
rect 10192 24772 10272 24800
rect 10140 24754 10192 24760
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9876 22001 9904 23122
rect 9862 21992 9918 22001
rect 9862 21927 9918 21936
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9600 20913 9628 21286
rect 9692 20942 9720 21286
rect 9680 20936 9732 20942
rect 9586 20904 9642 20913
rect 9680 20878 9732 20884
rect 9586 20839 9642 20848
rect 9404 20800 9456 20806
rect 9402 20768 9404 20777
rect 9456 20768 9458 20777
rect 9402 20703 9458 20712
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9416 18290 9444 20334
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9692 19145 9720 19654
rect 9876 19378 9904 20402
rect 9968 19854 9996 23190
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10060 22642 10088 23054
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 10060 19292 10088 22578
rect 10244 22522 10272 24772
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10152 22506 10272 22522
rect 10336 22506 10364 22986
rect 10428 22506 10456 24142
rect 10520 22545 10548 27950
rect 10612 24818 10640 28319
rect 10690 28248 10746 28257
rect 10796 28218 10824 28426
rect 10690 28183 10746 28192
rect 10784 28212 10836 28218
rect 10704 28082 10732 28183
rect 10784 28154 10836 28160
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10980 27674 11008 28727
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 11072 27402 11100 30670
rect 11164 30308 11192 30670
rect 11164 30280 11284 30308
rect 11152 29844 11204 29850
rect 11152 29786 11204 29792
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 11164 26897 11192 29786
rect 11256 28966 11284 30280
rect 11348 29850 11376 34478
rect 11440 34241 11468 36042
rect 11520 35284 11572 35290
rect 11520 35226 11572 35232
rect 11426 34232 11482 34241
rect 11426 34167 11482 34176
rect 11532 33658 11560 35226
rect 11624 34241 11652 36751
rect 11796 36644 11848 36650
rect 11796 36586 11848 36592
rect 11808 36530 11836 36586
rect 11808 36502 12112 36530
rect 12084 36378 12112 36502
rect 12072 36372 12124 36378
rect 12072 36314 12124 36320
rect 12176 36310 12204 36790
rect 12164 36304 12216 36310
rect 12164 36246 12216 36252
rect 12268 36009 12296 37023
rect 12346 36952 12402 36961
rect 12346 36887 12348 36896
rect 12400 36887 12402 36896
rect 12532 36916 12584 36922
rect 12348 36858 12400 36864
rect 12532 36858 12584 36864
rect 12544 36825 12572 36858
rect 12624 36848 12676 36854
rect 12530 36816 12586 36825
rect 12360 36774 12480 36802
rect 12360 36281 12388 36774
rect 12346 36272 12402 36281
rect 12346 36207 12402 36216
rect 12452 36174 12480 36774
rect 12624 36790 12676 36796
rect 12530 36751 12586 36760
rect 12636 36417 12664 36790
rect 12622 36408 12678 36417
rect 12622 36343 12678 36352
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 13174 36136 13230 36145
rect 12992 36100 13044 36106
rect 13174 36071 13230 36080
rect 12992 36042 13044 36048
rect 12440 36032 12492 36038
rect 11794 36000 11850 36009
rect 11794 35935 11850 35944
rect 12254 36000 12310 36009
rect 12440 35974 12492 35980
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12254 35935 12310 35944
rect 11702 34504 11758 34513
rect 11702 34439 11758 34448
rect 11610 34232 11666 34241
rect 11610 34167 11666 34176
rect 11610 33688 11666 33697
rect 11520 33652 11572 33658
rect 11610 33623 11666 33632
rect 11520 33594 11572 33600
rect 11518 33552 11574 33561
rect 11518 33487 11574 33496
rect 11532 33454 11560 33487
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11532 32502 11560 32914
rect 11520 32496 11572 32502
rect 11520 32438 11572 32444
rect 11624 31754 11652 33623
rect 11716 32337 11744 34439
rect 11808 32745 11836 35935
rect 12256 35828 12308 35834
rect 12256 35770 12308 35776
rect 12268 35737 12296 35770
rect 12254 35728 12310 35737
rect 12254 35663 12310 35672
rect 12072 35624 12124 35630
rect 11992 35572 12072 35578
rect 12452 35601 12480 35974
rect 12636 35737 12664 35974
rect 12622 35728 12678 35737
rect 12622 35663 12678 35672
rect 11992 35566 12124 35572
rect 12438 35592 12494 35601
rect 11992 35550 12112 35566
rect 11992 34542 12020 35550
rect 13004 35562 13032 36042
rect 13082 36000 13138 36009
rect 13082 35935 13138 35944
rect 12438 35527 12494 35536
rect 12992 35556 13044 35562
rect 12992 35498 13044 35504
rect 12808 35216 12860 35222
rect 12452 35164 12808 35170
rect 12452 35158 12860 35164
rect 12452 35142 12848 35158
rect 12072 34672 12124 34678
rect 12072 34614 12124 34620
rect 12084 34542 12112 34614
rect 12452 34542 12480 35142
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 12544 34649 12572 34954
rect 12530 34640 12586 34649
rect 12530 34575 12586 34584
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 12348 34400 12400 34406
rect 12348 34342 12400 34348
rect 12360 34066 12388 34342
rect 12438 34232 12494 34241
rect 12438 34167 12494 34176
rect 12348 34060 12400 34066
rect 12348 34002 12400 34008
rect 11888 33924 11940 33930
rect 11888 33866 11940 33872
rect 11900 33833 11928 33866
rect 11886 33824 11942 33833
rect 11886 33759 11942 33768
rect 12072 33448 12124 33454
rect 12072 33390 12124 33396
rect 12084 33318 12112 33390
rect 12072 33312 12124 33318
rect 12072 33254 12124 33260
rect 11794 32736 11850 32745
rect 11794 32671 11850 32680
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 11702 32328 11758 32337
rect 11702 32263 11758 32272
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11612 31748 11664 31754
rect 11532 31708 11612 31736
rect 11532 31226 11560 31708
rect 11612 31690 11664 31696
rect 11440 31198 11560 31226
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 11244 28960 11296 28966
rect 11244 28902 11296 28908
rect 11244 27668 11296 27674
rect 11244 27610 11296 27616
rect 11256 26926 11284 27610
rect 11244 26920 11296 26926
rect 11150 26888 11206 26897
rect 11244 26862 11296 26868
rect 11150 26823 11206 26832
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 10980 26586 11008 26726
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11256 26382 11284 26862
rect 11348 26518 11376 29038
rect 11440 28801 11468 31198
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11426 28792 11482 28801
rect 11426 28727 11482 28736
rect 11428 28688 11480 28694
rect 11428 28630 11480 28636
rect 11440 28257 11468 28630
rect 11426 28248 11482 28257
rect 11426 28183 11482 28192
rect 11532 27062 11560 30534
rect 11624 29646 11652 30806
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11716 29170 11744 31826
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11520 27056 11572 27062
rect 11520 26998 11572 27004
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 10966 25800 11022 25809
rect 10784 25764 10836 25770
rect 10784 25706 10836 25712
rect 10876 25764 10928 25770
rect 10966 25735 11022 25744
rect 10876 25706 10928 25712
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10704 23118 10732 24210
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10506 22536 10562 22545
rect 10140 22500 10272 22506
rect 10192 22494 10272 22500
rect 10140 22442 10192 22448
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 9968 19264 10088 19292
rect 10152 19281 10180 22034
rect 10138 19272 10194 19281
rect 9864 19236 9916 19242
rect 9968 19224 9996 19264
rect 9916 19196 9996 19224
rect 10138 19207 10194 19216
rect 9864 19178 9916 19184
rect 9678 19136 9734 19145
rect 9678 19071 9734 19080
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9692 17746 9720 18838
rect 9876 18766 9904 19178
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18970 10088 19110
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10046 18864 10102 18873
rect 10046 18799 10102 18808
rect 10060 18766 10088 18799
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9324 16114 9352 16526
rect 9876 16114 9904 18702
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18290 10088 18566
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 8864 14618 8892 16050
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15570 9352 15846
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9968 15502 9996 16390
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7944 10266 7972 13262
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 6380 2650 6408 5646
rect 8312 3738 8340 7822
rect 9140 5914 9168 15438
rect 10244 14482 10272 22494
rect 10324 22500 10376 22506
rect 10324 22442 10376 22448
rect 10416 22500 10468 22506
rect 10506 22471 10562 22480
rect 10416 22442 10468 22448
rect 10324 22160 10376 22166
rect 10322 22128 10324 22137
rect 10376 22128 10378 22137
rect 10322 22063 10378 22072
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10336 20890 10364 21966
rect 10428 21690 10456 22442
rect 10520 22080 10548 22471
rect 10520 22052 10640 22080
rect 10506 21992 10562 22001
rect 10506 21927 10508 21936
rect 10560 21927 10562 21936
rect 10508 21898 10560 21904
rect 10612 21894 10640 22052
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10520 21554 10548 21626
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10704 20942 10732 21966
rect 10796 21146 10824 25706
rect 10888 23186 10916 25706
rect 10980 24313 11008 25735
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10966 24304 11022 24313
rect 10966 24239 11022 24248
rect 11072 23322 11100 25230
rect 11164 24274 11192 25366
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22778 11100 23054
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11164 22658 11192 23666
rect 11072 22642 11192 22658
rect 11060 22636 11192 22642
rect 11112 22630 11192 22636
rect 11060 22578 11112 22584
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22234 11100 22374
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11058 22128 11114 22137
rect 11058 22063 11060 22072
rect 11112 22063 11114 22072
rect 11060 22034 11112 22040
rect 11256 21978 11284 25638
rect 11336 25288 11388 25294
rect 11624 25242 11652 28902
rect 11716 28529 11744 29106
rect 11702 28520 11758 28529
rect 11702 28455 11758 28464
rect 11716 28082 11744 28455
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11704 27940 11756 27946
rect 11704 27882 11756 27888
rect 11716 27674 11744 27882
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 11716 27402 11744 27610
rect 11704 27396 11756 27402
rect 11704 27338 11756 27344
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11716 25906 11744 27066
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11808 25294 11836 32166
rect 12070 31784 12126 31793
rect 12070 31719 12072 31728
rect 12124 31719 12126 31728
rect 12072 31690 12124 31696
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11992 30938 12020 31282
rect 12072 31204 12124 31210
rect 12072 31146 12124 31152
rect 11980 30932 12032 30938
rect 11980 30874 12032 30880
rect 11980 30796 12032 30802
rect 11980 30738 12032 30744
rect 11888 30728 11940 30734
rect 11888 30670 11940 30676
rect 11900 29578 11928 30670
rect 11992 30410 12020 30738
rect 12084 30598 12112 31146
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 12176 30410 12204 32506
rect 12346 32464 12402 32473
rect 12346 32399 12402 32408
rect 11992 30382 12204 30410
rect 12360 30394 12388 32399
rect 12452 30938 12480 34167
rect 12544 32230 12572 34478
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12636 33561 12664 33594
rect 12622 33552 12678 33561
rect 12622 33487 12678 33496
rect 12728 33454 12756 33798
rect 12716 33448 12768 33454
rect 12992 33448 13044 33454
rect 12716 33390 12768 33396
rect 12912 33408 12992 33436
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 31754 12756 32166
rect 12728 31726 12848 31754
rect 12624 31680 12676 31686
rect 12624 31622 12676 31628
rect 12530 31512 12586 31521
rect 12530 31447 12586 31456
rect 12544 31346 12572 31447
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12440 30932 12492 30938
rect 12636 30920 12664 31622
rect 12440 30874 12492 30880
rect 12544 30892 12664 30920
rect 12070 30016 12126 30025
rect 12070 29951 12126 29960
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11980 29572 12032 29578
rect 11980 29514 12032 29520
rect 11992 29073 12020 29514
rect 11978 29064 12034 29073
rect 11978 28999 12034 29008
rect 11980 28960 12032 28966
rect 11980 28902 12032 28908
rect 11992 28558 12020 28902
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11900 27062 11928 28358
rect 11992 28150 12020 28358
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 12084 26466 12112 29951
rect 12176 29850 12204 30382
rect 12348 30388 12400 30394
rect 12544 30376 12572 30892
rect 12820 30818 12848 31726
rect 12912 31278 12940 33408
rect 12992 33390 13044 33396
rect 13096 33266 13124 35935
rect 13188 34950 13216 36071
rect 13280 34950 13308 37674
rect 13556 37126 13584 39200
rect 13912 37460 13964 37466
rect 13912 37402 13964 37408
rect 13360 37120 13412 37126
rect 13360 37062 13412 37068
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 13372 36718 13400 37062
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 13360 36712 13412 36718
rect 13360 36654 13412 36660
rect 13176 34944 13228 34950
rect 13268 34944 13320 34950
rect 13176 34886 13228 34892
rect 13266 34912 13268 34921
rect 13320 34912 13322 34921
rect 13266 34847 13322 34856
rect 13174 34368 13230 34377
rect 13174 34303 13230 34312
rect 13188 33998 13216 34303
rect 13268 34196 13320 34202
rect 13268 34138 13320 34144
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13004 33238 13124 33266
rect 13004 31754 13032 33238
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 13084 31476 13136 31482
rect 13084 31418 13136 31424
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12348 30330 12400 30336
rect 12452 30348 12572 30376
rect 12636 30790 12848 30818
rect 12452 30122 12480 30348
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 12164 29844 12216 29850
rect 12164 29786 12216 29792
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 12268 29073 12296 29174
rect 12452 29102 12480 30058
rect 12544 29578 12572 30194
rect 12532 29572 12584 29578
rect 12532 29514 12584 29520
rect 12440 29096 12492 29102
rect 12254 29064 12310 29073
rect 12440 29038 12492 29044
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12254 28999 12310 29008
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 12360 28014 12388 28426
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12256 26852 12308 26858
rect 12256 26794 12308 26800
rect 12176 26625 12204 26794
rect 12162 26616 12218 26625
rect 12162 26551 12218 26560
rect 12268 26518 12296 26794
rect 11992 26438 12112 26466
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 11336 25230 11388 25236
rect 11348 24274 11376 25230
rect 11532 25214 11652 25242
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11348 23730 11376 24210
rect 11532 24070 11560 25214
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 22642 11376 23462
rect 11532 23322 11560 23530
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11440 22234 11468 22510
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11164 21950 11284 21978
rect 11164 21690 11192 21950
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 21350 11008 21490
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10692 20936 10744 20942
rect 10336 20874 10548 20890
rect 10692 20878 10744 20884
rect 10336 20868 10560 20874
rect 10336 20862 10508 20868
rect 10336 20466 10364 20862
rect 10508 20810 10560 20816
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10336 19224 10364 19858
rect 10428 19378 10456 20742
rect 10796 19990 10824 21082
rect 11072 20505 11100 21286
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11242 20768 11298 20777
rect 11242 20703 11298 20712
rect 11058 20496 11114 20505
rect 11058 20431 11114 20440
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10888 19922 10916 20198
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10980 19514 11008 19994
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19514 11100 19654
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10966 19408 11022 19417
rect 10416 19372 10468 19378
rect 10966 19343 10968 19352
rect 10416 19314 10468 19320
rect 11020 19343 11022 19352
rect 10968 19314 11020 19320
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10336 19196 10456 19224
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10336 16794 10364 17138
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10428 16590 10456 19196
rect 10612 18902 10640 19246
rect 11164 19242 11192 20266
rect 11256 19854 11284 20703
rect 11348 20466 11376 20946
rect 11532 20534 11560 23258
rect 11624 22778 11652 25094
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11716 23730 11744 24210
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11808 23186 11836 25094
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11900 23746 11928 24550
rect 11992 24290 12020 26438
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 12162 26344 12218 26353
rect 12084 25906 12112 26318
rect 12162 26279 12218 26288
rect 12176 26042 12204 26279
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12176 24954 12204 25842
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12256 24880 12308 24886
rect 12256 24822 12308 24828
rect 11992 24274 12204 24290
rect 11980 24268 12204 24274
rect 12032 24262 12204 24268
rect 11980 24210 12032 24216
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 11992 23866 12020 24074
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11900 23730 12020 23746
rect 11900 23724 12032 23730
rect 11900 23718 11980 23724
rect 11980 23666 12032 23672
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 12084 23118 12112 24074
rect 12176 23474 12204 24262
rect 12268 24206 12296 24822
rect 12360 24410 12388 27950
rect 12544 27010 12572 29038
rect 12452 26982 12572 27010
rect 12452 26625 12480 26982
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12438 26616 12494 26625
rect 12544 26586 12572 26862
rect 12438 26551 12494 26560
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12346 24304 12402 24313
rect 12346 24239 12402 24248
rect 12360 24206 12388 24239
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12360 23798 12388 24006
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12176 23446 12388 23474
rect 12162 23352 12218 23361
rect 12162 23287 12164 23296
rect 12216 23287 12218 23296
rect 12164 23258 12216 23264
rect 12360 23118 12388 23446
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12084 22098 12112 22170
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 11612 22024 11664 22030
rect 11610 21992 11612 22001
rect 11664 21992 11666 22001
rect 11610 21927 11666 21936
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11702 21448 11758 21457
rect 12084 21434 12112 21490
rect 11702 21383 11758 21392
rect 11992 21406 12112 21434
rect 11716 21146 11744 21383
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11900 20398 11928 20470
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11334 19272 11390 19281
rect 11152 19236 11204 19242
rect 11334 19207 11390 19216
rect 11152 19178 11204 19184
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10796 18426 10824 18770
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10520 17814 10548 18158
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10520 16998 10548 17750
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 15706 10364 16390
rect 10612 16250 10640 17614
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16250 10916 17070
rect 10980 16522 11008 18362
rect 11256 18086 11284 18634
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 16590 11100 17138
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 11164 15162 11192 17614
rect 11348 16726 11376 19207
rect 11532 18698 11560 19722
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11716 19174 11744 19382
rect 11992 19310 12020 21406
rect 12176 20806 12204 22578
rect 12256 22568 12308 22574
rect 12254 22536 12256 22545
rect 12308 22536 12310 22545
rect 12254 22471 12310 22480
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 22234 12296 22374
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12360 22166 12388 22918
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12254 21992 12310 22001
rect 12254 21927 12310 21936
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12268 19854 12296 21927
rect 12360 21622 12388 22102
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12360 21146 12388 21286
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19310 12480 19654
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11348 16114 11376 16662
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11440 15706 11468 16526
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 11532 10674 11560 18634
rect 11808 18358 11836 18838
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11808 17814 11836 18294
rect 12084 18222 12112 19246
rect 12544 18714 12572 25638
rect 12636 21894 12664 30790
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12728 29714 12756 29990
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12728 28218 12756 28494
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12728 23662 12756 27338
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12820 22982 12848 30670
rect 12912 29209 12940 31078
rect 12992 30864 13044 30870
rect 12992 30806 13044 30812
rect 13004 29782 13032 30806
rect 13096 30734 13124 31418
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12992 29776 13044 29782
rect 12992 29718 13044 29724
rect 13084 29776 13136 29782
rect 13084 29718 13136 29724
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 12898 29200 12954 29209
rect 12898 29135 12954 29144
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12912 28218 12940 28358
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 13004 27402 13032 29446
rect 12992 27396 13044 27402
rect 12992 27338 13044 27344
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12912 25906 12940 26726
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 13096 25673 13124 29718
rect 13188 29628 13216 33934
rect 13280 32774 13308 34138
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13280 29782 13308 32710
rect 13268 29776 13320 29782
rect 13268 29718 13320 29724
rect 13188 29600 13308 29628
rect 13174 29064 13230 29073
rect 13174 28999 13176 29008
rect 13228 28999 13230 29008
rect 13176 28970 13228 28976
rect 13176 27328 13228 27334
rect 13176 27270 13228 27276
rect 13188 26382 13216 27270
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 13082 25664 13138 25673
rect 13082 25599 13138 25608
rect 13188 25226 13216 26182
rect 13280 25702 13308 29600
rect 13372 25945 13400 36654
rect 13636 36576 13688 36582
rect 13634 36544 13636 36553
rect 13688 36544 13690 36553
rect 13634 36479 13690 36488
rect 13636 36168 13688 36174
rect 13636 36110 13688 36116
rect 13544 36032 13596 36038
rect 13544 35974 13596 35980
rect 13452 34944 13504 34950
rect 13452 34886 13504 34892
rect 13464 33930 13492 34886
rect 13556 34202 13584 35974
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13452 33924 13504 33930
rect 13452 33866 13504 33872
rect 13544 33380 13596 33386
rect 13544 33322 13596 33328
rect 13556 33289 13584 33322
rect 13542 33280 13598 33289
rect 13542 33215 13598 33224
rect 13648 31958 13676 36110
rect 13740 34785 13768 36790
rect 13726 34776 13782 34785
rect 13726 34711 13782 34720
rect 13924 34626 13952 37402
rect 15108 37256 15160 37262
rect 14370 37224 14426 37233
rect 15108 37198 15160 37204
rect 14370 37159 14426 37168
rect 14188 36712 14240 36718
rect 14188 36654 14240 36660
rect 14200 35154 14228 36654
rect 14280 36576 14332 36582
rect 14280 36518 14332 36524
rect 14292 36310 14320 36518
rect 14280 36304 14332 36310
rect 14280 36246 14332 36252
rect 14096 35148 14148 35154
rect 14096 35090 14148 35096
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 14002 34776 14058 34785
rect 14108 34746 14136 35090
rect 14278 35048 14334 35057
rect 14278 34983 14334 34992
rect 14002 34711 14004 34720
rect 14056 34711 14058 34720
rect 14096 34740 14148 34746
rect 14004 34682 14056 34688
rect 14096 34682 14148 34688
rect 13924 34598 14228 34626
rect 13728 34536 13780 34542
rect 13728 34478 13780 34484
rect 13740 33114 13768 34478
rect 14096 34400 14148 34406
rect 14096 34342 14148 34348
rect 14004 33924 14056 33930
rect 14004 33866 14056 33872
rect 14016 33658 14044 33866
rect 14108 33658 14136 34342
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 14096 33652 14148 33658
rect 14096 33594 14148 33600
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 13728 33108 13780 33114
rect 13728 33050 13780 33056
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13726 32736 13782 32745
rect 13726 32671 13782 32680
rect 13636 31952 13688 31958
rect 13636 31894 13688 31900
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13450 31376 13506 31385
rect 13450 31311 13452 31320
rect 13504 31311 13506 31320
rect 13452 31282 13504 31288
rect 13450 30424 13506 30433
rect 13450 30359 13506 30368
rect 13464 30326 13492 30359
rect 13452 30320 13504 30326
rect 13452 30262 13504 30268
rect 13450 27976 13506 27985
rect 13450 27911 13506 27920
rect 13358 25936 13414 25945
rect 13358 25871 13414 25880
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13096 24886 13124 25162
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13360 24336 13412 24342
rect 13360 24278 13412 24284
rect 13372 23730 13400 24278
rect 13464 24274 13492 27911
rect 13556 27674 13584 31758
rect 13636 31204 13688 31210
rect 13636 31146 13688 31152
rect 13648 28150 13676 31146
rect 13740 30938 13768 32671
rect 13832 32502 13860 33050
rect 13924 32842 13952 33458
rect 14016 33017 14044 33458
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 14002 33008 14058 33017
rect 14002 32943 14058 32952
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 13912 32836 13964 32842
rect 13912 32778 13964 32784
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13832 31278 13860 31758
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13832 30258 13860 31078
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13740 29646 13768 29990
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13728 27940 13780 27946
rect 13728 27882 13780 27888
rect 13544 27668 13596 27674
rect 13544 27610 13596 27616
rect 13740 26994 13768 27882
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13556 25362 13584 26182
rect 13648 25974 13676 26726
rect 13740 26382 13768 26930
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13636 25968 13688 25974
rect 13636 25910 13688 25916
rect 13832 25537 13860 29990
rect 13924 29170 13952 32778
rect 14016 32570 14044 32846
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 14016 30258 14044 31758
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14108 29238 14136 33254
rect 14200 32570 14228 34598
rect 14188 32564 14240 32570
rect 14188 32506 14240 32512
rect 14188 32292 14240 32298
rect 14188 32234 14240 32240
rect 14200 29866 14228 32234
rect 14292 31482 14320 34983
rect 14384 34490 14412 37159
rect 14830 36952 14886 36961
rect 14830 36887 14886 36896
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 14464 35692 14516 35698
rect 14464 35634 14516 35640
rect 14476 35476 14504 35634
rect 14556 35488 14608 35494
rect 14476 35448 14556 35476
rect 14556 35430 14608 35436
rect 14556 35012 14608 35018
rect 14556 34954 14608 34960
rect 14384 34462 14504 34490
rect 14372 34400 14424 34406
rect 14372 34342 14424 34348
rect 14384 34066 14412 34342
rect 14372 34060 14424 34066
rect 14372 34002 14424 34008
rect 14476 32774 14504 34462
rect 14372 32768 14424 32774
rect 14372 32710 14424 32716
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14384 32502 14412 32710
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14372 32496 14424 32502
rect 14372 32438 14424 32444
rect 14372 32360 14424 32366
rect 14370 32328 14372 32337
rect 14424 32328 14426 32337
rect 14370 32263 14426 32272
rect 14476 32042 14504 32506
rect 14568 32230 14596 34954
rect 14660 32570 14688 36110
rect 14740 36100 14792 36106
rect 14740 36042 14792 36048
rect 14752 35834 14780 36042
rect 14740 35828 14792 35834
rect 14740 35770 14792 35776
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14752 33522 14780 34546
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14752 32230 14780 33458
rect 14844 32842 14872 36887
rect 15120 35834 15148 37198
rect 15488 37126 15516 39200
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 16672 37256 16724 37262
rect 16672 37198 16724 37204
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15476 36644 15528 36650
rect 15476 36586 15528 36592
rect 15488 36378 15516 36586
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15384 36032 15436 36038
rect 15580 36009 15608 36722
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15384 35974 15436 35980
rect 15566 36000 15622 36009
rect 15108 35828 15160 35834
rect 15108 35770 15160 35776
rect 15292 35828 15344 35834
rect 15292 35770 15344 35776
rect 15304 35714 15332 35770
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 15120 35686 15332 35714
rect 15396 35698 15424 35974
rect 15566 35935 15622 35944
rect 15384 35692 15436 35698
rect 14832 32836 14884 32842
rect 14832 32778 14884 32784
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14740 32224 14792 32230
rect 14740 32166 14792 32172
rect 14476 32014 14596 32042
rect 14370 31920 14426 31929
rect 14370 31855 14372 31864
rect 14424 31855 14426 31864
rect 14372 31826 14424 31832
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30734 14320 31282
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14200 29838 14320 29866
rect 14188 29708 14240 29714
rect 14188 29650 14240 29656
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14200 29170 14228 29650
rect 14292 29306 14320 29838
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14476 29238 14504 29446
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 13912 29164 13964 29170
rect 13912 29106 13964 29112
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14280 29028 14332 29034
rect 14280 28970 14332 28976
rect 14096 28688 14148 28694
rect 14096 28630 14148 28636
rect 13912 27532 13964 27538
rect 13912 27474 13964 27480
rect 13924 26625 13952 27474
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 13910 26616 13966 26625
rect 13910 26551 13966 26560
rect 13818 25528 13874 25537
rect 13818 25463 13874 25472
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13450 24168 13506 24177
rect 13450 24103 13506 24112
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22098 12848 22918
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 12912 20806 12940 21354
rect 13096 21078 13124 21354
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 13188 21010 13216 21422
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13096 20602 13124 20810
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12992 20528 13044 20534
rect 13188 20482 13216 20538
rect 12992 20470 13044 20476
rect 13004 20330 13032 20470
rect 13096 20454 13216 20482
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 12716 19848 12768 19854
rect 12768 19808 12848 19836
rect 12716 19790 12768 19796
rect 12820 19514 12848 19808
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12820 18884 12848 19450
rect 12622 18864 12678 18873
rect 12622 18799 12678 18808
rect 12728 18856 12848 18884
rect 12452 18686 12572 18714
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11716 15706 11744 15914
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 9140 2446 9168 5510
rect 9508 2650 9536 8434
rect 9692 5710 9720 9862
rect 11808 6458 11836 17070
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 11164 2650 11192 6258
rect 11900 5234 11928 10406
rect 12084 10062 12112 18158
rect 12452 16590 12480 18686
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18426 12572 18566
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12544 17542 12572 17750
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12360 16017 12388 16050
rect 12346 16008 12402 16017
rect 12346 15943 12402 15952
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 15162 12480 15438
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12544 12434 12572 16594
rect 12636 15502 12664 18799
rect 12728 17354 12756 18856
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12820 17610 12848 18158
rect 12912 18086 12940 20266
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12728 17326 12940 17354
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12728 15434 12756 16526
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16250 12848 16390
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12912 16130 12940 17326
rect 13004 16658 13032 20266
rect 13096 19514 13124 20454
rect 13280 19990 13308 23598
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13372 23186 13400 23462
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 21554 13400 21830
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13464 21418 13492 24103
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 23050 13584 23666
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13542 22264 13598 22273
rect 13542 22199 13598 22208
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13358 20904 13414 20913
rect 13358 20839 13414 20848
rect 13372 20806 13400 20839
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 20058 13400 20334
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13188 19310 13216 19926
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13188 18222 13216 19110
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13096 17338 13124 18158
rect 13176 18080 13228 18086
rect 13464 18034 13492 20946
rect 13556 19854 13584 22199
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13648 20398 13676 21354
rect 13740 21010 13768 25162
rect 13924 24614 13952 26551
rect 14016 25906 14044 26794
rect 14108 25906 14136 28630
rect 14292 26994 14320 28970
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 27878 14412 28494
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14476 27470 14504 27950
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14568 27062 14596 32014
rect 14752 31346 14780 32166
rect 14936 31754 14964 35634
rect 15120 35494 15148 35686
rect 15384 35634 15436 35640
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 15488 35578 15516 35634
rect 15304 35550 15516 35578
rect 15108 35488 15160 35494
rect 15108 35430 15160 35436
rect 15014 34776 15070 34785
rect 15014 34711 15016 34720
rect 15068 34711 15070 34720
rect 15016 34682 15068 34688
rect 15304 34610 15332 35550
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15476 34604 15528 34610
rect 15476 34546 15528 34552
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 15120 34202 15148 34342
rect 15108 34196 15160 34202
rect 15108 34138 15160 34144
rect 15198 33824 15254 33833
rect 15304 33810 15332 34546
rect 15254 33782 15332 33810
rect 15198 33759 15254 33768
rect 15212 33522 15240 33759
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15212 33386 15240 33458
rect 15200 33380 15252 33386
rect 15200 33322 15252 33328
rect 15488 33046 15516 34546
rect 15672 33969 15700 36654
rect 15764 36378 15792 37198
rect 15844 37188 15896 37194
rect 15844 37130 15896 37136
rect 15856 36786 15884 37130
rect 16212 36916 16264 36922
rect 16212 36858 16264 36864
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15844 36168 15896 36174
rect 15844 36110 15896 36116
rect 15856 34134 15884 36110
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15948 35290 15976 35430
rect 15936 35284 15988 35290
rect 15936 35226 15988 35232
rect 16120 35080 16172 35086
rect 16120 35022 16172 35028
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15844 34128 15896 34134
rect 15844 34070 15896 34076
rect 15658 33960 15714 33969
rect 15658 33895 15714 33904
rect 15948 33697 15976 34886
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 15934 33688 15990 33697
rect 15844 33652 15896 33658
rect 16040 33658 16068 33934
rect 15934 33623 15990 33632
rect 16028 33652 16080 33658
rect 15844 33594 15896 33600
rect 16028 33594 16080 33600
rect 15856 33318 15884 33594
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15476 33040 15528 33046
rect 15476 32982 15528 32988
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 15028 32434 15056 32846
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15658 32600 15714 32609
rect 15658 32535 15714 32544
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15028 31822 15056 32370
rect 15396 32314 15424 32370
rect 15396 32298 15516 32314
rect 15396 32292 15528 32298
rect 15396 32286 15476 32292
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 14844 31726 14964 31754
rect 14740 31340 14792 31346
rect 14740 31282 14792 31288
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14660 28150 14688 28630
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14004 25220 14056 25226
rect 14004 25162 14056 25168
rect 14016 24750 14044 25162
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13648 19786 13676 20198
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13544 19712 13596 19718
rect 13740 19666 13768 20334
rect 13832 20262 13860 23802
rect 14016 21418 14044 24686
rect 14108 24206 14136 25638
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14200 24410 14228 24686
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14200 23730 14228 24006
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 20058 13860 20198
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13544 19654 13596 19660
rect 13556 19174 13584 19654
rect 13648 19638 13768 19666
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13648 18290 13676 19638
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 19009 13768 19110
rect 13726 19000 13782 19009
rect 13726 18935 13782 18944
rect 13740 18698 13768 18935
rect 14200 18766 14228 22510
rect 14292 20398 14320 26318
rect 14384 25362 14412 26386
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14476 25226 14504 26182
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14370 23216 14426 23225
rect 14370 23151 14426 23160
rect 14384 23118 14412 23151
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14384 19394 14412 23054
rect 14568 22148 14596 26862
rect 14660 26450 14688 27814
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14752 26353 14780 30670
rect 14844 27334 14872 31726
rect 15212 30870 15240 32166
rect 15396 31346 15424 32286
rect 15476 32234 15528 32240
rect 15672 32026 15700 32535
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15200 30864 15252 30870
rect 15200 30806 15252 30812
rect 15014 30288 15070 30297
rect 15014 30223 15070 30232
rect 15028 29646 15056 30223
rect 15108 29776 15160 29782
rect 15108 29718 15160 29724
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 15028 29322 15056 29582
rect 14936 29294 15056 29322
rect 14936 28082 14964 29294
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 15028 28558 15056 29106
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 14738 26344 14794 26353
rect 14738 26279 14794 26288
rect 14844 26194 14872 26862
rect 15028 26489 15056 28154
rect 15120 27402 15148 29718
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15212 28082 15240 28970
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15304 27674 15332 31078
rect 15566 30832 15622 30841
rect 15566 30767 15622 30776
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 15396 30258 15424 30534
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15488 27946 15516 28494
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15292 27668 15344 27674
rect 15292 27610 15344 27616
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15476 26920 15528 26926
rect 15474 26888 15476 26897
rect 15528 26888 15530 26897
rect 15474 26823 15530 26832
rect 15014 26480 15070 26489
rect 15014 26415 15070 26424
rect 15580 26382 15608 30767
rect 15856 30122 15884 32370
rect 15948 32026 15976 32778
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15856 29782 15884 30058
rect 15844 29776 15896 29782
rect 15844 29718 15896 29724
rect 15660 28416 15712 28422
rect 15660 28358 15712 28364
rect 15844 28416 15896 28422
rect 15844 28358 15896 28364
rect 15672 27538 15700 28358
rect 15856 28082 15884 28358
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 16040 28014 16068 32710
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15764 27062 15792 27814
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15672 26246 15700 26998
rect 14752 26166 14872 26194
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 14568 22120 14688 22148
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14568 21457 14596 21558
rect 14554 21448 14610 21457
rect 14554 21383 14610 21392
rect 14660 20262 14688 22120
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14292 19366 14412 19394
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13176 18022 13228 18028
rect 13188 17610 13216 18022
rect 13372 18006 13492 18034
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13372 17218 13400 18006
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13096 17190 13400 17218
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12820 16102 12940 16130
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12728 15026 12756 15370
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12544 12406 12664 12434
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12636 8566 12664 12406
rect 12820 8634 12848 16102
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12912 6390 12940 15982
rect 13096 12850 13124 17190
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 15570 13216 15982
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13280 15094 13308 15914
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13372 14906 13400 17070
rect 13280 14878 13400 14906
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13280 11830 13308 14878
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13464 11762 13492 17546
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13556 15706 13584 16662
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11716 2446 11744 4966
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 1465 1808 2246
rect 1766 1456 1822 1465
rect 1766 1391 1822 1400
rect 2608 800 2636 2382
rect 4540 800 4568 2382
rect 5828 800 5856 2382
rect 7116 800 7144 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 800 9076 2246
rect 10336 800 10364 2382
rect 13188 2378 13216 8910
rect 13648 8090 13676 18226
rect 13832 15706 13860 18566
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14016 17338 14044 18090
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14292 17134 14320 19366
rect 14370 19136 14426 19145
rect 14370 19071 14426 19080
rect 14384 18834 14412 19071
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18290 14596 18566
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14660 17814 14688 20198
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14370 16960 14426 16969
rect 14370 16895 14426 16904
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14200 15978 14228 16118
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14521 13768 14826
rect 13726 14512 13782 14521
rect 13726 14447 13782 14456
rect 13740 14414 13768 14447
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13924 13938 13952 15846
rect 14384 15502 14412 16895
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14476 14074 14504 16594
rect 14752 14958 14780 26166
rect 15566 26072 15622 26081
rect 15200 26036 15252 26042
rect 15566 26007 15622 26016
rect 15200 25978 15252 25984
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14844 24886 14872 25162
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 15028 23662 15056 23734
rect 15016 23656 15068 23662
rect 15016 23598 15068 23604
rect 14924 23248 14976 23254
rect 14924 23190 14976 23196
rect 14936 22098 14964 23190
rect 15120 22166 15148 25298
rect 15212 24750 15240 25978
rect 15292 25900 15344 25906
rect 15476 25900 15528 25906
rect 15344 25860 15424 25888
rect 15292 25842 15344 25848
rect 15396 25158 15424 25860
rect 15476 25842 15528 25848
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15304 23866 15332 24006
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15212 20942 15240 21830
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19446 14872 19790
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 15212 19378 15240 20878
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15304 19310 15332 23598
rect 15396 22710 15424 25094
rect 15488 23594 15516 25842
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15580 23118 15608 26007
rect 16132 25702 16160 35022
rect 16224 34542 16252 36858
rect 16580 36168 16632 36174
rect 16580 36110 16632 36116
rect 16304 36032 16356 36038
rect 16304 35974 16356 35980
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 16212 33924 16264 33930
rect 16212 33866 16264 33872
rect 16224 33658 16252 33866
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 16212 33380 16264 33386
rect 16212 33322 16264 33328
rect 16224 32570 16252 33322
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16316 30682 16344 35974
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16396 35080 16448 35086
rect 16396 35022 16448 35028
rect 16408 34610 16436 35022
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16408 33930 16436 34546
rect 16500 34474 16528 35634
rect 16592 35562 16620 36110
rect 16580 35556 16632 35562
rect 16580 35498 16632 35504
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16488 34128 16540 34134
rect 16488 34070 16540 34076
rect 16396 33924 16448 33930
rect 16396 33866 16448 33872
rect 16408 33266 16436 33866
rect 16500 33386 16528 34070
rect 16488 33380 16540 33386
rect 16488 33322 16540 33328
rect 16408 33238 16528 33266
rect 16500 32910 16528 33238
rect 16684 33046 16712 37198
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16764 36576 16816 36582
rect 16764 36518 16816 36524
rect 16776 36378 16804 36518
rect 16764 36372 16816 36378
rect 16764 36314 16816 36320
rect 16868 36310 16896 37198
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 16856 36304 16908 36310
rect 16856 36246 16908 36252
rect 17512 36174 17540 36722
rect 17592 36576 17644 36582
rect 17592 36518 17644 36524
rect 17604 36242 17632 36518
rect 17592 36236 17644 36242
rect 17592 36178 17644 36184
rect 17500 36168 17552 36174
rect 17130 36136 17186 36145
rect 17500 36110 17552 36116
rect 17130 36071 17132 36080
rect 17184 36071 17186 36080
rect 17132 36042 17184 36048
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16960 34678 16988 35430
rect 16948 34672 17000 34678
rect 16948 34614 17000 34620
rect 16948 34536 17000 34542
rect 16948 34478 17000 34484
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16672 33040 16724 33046
rect 16672 32982 16724 32988
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16396 32564 16448 32570
rect 16396 32506 16448 32512
rect 16408 31346 16436 32506
rect 16500 32298 16528 32846
rect 16488 32292 16540 32298
rect 16488 32234 16540 32240
rect 16868 32026 16896 34342
rect 16960 32978 16988 34478
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 16948 32768 17000 32774
rect 16948 32710 17000 32716
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16396 31340 16448 31346
rect 16396 31282 16448 31288
rect 16316 30654 16436 30682
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16316 29714 16344 30534
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16224 26382 16252 27406
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15948 24954 15976 25230
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16408 24834 16436 30654
rect 16960 30161 16988 32710
rect 17144 31482 17172 35770
rect 17512 35698 17540 36110
rect 17592 36032 17644 36038
rect 17592 35974 17644 35980
rect 17604 35766 17632 35974
rect 17592 35760 17644 35766
rect 17592 35702 17644 35708
rect 17500 35692 17552 35698
rect 17500 35634 17552 35640
rect 17512 34746 17540 35634
rect 17592 35488 17644 35494
rect 17592 35430 17644 35436
rect 17604 35193 17632 35430
rect 17590 35184 17646 35193
rect 17590 35119 17646 35128
rect 17868 35148 17920 35154
rect 17868 35090 17920 35096
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17592 34400 17644 34406
rect 17592 34342 17644 34348
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17328 33590 17356 33934
rect 17316 33584 17368 33590
rect 17316 33526 17368 33532
rect 17604 33454 17632 34342
rect 17592 33448 17644 33454
rect 17592 33390 17644 33396
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17512 32230 17540 32846
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17696 30326 17724 35022
rect 17880 34202 17908 35090
rect 17868 34196 17920 34202
rect 17868 34138 17920 34144
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17880 33590 17908 33798
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 18156 32842 18184 37062
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 18236 35624 18288 35630
rect 18236 35566 18288 35572
rect 18248 34746 18276 35566
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 18144 32836 18196 32842
rect 18144 32778 18196 32784
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17788 31754 17816 32370
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 31754 18092 32302
rect 17788 31726 17908 31754
rect 17684 30320 17736 30326
rect 17684 30262 17736 30268
rect 17880 30258 17908 31726
rect 17972 31726 18092 31754
rect 18432 31754 18460 35974
rect 19260 35873 19288 37198
rect 19352 36786 19380 37606
rect 19996 37126 20024 39200
rect 21284 37262 21312 39200
rect 22572 37262 22600 39200
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19246 35864 19302 35873
rect 19246 35799 19302 35808
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18616 33998 18644 34546
rect 19156 34128 19208 34134
rect 19156 34070 19208 34076
rect 18604 33992 18656 33998
rect 18604 33934 18656 33940
rect 18696 33856 18748 33862
rect 18696 33798 18748 33804
rect 18708 33114 18736 33798
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 18604 32292 18656 32298
rect 18604 32234 18656 32240
rect 18432 31726 18552 31754
rect 17972 31346 18000 31726
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 16946 30152 17002 30161
rect 16946 30087 17002 30096
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 17052 29170 17080 29446
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16776 28082 16804 28970
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16868 28121 16896 28494
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 16854 28112 16910 28121
rect 16764 28076 16816 28082
rect 16854 28047 16910 28056
rect 16764 28018 16816 28024
rect 16580 27872 16632 27878
rect 16580 27814 16632 27820
rect 16592 25498 16620 27814
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16672 27056 16724 27062
rect 16672 26998 16724 27004
rect 16684 26382 16712 26998
rect 16776 26858 16804 27270
rect 16764 26852 16816 26858
rect 16764 26794 16816 26800
rect 16762 26616 16818 26625
rect 16762 26551 16818 26560
rect 16776 26518 16804 26551
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16316 24806 16436 24834
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 16040 24138 16068 24550
rect 16316 24342 16344 24806
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16408 24342 16436 24686
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15474 22672 15530 22681
rect 15474 22607 15476 22616
rect 15528 22607 15530 22616
rect 15476 22578 15528 22584
rect 15488 20942 15516 22578
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15580 21350 15608 21898
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 16040 21554 16068 21830
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 16224 21010 16252 22714
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15474 20496 15530 20505
rect 15474 20431 15476 20440
rect 15528 20431 15530 20440
rect 15476 20402 15528 20408
rect 15580 19514 15608 20946
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 14414 14780 14894
rect 14844 14618 14872 17546
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14936 15162 14964 17070
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 2650 14320 7822
rect 15028 5778 15056 19178
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 16998 15148 17478
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15212 16794 15240 18022
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15120 16454 15148 16594
rect 15304 16590 15332 18702
rect 15764 18086 15792 20198
rect 16132 19922 16160 20470
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16250 15148 16390
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15304 14074 15332 15438
rect 15396 14890 15424 16458
rect 15488 15706 15516 17546
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15580 15094 15608 16118
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15488 14618 15516 14962
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15672 14414 15700 15370
rect 15856 14618 15884 18226
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15948 14074 15976 15506
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15198 13696 15254 13705
rect 15198 13631 15254 13640
rect 15212 13326 15240 13631
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 16040 10674 16068 15302
rect 16132 15162 16160 19178
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16316 18426 16344 18566
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16408 16574 16436 24278
rect 16592 24070 16620 25434
rect 17052 25294 17080 25774
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17144 24342 17172 28426
rect 17512 27878 17540 30194
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17696 28626 17724 30126
rect 17774 29744 17830 29753
rect 17774 29679 17830 29688
rect 17684 28620 17736 28626
rect 17684 28562 17736 28568
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17512 27130 17540 27814
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17328 26382 17356 26726
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17316 26240 17368 26246
rect 17316 26182 17368 26188
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17236 25362 17264 25706
rect 17328 25498 17356 26182
rect 17420 25906 17448 26930
rect 17590 26888 17646 26897
rect 17590 26823 17592 26832
rect 17644 26823 17646 26832
rect 17592 26794 17644 26800
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17512 25362 17540 26726
rect 17590 26072 17646 26081
rect 17590 26007 17646 26016
rect 17604 25906 17632 26007
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17512 24410 17540 24686
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16592 23322 16620 23598
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16684 23254 16712 24074
rect 16868 23254 16896 24142
rect 17144 23730 17172 24278
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16856 23248 16908 23254
rect 16856 23190 16908 23196
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16486 22808 16542 22817
rect 16486 22743 16542 22752
rect 16500 21622 16528 22743
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16500 17746 16528 19314
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16500 17270 16528 17682
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16408 16546 16620 16574
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16316 15026 16344 16390
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16408 13530 16436 15438
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16592 12238 16620 16546
rect 16684 16114 16712 23054
rect 16868 22982 16896 23190
rect 17052 23050 17080 23462
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16868 21962 16896 22442
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16960 21146 16988 22986
rect 17132 22976 17184 22982
rect 17052 22924 17132 22930
rect 17052 22918 17184 22924
rect 17052 22902 17172 22918
rect 17052 22642 17080 22902
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17052 22234 17080 22578
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 21690 17172 21830
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 20466 16804 20742
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 17236 20398 17264 23530
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17328 21554 17356 22374
rect 17604 22166 17632 25434
rect 17696 24682 17724 28562
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17788 24562 17816 29679
rect 17880 28694 17908 30194
rect 17868 28688 17920 28694
rect 17868 28630 17920 28636
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17880 25294 17908 27406
rect 17972 27033 18000 31282
rect 18236 30864 18288 30870
rect 18236 30806 18288 30812
rect 18248 30666 18276 30806
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18328 30660 18380 30666
rect 18328 30602 18380 30608
rect 18248 29186 18276 30602
rect 18340 30394 18368 30602
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18052 29164 18104 29170
rect 18248 29158 18368 29186
rect 18052 29106 18104 29112
rect 18064 28558 18092 29106
rect 18236 29028 18288 29034
rect 18236 28970 18288 28976
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18064 28150 18092 28494
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 17958 27024 18014 27033
rect 17958 26959 18014 26968
rect 18064 26382 18092 28086
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18156 25498 18184 27542
rect 18248 26926 18276 28970
rect 18340 26994 18368 29158
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18432 26586 18460 29038
rect 18524 28218 18552 31726
rect 18616 31414 18644 32234
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18892 31822 18920 32166
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18788 31272 18840 31278
rect 18788 31214 18840 31220
rect 18972 31272 19024 31278
rect 18972 31214 19024 31220
rect 18800 30938 18828 31214
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18984 30666 19012 31214
rect 19168 31210 19196 34070
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 19260 32910 19288 34002
rect 19352 33153 19380 36518
rect 19338 33144 19394 33153
rect 19338 33079 19394 33088
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19156 31204 19208 31210
rect 19156 31146 19208 31152
rect 18972 30660 19024 30666
rect 18972 30602 19024 30608
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18892 28762 18920 29582
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18512 28008 18564 28014
rect 18512 27950 18564 27956
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18340 26042 18368 26318
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17696 24534 17816 24562
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 17696 22094 17724 24534
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17788 23730 17816 24006
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17880 22642 17908 23462
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17696 22066 17908 22094
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17236 20058 17264 20334
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17604 19922 17632 20266
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16960 19310 16988 19654
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17270 16804 18158
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 14414 16712 16050
rect 16776 15570 16804 17206
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15304 5234 15332 10406
rect 16960 9178 16988 15506
rect 17038 13968 17094 13977
rect 17038 13903 17040 13912
rect 17092 13903 17094 13912
rect 17040 13874 17092 13880
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17144 7750 17172 19790
rect 17696 19718 17724 20878
rect 17880 19786 17908 22066
rect 18064 21962 18092 23802
rect 18156 23186 18184 24074
rect 18248 23730 18276 25638
rect 18524 24818 18552 27950
rect 18616 27538 18644 28358
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18708 27130 18736 27338
rect 18800 27130 18828 27406
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 18708 24818 18736 26454
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18892 24682 18920 25434
rect 18984 25226 19012 30602
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 19168 29306 19196 29582
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19076 26994 19104 27270
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19168 25906 19196 29242
rect 19260 27402 19288 29446
rect 19352 29238 19380 31826
rect 19444 30802 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20088 35222 20116 37198
rect 20628 37188 20680 37194
rect 20628 37130 20680 37136
rect 23940 37188 23992 37194
rect 23940 37130 23992 37136
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20166 36680 20222 36689
rect 20166 36615 20222 36624
rect 20076 35216 20128 35222
rect 20076 35158 20128 35164
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19984 33448 20036 33454
rect 19984 33390 20036 33396
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19524 32564 19576 32570
rect 19524 32506 19576 32512
rect 19536 31822 19564 32506
rect 19996 32026 20024 33390
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 20076 31952 20128 31958
rect 20076 31894 20128 31900
rect 19524 31816 19576 31822
rect 19524 31758 19576 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19628 30734 19656 31078
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 30326 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19444 29050 19472 30126
rect 19616 29776 19668 29782
rect 19522 29744 19578 29753
rect 19616 29718 19668 29724
rect 19522 29679 19524 29688
rect 19576 29679 19578 29688
rect 19524 29650 19576 29656
rect 19628 29617 19656 29718
rect 19800 29640 19852 29646
rect 19614 29608 19670 29617
rect 19800 29582 19852 29588
rect 19614 29543 19670 29552
rect 19812 29510 19840 29582
rect 19800 29504 19852 29510
rect 19800 29446 19852 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19522 29200 19578 29209
rect 19522 29135 19578 29144
rect 19352 29022 19472 29050
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19352 25294 19380 29022
rect 19536 28506 19564 29135
rect 19996 28626 20024 31418
rect 20088 31414 20116 31894
rect 20076 31408 20128 31414
rect 20076 31350 20128 31356
rect 20180 29594 20208 36615
rect 20364 33522 20392 37062
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20260 33312 20312 33318
rect 20260 33254 20312 33260
rect 20088 29566 20208 29594
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19444 28478 19564 28506
rect 19444 25974 19472 28478
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19628 27470 19656 27814
rect 19996 27606 20024 28562
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19536 26314 19564 26522
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19444 25294 19472 25910
rect 19996 25770 20024 26794
rect 19984 25764 20036 25770
rect 19984 25706 20036 25712
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 18972 25220 19024 25226
rect 18972 25162 19024 25168
rect 18880 24676 18932 24682
rect 18880 24618 18932 24624
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23866 18552 24006
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 18156 22234 18184 23122
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18432 22710 18460 23054
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18524 22574 18552 23802
rect 18512 22568 18564 22574
rect 18512 22510 18564 22516
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 17972 21690 18000 21898
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17972 21146 18000 21626
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18248 20262 18276 22034
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 18340 19514 18368 20402
rect 18708 19854 18736 21558
rect 18880 20528 18932 20534
rect 18880 20470 18932 20476
rect 18892 19854 18920 20470
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18432 19378 18460 19722
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17236 16658 17264 17546
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17328 16114 17356 19110
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17420 17338 17448 18634
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16794 17448 16934
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17328 5778 17356 14894
rect 17420 10674 17448 15982
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17512 14074 17540 14894
rect 17696 14618 17724 16594
rect 17880 14618 17908 17070
rect 18064 16998 18092 17478
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18156 15706 18184 18838
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18248 16794 18276 17614
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18340 16250 18368 18838
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 18616 18426 18644 18634
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18892 18290 18920 19790
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18694 17776 18750 17785
rect 18694 17711 18750 17720
rect 18708 17678 18736 17711
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17354 18736 17614
rect 18708 17326 18828 17354
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18708 16182 18736 17002
rect 18800 16590 18828 17326
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18984 16250 19012 17070
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18248 15502 18276 15846
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15162 18000 15370
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 18064 14414 18092 14758
rect 18616 14482 18644 14962
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 19076 12850 19104 22442
rect 19352 22094 19380 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 24342 19472 24754
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19432 24336 19484 24342
rect 19720 24313 19748 24346
rect 19432 24278 19484 24284
rect 19706 24304 19762 24313
rect 19444 22982 19472 24278
rect 19706 24239 19762 24248
rect 19720 24206 19748 24239
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22710 20024 24006
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19352 22066 19472 22094
rect 19444 21554 19472 22066
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19260 20210 19288 21422
rect 19352 20330 19380 21422
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19260 20182 19380 20210
rect 19352 19530 19380 20182
rect 19260 19502 19380 19530
rect 19260 18714 19288 19502
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19352 18834 19380 19382
rect 19444 19378 19472 20878
rect 19536 20806 19564 21286
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19996 19242 20024 19722
rect 20088 19378 20116 29566
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 29170 20208 29446
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 20272 28626 20300 33254
rect 20640 32570 20668 37130
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 21272 33380 21324 33386
rect 21272 33322 21324 33328
rect 21088 33040 21140 33046
rect 21088 32982 21140 32988
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20352 32224 20404 32230
rect 20352 32166 20404 32172
rect 20364 31754 20392 32166
rect 21100 31958 21128 32982
rect 21088 31952 21140 31958
rect 21088 31894 21140 31900
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20548 31754 20576 31826
rect 20352 31748 20404 31754
rect 20352 31690 20404 31696
rect 20456 31726 20576 31754
rect 21284 31754 21312 33322
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 22560 32768 22612 32774
rect 22560 32710 22612 32716
rect 22204 31890 22232 32710
rect 22572 32434 22600 32710
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22744 32292 22796 32298
rect 22744 32234 22796 32240
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21284 31726 21404 31754
rect 20456 30122 20484 31726
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20444 30116 20496 30122
rect 20444 30058 20496 30064
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 20364 28014 20392 29582
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20272 25362 20300 26862
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20364 26042 20392 26318
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20180 23118 20208 24686
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20180 20942 20208 22442
rect 20272 22438 20300 23598
rect 20364 23186 20392 24006
rect 20456 23798 20484 30058
rect 20732 28218 20760 31078
rect 21180 30932 21232 30938
rect 21180 30874 21232 30880
rect 20812 29572 20864 29578
rect 20812 29514 20864 29520
rect 20824 28626 20852 29514
rect 20996 29028 21048 29034
rect 20996 28970 21048 28976
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 21008 27946 21036 28970
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 20996 27940 21048 27946
rect 20996 27882 21048 27888
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20640 25362 20668 26182
rect 20732 26042 20760 26862
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20824 25974 20852 26182
rect 20916 25974 20944 26726
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 21008 25498 21036 27882
rect 20996 25492 21048 25498
rect 20996 25434 21048 25440
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20824 24818 20852 25094
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20548 24206 20576 24550
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 21008 23730 21036 24550
rect 21100 23866 21128 28358
rect 21192 25226 21220 30874
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 21284 27470 21312 29446
rect 21376 29170 21404 31726
rect 21638 29744 21694 29753
rect 21638 29679 21694 29688
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21376 26518 21404 29106
rect 21652 28218 21680 29679
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21652 27606 21680 28154
rect 21836 28082 21864 31758
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 21914 28656 21970 28665
rect 21914 28591 21970 28600
rect 21928 28558 21956 28591
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21560 27130 21588 27270
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21364 26512 21416 26518
rect 21364 26454 21416 26460
rect 21456 26308 21508 26314
rect 21456 26250 21508 26256
rect 21468 25974 21496 26250
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21468 25702 21496 25910
rect 21744 25770 21772 27950
rect 21836 27062 21864 28018
rect 21928 27946 21956 28494
rect 21916 27940 21968 27946
rect 21916 27882 21968 27888
rect 22020 27538 22048 28970
rect 22204 28082 22232 29446
rect 22756 28626 22784 32234
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22848 32026 22876 32166
rect 22836 32020 22888 32026
rect 22836 31962 22888 31968
rect 22940 29306 22968 35022
rect 23952 32434 23980 37130
rect 24504 37126 24532 39200
rect 25792 37262 25820 39200
rect 27724 37262 27752 39200
rect 29012 37262 29040 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 29000 37256 29052 37262
rect 30300 37244 30328 39200
rect 32232 37262 32260 39200
rect 33520 37262 33548 39200
rect 34808 37262 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36740 37262 36768 39200
rect 37186 38176 37242 38185
rect 37186 38111 37242 38120
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 29000 37198 29052 37204
rect 30380 37198 30432 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24596 35290 24624 37198
rect 31484 37188 31536 37194
rect 31484 37130 31536 37136
rect 27804 37120 27856 37126
rect 27804 37062 27856 37068
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30656 37120 30708 37126
rect 30656 37062 30708 37068
rect 27816 36922 27844 37062
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 24688 30734 24716 36858
rect 29000 33312 29052 33318
rect 29000 33254 29052 33260
rect 26148 32292 26200 32298
rect 26148 32234 26200 32240
rect 25134 31920 25190 31929
rect 25134 31855 25190 31864
rect 25148 31822 25176 31855
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24872 30938 24900 31622
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24676 30728 24728 30734
rect 24398 30696 24454 30705
rect 24676 30670 24728 30676
rect 24398 30631 24454 30640
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 23584 29238 23612 29786
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22848 28626 22876 28902
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 21824 27056 21876 27062
rect 21824 26998 21876 27004
rect 22204 26926 22232 27814
rect 22744 27600 22796 27606
rect 22744 27542 22796 27548
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 22652 26240 22704 26246
rect 22652 26182 22704 26188
rect 21928 25838 21956 26182
rect 21916 25832 21968 25838
rect 21916 25774 21968 25780
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 22664 25362 22692 26182
rect 22756 25498 22784 27542
rect 23308 27334 23336 28970
rect 23400 27606 23428 29106
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23492 27470 23520 27950
rect 23584 27470 23612 29174
rect 24032 28756 24084 28762
rect 24032 28698 24084 28704
rect 23664 28416 23716 28422
rect 23664 28358 23716 28364
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20904 23520 20956 23526
rect 20904 23462 20956 23468
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20824 22574 20852 23190
rect 20916 22710 20944 23462
rect 21100 22778 21128 23802
rect 21192 23254 21220 25162
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21192 22778 21220 23054
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20272 22166 20300 22374
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20732 21622 20760 21966
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19984 19236 20036 19242
rect 20180 19224 20208 20742
rect 20272 20398 20300 21286
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20272 19990 20300 20334
rect 20364 20058 20392 20470
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20548 19514 20576 20878
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 19984 19178 20036 19184
rect 20088 19196 20208 19224
rect 20444 19236 20496 19242
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19260 18686 19380 18714
rect 19628 18698 19656 18838
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19260 14482 19288 16662
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14936 2446 14964 4966
rect 16868 2446 16896 4966
rect 18156 2650 18184 8910
rect 18340 5710 18368 12038
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18708 5234 18736 12582
rect 19352 8634 19380 18686
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19444 17882 19472 18158
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19536 16794 19564 17070
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19628 16590 19656 17138
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19904 16454 19932 17002
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15502 19656 15846
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20088 12434 20116 19196
rect 20444 19178 20496 19184
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20180 18358 20208 18634
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20272 17882 20300 18158
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20456 17202 20484 19178
rect 20732 18970 20760 20878
rect 20824 20602 20852 21422
rect 21008 21146 21036 21422
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21284 21010 21312 22986
rect 21376 22030 21404 24618
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21468 23730 21496 24006
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 21284 20058 21312 20946
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21376 19922 21404 21966
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20824 18766 20852 19314
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20916 18630 20944 19790
rect 21192 19514 21220 19790
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20364 14890 20392 16526
rect 20548 16250 20576 17614
rect 20824 17202 20852 17750
rect 21008 17270 21036 18294
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21100 17338 21128 17614
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20456 13938 20484 16050
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20088 12406 20576 12434
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20548 11150 20576 12406
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 19444 2446 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20272 5234 20300 10406
rect 21192 5710 21220 11018
rect 21376 9178 21404 19858
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21468 7002 21496 21898
rect 21560 20058 21588 25230
rect 22284 24608 22336 24614
rect 22284 24550 22336 24556
rect 22296 23050 22324 24550
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21652 21690 21680 22918
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21652 21010 21680 21626
rect 22112 21554 22140 22510
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 19378 22140 19654
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22204 18766 22232 19178
rect 22296 18902 22324 19790
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22112 17746 22140 18158
rect 22204 17882 22232 18294
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22388 17814 22416 23598
rect 22756 22982 22784 24006
rect 22848 23798 22876 26998
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23308 26586 23336 26862
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 23492 26382 23520 27270
rect 23584 26450 23612 27270
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23112 25968 23164 25974
rect 23112 25910 23164 25916
rect 23124 25770 23152 25910
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 23676 25498 23704 28358
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23768 25906 23796 26386
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23676 24750 23704 25434
rect 23768 25430 23796 25842
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23756 25424 23808 25430
rect 23756 25366 23808 25372
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23756 24676 23808 24682
rect 23756 24618 23808 24624
rect 22836 23792 22888 23798
rect 22836 23734 22888 23740
rect 22848 23186 22876 23734
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22664 21690 22692 21898
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22848 21162 22876 21354
rect 22848 21146 23060 21162
rect 22848 21140 23072 21146
rect 22848 21134 23020 21140
rect 23020 21082 23072 21088
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 20330 22600 20878
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21928 12102 21956 17682
rect 22388 17066 22416 17750
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 22020 10742 22048 16934
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 22388 8634 22416 11766
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 22020 2650 22048 8434
rect 22480 7206 22508 19858
rect 22572 16114 22600 20266
rect 22756 19990 22784 20334
rect 22848 20058 22876 20470
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22756 19514 22784 19926
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22940 18970 22968 19246
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22848 17338 22876 17614
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22664 2446 22692 4966
rect 23124 4146 23152 18158
rect 23216 5710 23244 19790
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23308 19378 23336 19722
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23308 18766 23336 19314
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23400 18086 23428 22510
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 21962 23520 22374
rect 23768 21962 23796 24618
rect 23860 24274 23888 25638
rect 23952 24410 23980 27338
rect 24044 26790 24072 28698
rect 24216 27464 24268 27470
rect 24216 27406 24268 27412
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23952 23730 23980 24346
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 22710 23888 23122
rect 24044 22778 24072 26726
rect 24124 26240 24176 26246
rect 24124 26182 24176 26188
rect 24136 25362 24164 26182
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24032 22772 24084 22778
rect 24032 22714 24084 22720
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 18970 23520 19790
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23676 18766 23704 19450
rect 23768 18766 23796 21898
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 10674 23612 16594
rect 23860 12850 23888 22646
rect 24228 21622 24256 27406
rect 24320 24342 24348 27406
rect 24412 24818 24440 30631
rect 24872 30258 24900 30874
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 25056 30122 25084 31282
rect 25044 30116 25096 30122
rect 25044 30058 25096 30064
rect 25148 29646 25176 31758
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25240 31346 25268 31622
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25320 31204 25372 31210
rect 25320 31146 25372 31152
rect 25332 30666 25360 31146
rect 25320 30660 25372 30666
rect 25320 30602 25372 30608
rect 25136 29640 25188 29646
rect 25136 29582 25188 29588
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24584 28688 24636 28694
rect 24584 28630 24636 28636
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24308 24336 24360 24342
rect 24308 24278 24360 24284
rect 24412 23866 24440 24550
rect 24504 24274 24532 26862
rect 24596 25906 24624 28630
rect 24964 28082 24992 29446
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24780 26994 24808 27814
rect 25332 27130 25360 30602
rect 25516 30326 25544 31758
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 30326 25636 31078
rect 26160 30802 26188 32234
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 26160 30326 26188 30738
rect 25504 30320 25556 30326
rect 25504 30262 25556 30268
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 26148 30320 26200 30326
rect 26148 30262 26200 30268
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 26344 26518 26372 32166
rect 29012 31278 29040 33254
rect 29748 32910 29776 37062
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29000 31272 29052 31278
rect 29000 31214 29052 31220
rect 26608 30932 26660 30938
rect 26608 30874 26660 30880
rect 26620 30734 26648 30874
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 30392 29170 30420 37062
rect 30668 30734 30696 37062
rect 31496 33522 31524 37130
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 32416 35894 32444 37062
rect 32232 35866 32444 35894
rect 34532 35894 34560 37062
rect 35900 36644 35952 36650
rect 35900 36586 35952 36592
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34532 35866 34652 35894
rect 31484 33516 31536 33522
rect 31484 33458 31536 33464
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31772 31482 31800 32710
rect 32232 32434 32260 35866
rect 34244 35080 34296 35086
rect 34244 35022 34296 35028
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32404 32224 32456 32230
rect 32404 32166 32456 32172
rect 32416 31890 32444 32166
rect 32404 31884 32456 31890
rect 32404 31826 32456 31832
rect 31760 31476 31812 31482
rect 31760 31418 31812 31424
rect 32404 31136 32456 31142
rect 32404 31078 32456 31084
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 32416 29238 32444 31078
rect 34256 30122 34284 35022
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34532 32502 34560 33934
rect 34520 32496 34572 32502
rect 34520 32438 34572 32444
rect 34624 30326 34652 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35912 32910 35940 36586
rect 35992 36576 36044 36582
rect 35992 36518 36044 36524
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 36004 32366 36032 36518
rect 37200 36174 37228 38111
rect 37280 37256 37332 37262
rect 37280 37198 37332 37204
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 35992 32360 36044 32366
rect 35992 32302 36044 32308
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36096 31346 36124 35974
rect 37292 34202 37320 37198
rect 38028 36786 38056 39200
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 38212 36825 38240 37062
rect 39316 36854 39344 39200
rect 39304 36848 39356 36854
rect 38198 36816 38254 36825
rect 38016 36780 38068 36786
rect 39304 36790 39356 36796
rect 38198 36751 38254 36760
rect 38016 36722 38068 36728
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 37280 34196 37332 34202
rect 37280 34138 37332 34144
rect 37924 33516 37976 33522
rect 37924 33458 37976 33464
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34612 30320 34664 30326
rect 34612 30262 34664 30268
rect 34428 30252 34480 30258
rect 34428 30194 34480 30200
rect 34244 30116 34296 30122
rect 34244 30058 34296 30064
rect 32404 29232 32456 29238
rect 32404 29174 32456 29180
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31772 26858 31800 27270
rect 34440 27130 34468 30194
rect 37004 30048 37056 30054
rect 37004 29990 37056 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35452 27470 35480 28970
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 34428 27124 34480 27130
rect 34428 27066 34480 27072
rect 37016 26994 37044 29990
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 31760 26852 31812 26858
rect 31760 26794 31812 26800
rect 32588 26784 32640 26790
rect 32588 26726 32640 26732
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24584 25288 24636 25294
rect 24582 25256 24584 25265
rect 24636 25256 24638 25265
rect 24582 25191 24638 25200
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24688 24886 24716 25094
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24492 24268 24544 24274
rect 24492 24210 24544 24216
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24504 22094 24532 24210
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24596 23322 24624 23666
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24780 23118 24808 25366
rect 24964 24410 24992 26250
rect 26608 25968 26660 25974
rect 26608 25910 26660 25916
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 24964 23254 24992 24346
rect 25608 24274 25636 24550
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25884 24206 25912 25230
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26344 24410 26372 24754
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 26620 24206 26648 25910
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 27540 24138 27568 24754
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 24952 23248 25004 23254
rect 24952 23190 25004 23196
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22642 24808 23054
rect 25700 22710 25728 24006
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 30208 22574 30236 24006
rect 32600 23526 32628 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 34532 24818 34560 26318
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 37936 24313 37964 33458
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 32065 38332 32370
rect 38290 32056 38346 32065
rect 38290 31991 38346 32000
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 38304 30025 38332 30194
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 26586 38056 27406
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38016 26580 38068 26586
rect 38016 26522 38068 26528
rect 38016 25696 38068 25702
rect 38016 25638 38068 25644
rect 38028 25294 38056 25638
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 38198 25256 38254 25265
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 37922 24304 37978 24313
rect 37922 24239 37978 24248
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38108 24064 38160 24070
rect 38108 24006 38160 24012
rect 32588 23520 32640 23526
rect 32588 23462 32640 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 38120 22710 38148 24006
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 38108 22704 38160 22710
rect 38108 22646 38160 22652
rect 30196 22568 30248 22574
rect 30196 22510 30248 22516
rect 28264 22432 28316 22438
rect 28264 22374 28316 22380
rect 38016 22432 38068 22438
rect 38016 22374 38068 22380
rect 24412 22066 24532 22094
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20534 24072 20742
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23952 19514 23980 20334
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 24136 8090 24164 18022
rect 24412 11558 24440 22066
rect 24582 21312 24638 21321
rect 24582 21247 24638 21256
rect 24596 20466 24624 21247
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25056 20602 25084 20878
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24504 19378 24532 20266
rect 24596 19854 24624 20402
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26252 16658 26280 18362
rect 26344 17678 26372 20198
rect 28276 19718 28304 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 38028 20942 38056 22374
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38016 20936 38068 20942
rect 38016 20878 38068 20884
rect 38200 20800 38252 20806
rect 38200 20742 38252 20748
rect 38212 20505 38240 20742
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30300 18766 30328 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 34796 18692 34848 18698
rect 34796 18634 34848 18640
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 33060 15502 33088 18566
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 33508 16448 33560 16454
rect 33508 16390 33560 16396
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33520 16114 33548 16390
rect 33704 16250 33732 16390
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33508 16108 33560 16114
rect 33508 16050 33560 16056
rect 33324 15904 33376 15910
rect 33324 15846 33376 15852
rect 33048 15496 33100 15502
rect 33048 15438 33100 15444
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24688 5710 24716 12582
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23216 2446 23244 5510
rect 24872 2650 24900 8434
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25424 2514 25452 6734
rect 25608 5234 25636 10406
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25412 2508 25464 2514
rect 25412 2450 25464 2456
rect 25884 2446 25912 5510
rect 28368 4622 28396 10406
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28644 2650 28672 7822
rect 28920 6458 28948 14418
rect 33336 12850 33364 15846
rect 34532 14414 34560 17478
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 34808 7886 34836 18634
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 38028 17202 38056 18566
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35808 16652 35860 16658
rect 35808 16594 35860 16600
rect 35820 16250 35848 16594
rect 35808 16244 35860 16250
rect 35808 16186 35860 16192
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14414 35388 15846
rect 38304 15745 38332 16050
rect 38290 15736 38346 15745
rect 38290 15671 38346 15680
rect 38016 15360 38068 15366
rect 38016 15302 38068 15308
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 37280 14272 37332 14278
rect 37280 14214 37332 14220
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35348 12640 35400 12646
rect 35348 12582 35400 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 8974 35388 12582
rect 37292 11150 37320 14214
rect 38028 12850 38056 15302
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 37096 7744 37148 7750
rect 37096 7686 37148 7692
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 30300 2582 30328 6258
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 32588 5704 32640 5710
rect 32588 5646 32640 5652
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 31680 2446 31708 4966
rect 32600 2650 32628 5646
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 32588 2644 32640 2650
rect 32588 2586 32640 2592
rect 33980 2514 34008 4422
rect 34532 3738 34560 5646
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 35820 3194 35848 7346
rect 37108 5710 37136 7686
rect 37278 6216 37334 6225
rect 37278 6151 37334 6160
rect 37292 6118 37320 6151
rect 37280 6112 37332 6118
rect 37280 6054 37332 6060
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 37832 5568 37884 5574
rect 37832 5510 37884 5516
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37476 3534 37504 3878
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 37844 3058 37872 5510
rect 37936 4826 37964 11698
rect 38120 8090 38148 12174
rect 38200 11280 38252 11286
rect 38200 11222 38252 11228
rect 38212 10985 38240 11222
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38108 8084 38160 8090
rect 38108 8026 38160 8032
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38108 6316 38160 6322
rect 38108 6258 38160 6264
rect 38120 6225 38148 6258
rect 38106 6216 38162 6225
rect 38106 6151 38162 6160
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4185 38332 4558
rect 38290 4176 38346 4185
rect 38290 4111 38346 4120
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33968 2508 34020 2514
rect 33968 2450 34020 2456
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 800 11652 2246
rect 13556 800 13584 2382
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 14844 800 14872 2246
rect 16776 800 16804 2246
rect 18064 800 18092 2382
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 22572 800 22600 2246
rect 23860 800 23888 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2382
rect 29012 800 29040 2382
rect 30300 800 30328 2382
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 800 31616 2246
rect 33520 800 33548 2382
rect 34808 800 34836 2382
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 36096 800 36124 2246
rect 36924 1465 36952 2994
rect 38028 2446 38056 3334
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38120 1986 38148 3470
rect 38200 2848 38252 2854
rect 38198 2816 38200 2825
rect 38252 2816 38254 2825
rect 38198 2751 38254 2760
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 38028 1958 38148 1986
rect 36910 1456 36966 1465
rect 36910 1391 36966 1400
rect 38028 800 38056 1958
rect 39316 800 39344 2246
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 1306 35808 1362 35864
rect 1766 33360 1822 33416
rect 1858 31728 1914 31784
rect 1674 30640 1730 30696
rect 1858 29588 1860 29608
rect 1860 29588 1912 29608
rect 1912 29588 1914 29608
rect 1858 29552 1914 29588
rect 1858 28092 1860 28112
rect 1860 28092 1912 28112
rect 1912 28092 1914 28112
rect 1858 28056 1914 28092
rect 1858 27668 1914 27704
rect 1858 27648 1860 27668
rect 1860 27648 1912 27668
rect 1912 27648 1914 27668
rect 1766 27240 1822 27296
rect 1766 25200 1822 25256
rect 1766 23840 1822 23896
rect 1766 22480 1822 22536
rect 1766 20440 1822 20496
rect 1766 19080 1822 19136
rect 2318 33532 2320 33552
rect 2320 33532 2372 33552
rect 2372 33532 2374 33552
rect 2318 33496 2374 33532
rect 2318 28908 2320 28928
rect 2320 28908 2372 28928
rect 2372 28908 2374 28928
rect 2318 28872 2374 28908
rect 2870 32272 2926 32328
rect 3330 35572 3332 35592
rect 3332 35572 3384 35592
rect 3384 35572 3386 35592
rect 3330 35536 3386 35572
rect 3238 34992 3294 35048
rect 4066 38120 4122 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4434 36796 4436 36816
rect 4436 36796 4488 36816
rect 4488 36796 4490 36816
rect 4434 36760 4490 36796
rect 3606 36216 3662 36272
rect 3882 36216 3938 36272
rect 4618 36488 4674 36544
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 5722 37068 5724 37088
rect 5724 37068 5776 37088
rect 5776 37068 5778 37088
rect 5722 37032 5778 37068
rect 4802 35944 4858 36000
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3330 34892 3332 34912
rect 3332 34892 3384 34912
rect 3384 34892 3386 34912
rect 3330 34856 3386 34892
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4526 33396 4528 33416
rect 4528 33396 4580 33416
rect 4580 33396 4582 33416
rect 2686 28056 2742 28112
rect 2410 27920 2466 27976
rect 3146 28600 3202 28656
rect 3422 26968 3478 27024
rect 3606 27512 3662 27568
rect 3606 26832 3662 26888
rect 4526 33360 4582 33396
rect 4618 33224 4674 33280
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4066 32272 4122 32328
rect 3974 31864 4030 31920
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4526 31864 4582 31920
rect 3790 29008 3846 29064
rect 3790 28192 3846 28248
rect 3606 23840 3662 23896
rect 2318 23044 2374 23080
rect 2318 23024 2320 23044
rect 2320 23024 2372 23044
rect 2372 23024 2374 23044
rect 4986 33360 5042 33416
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4526 30368 4582 30424
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4526 29572 4582 29608
rect 4526 29552 4528 29572
rect 4528 29552 4580 29572
rect 4580 29552 4582 29572
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4434 28600 4490 28656
rect 3974 28192 4030 28248
rect 4342 28328 4398 28384
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3974 25336 4030 25392
rect 4618 26968 4674 27024
rect 4802 32000 4858 32056
rect 4986 31184 5042 31240
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4066 24656 4122 24712
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5538 34448 5594 34504
rect 5262 32680 5318 32736
rect 5170 30640 5226 30696
rect 5078 30096 5134 30152
rect 5446 30232 5502 30288
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 5078 25064 5134 25120
rect 7378 36352 7434 36408
rect 7286 35944 7342 36000
rect 7010 35672 7066 35728
rect 5538 24812 5594 24848
rect 5538 24792 5540 24812
rect 5540 24792 5592 24812
rect 5592 24792 5594 24812
rect 5722 25472 5778 25528
rect 6182 26424 6238 26480
rect 6734 34196 6790 34232
rect 6734 34176 6736 34196
rect 6736 34176 6788 34196
rect 6788 34176 6790 34196
rect 6550 33224 6606 33280
rect 6826 32272 6882 32328
rect 8482 37068 8484 37088
rect 8484 37068 8536 37088
rect 8536 37068 8538 37088
rect 8482 37032 8538 37068
rect 8850 37032 8906 37088
rect 8666 36896 8722 36952
rect 6550 26560 6606 26616
rect 7470 29688 7526 29744
rect 8758 36660 8760 36680
rect 8760 36660 8812 36680
rect 8812 36660 8814 36680
rect 7746 29144 7802 29200
rect 7654 27648 7710 27704
rect 7286 25608 7342 25664
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1766 17720 1822 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1766 15680 1822 15736
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1766 12280 1822 12336
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1766 10920 1822 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 7562 24656 7618 24712
rect 7746 24556 7748 24576
rect 7748 24556 7800 24576
rect 7800 24556 7802 24576
rect 7746 24520 7802 24556
rect 8390 35264 8446 35320
rect 8298 34040 8354 34096
rect 8206 33940 8208 33960
rect 8208 33940 8260 33960
rect 8260 33940 8262 33960
rect 8206 33904 8262 33940
rect 8758 36624 8814 36660
rect 8942 36216 8998 36272
rect 8942 35944 8998 36000
rect 8574 35672 8630 35728
rect 9586 36896 9642 36952
rect 9402 36624 9458 36680
rect 9218 36216 9274 36272
rect 9586 35672 9642 35728
rect 9494 34856 9550 34912
rect 8390 33088 8446 33144
rect 8114 32020 8170 32056
rect 8114 32000 8116 32020
rect 8116 32000 8168 32020
rect 8168 32000 8170 32020
rect 8666 32272 8722 32328
rect 7930 26288 7986 26344
rect 7654 22208 7710 22264
rect 9218 32272 9274 32328
rect 8206 29960 8262 30016
rect 8298 24928 8354 24984
rect 8758 29008 8814 29064
rect 9126 31320 9182 31376
rect 9126 29552 9182 29608
rect 8942 27920 8998 27976
rect 8850 26832 8906 26888
rect 8942 26152 8998 26208
rect 9126 25880 9182 25936
rect 8758 24384 8814 24440
rect 10046 36080 10102 36136
rect 9954 35400 10010 35456
rect 9770 33632 9826 33688
rect 9586 32988 9588 33008
rect 9588 32988 9640 33008
rect 9640 32988 9642 33008
rect 9586 32952 9642 32988
rect 9402 32852 9404 32872
rect 9404 32852 9456 32872
rect 9456 32852 9458 32872
rect 9402 32816 9458 32852
rect 9402 32716 9404 32736
rect 9404 32716 9456 32736
rect 9456 32716 9458 32736
rect 9402 32680 9458 32716
rect 9402 29280 9458 29336
rect 9678 31728 9734 31784
rect 9954 33224 10010 33280
rect 9862 32000 9918 32056
rect 9770 29552 9826 29608
rect 9954 29280 10010 29336
rect 10506 35128 10562 35184
rect 12346 37168 12402 37224
rect 12254 37032 12310 37088
rect 11610 36760 11666 36816
rect 10966 36488 11022 36544
rect 10598 34992 10654 35048
rect 10138 30096 10194 30152
rect 9586 26560 9642 26616
rect 9862 28736 9918 28792
rect 10046 28464 10102 28520
rect 9310 25200 9366 25256
rect 9218 21936 9274 21992
rect 9126 19372 9182 19408
rect 9126 19352 9128 19372
rect 9128 19352 9180 19372
rect 9180 19352 9182 19372
rect 8390 17992 8446 18048
rect 1766 9560 1822 9616
rect 1766 7520 1822 7576
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1858 5344 1914 5400
rect 1674 4800 1730 4856
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1766 2760 1822 2816
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9862 24520 9918 24576
rect 9586 24384 9642 24440
rect 10414 33224 10470 33280
rect 10598 33632 10654 33688
rect 11150 36080 11206 36136
rect 10874 35436 10876 35456
rect 10876 35436 10928 35456
rect 10928 35436 10930 35456
rect 10874 35400 10930 35436
rect 10782 32544 10838 32600
rect 10506 31456 10562 31512
rect 10598 31320 10654 31376
rect 10414 30776 10470 30832
rect 11150 35264 11206 35320
rect 11150 34856 11206 34912
rect 11150 34720 11206 34776
rect 11242 34312 11298 34368
rect 10690 30776 10746 30832
rect 10598 29280 10654 29336
rect 10874 30368 10930 30424
rect 10782 28872 10838 28928
rect 10966 28736 11022 28792
rect 10322 28328 10378 28384
rect 10598 28328 10654 28384
rect 10322 26016 10378 26072
rect 9862 21936 9918 21992
rect 9586 20848 9642 20904
rect 9402 20748 9404 20768
rect 9404 20748 9456 20768
rect 9456 20748 9458 20768
rect 9402 20712 9458 20748
rect 10690 28192 10746 28248
rect 11426 34176 11482 34232
rect 12346 36916 12402 36952
rect 12346 36896 12348 36916
rect 12348 36896 12400 36916
rect 12400 36896 12402 36916
rect 12346 36216 12402 36272
rect 12530 36760 12586 36816
rect 12622 36352 12678 36408
rect 13174 36080 13230 36136
rect 11794 35944 11850 36000
rect 12254 35944 12310 36000
rect 11702 34448 11758 34504
rect 11610 34176 11666 34232
rect 11610 33632 11666 33688
rect 11518 33496 11574 33552
rect 12254 35672 12310 35728
rect 12622 35672 12678 35728
rect 12438 35536 12494 35592
rect 13082 35944 13138 36000
rect 12530 34584 12586 34640
rect 12438 34176 12494 34232
rect 11886 33768 11942 33824
rect 11794 32680 11850 32736
rect 11702 32272 11758 32328
rect 11150 26832 11206 26888
rect 11426 28736 11482 28792
rect 11426 28192 11482 28248
rect 10966 25744 11022 25800
rect 10138 19216 10194 19272
rect 9678 19080 9734 19136
rect 10046 18808 10102 18864
rect 10506 22480 10562 22536
rect 10322 22108 10324 22128
rect 10324 22108 10376 22128
rect 10376 22108 10378 22128
rect 10322 22072 10378 22108
rect 10506 21956 10562 21992
rect 10506 21936 10508 21956
rect 10508 21936 10560 21956
rect 10560 21936 10562 21956
rect 10966 24248 11022 24304
rect 11058 22092 11114 22128
rect 11058 22072 11060 22092
rect 11060 22072 11112 22092
rect 11112 22072 11114 22092
rect 11702 28464 11758 28520
rect 12070 31748 12126 31784
rect 12070 31728 12072 31748
rect 12072 31728 12124 31748
rect 12124 31728 12126 31748
rect 12346 32408 12402 32464
rect 12622 33496 12678 33552
rect 12530 31456 12586 31512
rect 12070 29960 12126 30016
rect 11978 29008 12034 29064
rect 13266 34892 13268 34912
rect 13268 34892 13320 34912
rect 13320 34892 13322 34912
rect 13266 34856 13322 34892
rect 13174 34312 13230 34368
rect 12254 29008 12310 29064
rect 12162 26560 12218 26616
rect 11242 20712 11298 20768
rect 11058 20440 11114 20496
rect 10966 19372 11022 19408
rect 10966 19352 10968 19372
rect 10968 19352 11020 19372
rect 11020 19352 11022 19372
rect 12162 26288 12218 26344
rect 12438 26560 12494 26616
rect 12346 24248 12402 24304
rect 12162 23316 12218 23352
rect 12162 23296 12164 23316
rect 12164 23296 12216 23316
rect 12216 23296 12218 23316
rect 11610 21972 11612 21992
rect 11612 21972 11664 21992
rect 11664 21972 11666 21992
rect 11610 21936 11666 21972
rect 11702 21392 11758 21448
rect 11334 19216 11390 19272
rect 12254 22516 12256 22536
rect 12256 22516 12308 22536
rect 12308 22516 12310 22536
rect 12254 22480 12310 22516
rect 12254 21936 12310 21992
rect 12898 29144 12954 29200
rect 13174 29028 13230 29064
rect 13174 29008 13176 29028
rect 13176 29008 13228 29028
rect 13228 29008 13230 29028
rect 13082 25608 13138 25664
rect 13634 36524 13636 36544
rect 13636 36524 13688 36544
rect 13688 36524 13690 36544
rect 13634 36488 13690 36524
rect 13542 33224 13598 33280
rect 13726 34720 13782 34776
rect 14370 37168 14426 37224
rect 14002 34740 14058 34776
rect 14278 34992 14334 35048
rect 14002 34720 14004 34740
rect 14004 34720 14056 34740
rect 14056 34720 14058 34740
rect 13726 32680 13782 32736
rect 13450 31340 13506 31376
rect 13450 31320 13452 31340
rect 13452 31320 13504 31340
rect 13504 31320 13506 31340
rect 13450 30368 13506 30424
rect 13450 27920 13506 27976
rect 13358 25880 13414 25936
rect 14002 32952 14058 33008
rect 14830 36896 14886 36952
rect 14370 32308 14372 32328
rect 14372 32308 14424 32328
rect 14424 32308 14426 32328
rect 14370 32272 14426 32308
rect 15566 35944 15622 36000
rect 14370 31884 14426 31920
rect 14370 31864 14372 31884
rect 14372 31864 14424 31884
rect 14424 31864 14426 31884
rect 13910 26560 13966 26616
rect 13818 25472 13874 25528
rect 13450 24112 13506 24168
rect 12622 18808 12678 18864
rect 12346 15952 12402 16008
rect 13542 22208 13598 22264
rect 13358 20848 13414 20904
rect 15014 34740 15070 34776
rect 15014 34720 15016 34740
rect 15016 34720 15068 34740
rect 15068 34720 15070 34740
rect 15198 33768 15254 33824
rect 15658 33904 15714 33960
rect 15934 33632 15990 33688
rect 15658 32544 15714 32600
rect 13726 18944 13782 19000
rect 14370 23160 14426 23216
rect 15014 30232 15070 30288
rect 14738 26288 14794 26344
rect 15566 30776 15622 30832
rect 15474 26868 15476 26888
rect 15476 26868 15528 26888
rect 15528 26868 15530 26888
rect 15474 26832 15530 26868
rect 15014 26424 15070 26480
rect 14554 21392 14610 21448
rect 1766 1400 1822 1456
rect 14370 19080 14426 19136
rect 14370 16904 14426 16960
rect 13726 14456 13782 14512
rect 15566 26016 15622 26072
rect 17130 36100 17186 36136
rect 17130 36080 17132 36100
rect 17132 36080 17184 36100
rect 17184 36080 17186 36100
rect 17590 35128 17646 35184
rect 19246 35808 19302 35864
rect 16946 30096 17002 30152
rect 16854 28056 16910 28112
rect 16762 26560 16818 26616
rect 15474 22636 15530 22672
rect 15474 22616 15476 22636
rect 15476 22616 15528 22636
rect 15528 22616 15530 22636
rect 15474 20460 15530 20496
rect 15474 20440 15476 20460
rect 15476 20440 15528 20460
rect 15528 20440 15530 20460
rect 15198 13640 15254 13696
rect 17774 29688 17830 29744
rect 17590 26852 17646 26888
rect 17590 26832 17592 26852
rect 17592 26832 17644 26852
rect 17644 26832 17646 26852
rect 17590 26016 17646 26072
rect 16486 22752 16542 22808
rect 17958 26968 18014 27024
rect 19338 33088 19394 33144
rect 17038 13932 17094 13968
rect 17038 13912 17040 13932
rect 17040 13912 17092 13932
rect 17092 13912 17094 13932
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20166 36624 20222 36680
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19522 29708 19578 29744
rect 19522 29688 19524 29708
rect 19524 29688 19576 29708
rect 19576 29688 19578 29708
rect 19614 29552 19670 29608
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19522 29144 19578 29200
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18694 17720 18750 17776
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19706 24248 19762 24304
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 21638 29688 21694 29744
rect 21914 28600 21970 28656
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38120 37242 38176
rect 25134 31864 25190 31920
rect 24398 30640 24454 30696
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 38198 36760 38254 36816
rect 38198 34720 38254 34776
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 24582 25236 24584 25256
rect 24584 25236 24636 25256
rect 24636 25236 24638 25256
rect 24582 25200 24638 25236
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 32000 38346 32056
rect 38290 29960 38346 30016
rect 38290 28600 38346 28656
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38198 25200 38254 25256
rect 37922 24248 37978 24304
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 38290 23840 38346 23896
rect 24582 21256 24638 21312
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 38290 21800 38346 21856
rect 38198 20440 38254 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38290 15680 38346 15736
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38198 14320 38254 14376
rect 38198 12280 38254 12336
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 37278 6160 37334 6216
rect 38198 10920 38254 10976
rect 38198 8880 38254 8936
rect 38290 7520 38346 7576
rect 38106 6160 38162 6216
rect 38290 4120 38346 4176
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38198 2796 38200 2816
rect 38200 2796 38252 2816
rect 38252 2796 38254 2816
rect 38198 2760 38254 2796
rect 36910 1400 36966 1456
<< metal3 >>
rect 200 38178 800 38208
rect 4061 38178 4127 38181
rect 200 38176 4127 38178
rect 200 38120 4066 38176
rect 4122 38120 4127 38176
rect 200 38118 4127 38120
rect 200 38088 800 38118
rect 4061 38115 4127 38118
rect 37181 38178 37247 38181
rect 39200 38178 39800 38208
rect 37181 38176 39800 38178
rect 37181 38120 37186 38176
rect 37242 38120 39800 38176
rect 37181 38118 39800 38120
rect 37181 38115 37247 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 12341 37226 12407 37229
rect 14365 37226 14431 37229
rect 12341 37224 14431 37226
rect 12341 37168 12346 37224
rect 12402 37168 14370 37224
rect 14426 37168 14431 37224
rect 12341 37166 14431 37168
rect 12341 37163 12407 37166
rect 14365 37163 14431 37166
rect 5717 37092 5783 37093
rect 8477 37092 8543 37093
rect 5717 37090 5764 37092
rect 5672 37088 5764 37090
rect 5672 37032 5722 37088
rect 5672 37030 5764 37032
rect 5717 37028 5764 37030
rect 5828 37028 5834 37092
rect 8477 37090 8524 37092
rect 8432 37088 8524 37090
rect 8432 37032 8482 37088
rect 8432 37030 8524 37032
rect 8477 37028 8524 37030
rect 8588 37028 8594 37092
rect 8845 37090 8911 37093
rect 12249 37090 12315 37093
rect 8845 37088 12315 37090
rect 8845 37032 8850 37088
rect 8906 37032 12254 37088
rect 12310 37032 12315 37088
rect 8845 37030 12315 37032
rect 5717 37027 5783 37028
rect 8477 37027 8543 37028
rect 8845 37027 8911 37030
rect 12249 37027 12315 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 8661 36954 8727 36957
rect 4294 36952 8727 36954
rect 4294 36896 8666 36952
rect 8722 36896 8727 36952
rect 4294 36894 8727 36896
rect 200 36818 800 36848
rect 4294 36818 4354 36894
rect 8661 36891 8727 36894
rect 9581 36954 9647 36957
rect 12341 36954 12407 36957
rect 14825 36954 14891 36957
rect 9581 36952 12082 36954
rect 9581 36896 9586 36952
rect 9642 36896 12082 36952
rect 9581 36894 12082 36896
rect 9581 36891 9647 36894
rect 200 36758 4354 36818
rect 4429 36818 4495 36821
rect 11605 36818 11671 36821
rect 4429 36816 11671 36818
rect 4429 36760 4434 36816
rect 4490 36760 11610 36816
rect 11666 36760 11671 36816
rect 4429 36758 11671 36760
rect 12022 36818 12082 36894
rect 12341 36952 14891 36954
rect 12341 36896 12346 36952
rect 12402 36896 14830 36952
rect 14886 36896 14891 36952
rect 12341 36894 14891 36896
rect 12341 36891 12407 36894
rect 14825 36891 14891 36894
rect 12525 36818 12591 36821
rect 12022 36816 12591 36818
rect 12022 36760 12530 36816
rect 12586 36760 12591 36816
rect 12022 36758 12591 36760
rect 200 36728 800 36758
rect 4429 36755 4495 36758
rect 11605 36755 11671 36758
rect 12525 36755 12591 36758
rect 38193 36818 38259 36821
rect 39200 36818 39800 36848
rect 38193 36816 39800 36818
rect 38193 36760 38198 36816
rect 38254 36760 39800 36816
rect 38193 36758 39800 36760
rect 38193 36755 38259 36758
rect 39200 36728 39800 36758
rect 8753 36682 8819 36685
rect 9397 36682 9463 36685
rect 20161 36682 20227 36685
rect 8753 36680 20227 36682
rect 8753 36624 8758 36680
rect 8814 36624 9402 36680
rect 9458 36624 20166 36680
rect 20222 36624 20227 36680
rect 8753 36622 20227 36624
rect 8753 36619 8819 36622
rect 9397 36619 9463 36622
rect 20161 36619 20227 36622
rect 4613 36546 4679 36549
rect 8518 36546 8524 36548
rect 4613 36544 8524 36546
rect 4613 36488 4618 36544
rect 4674 36488 8524 36544
rect 4613 36486 8524 36488
rect 4613 36483 4679 36486
rect 8518 36484 8524 36486
rect 8588 36484 8594 36548
rect 10961 36546 11027 36549
rect 13486 36546 13492 36548
rect 10961 36544 13492 36546
rect 10961 36488 10966 36544
rect 11022 36488 13492 36544
rect 10961 36486 13492 36488
rect 10961 36483 11027 36486
rect 13486 36484 13492 36486
rect 13556 36546 13562 36548
rect 13629 36546 13695 36549
rect 13556 36544 13695 36546
rect 13556 36488 13634 36544
rect 13690 36488 13695 36544
rect 13556 36486 13695 36488
rect 13556 36484 13562 36486
rect 13629 36483 13695 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 7373 36410 7439 36413
rect 12617 36410 12683 36413
rect 7373 36408 12683 36410
rect 7373 36352 7378 36408
rect 7434 36352 12622 36408
rect 12678 36352 12683 36408
rect 7373 36350 12683 36352
rect 7373 36347 7439 36350
rect 12617 36347 12683 36350
rect 2078 36212 2084 36276
rect 2148 36274 2154 36276
rect 3601 36274 3667 36277
rect 2148 36272 3667 36274
rect 2148 36216 3606 36272
rect 3662 36216 3667 36272
rect 2148 36214 3667 36216
rect 2148 36212 2154 36214
rect 3601 36211 3667 36214
rect 3877 36274 3943 36277
rect 8937 36274 9003 36277
rect 3877 36272 9003 36274
rect 3877 36216 3882 36272
rect 3938 36216 8942 36272
rect 8998 36216 9003 36272
rect 3877 36214 9003 36216
rect 3877 36211 3943 36214
rect 8937 36211 9003 36214
rect 9213 36274 9279 36277
rect 12341 36274 12407 36277
rect 9213 36272 12407 36274
rect 9213 36216 9218 36272
rect 9274 36216 12346 36272
rect 12402 36216 12407 36272
rect 9213 36214 12407 36216
rect 9213 36211 9279 36214
rect 12341 36211 12407 36214
rect 5206 36076 5212 36140
rect 5276 36138 5282 36140
rect 10041 36138 10107 36141
rect 11145 36140 11211 36141
rect 11094 36138 11100 36140
rect 5276 36136 10107 36138
rect 5276 36080 10046 36136
rect 10102 36080 10107 36136
rect 5276 36078 10107 36080
rect 11054 36078 11100 36138
rect 11164 36136 11211 36140
rect 11206 36080 11211 36136
rect 5276 36076 5282 36078
rect 10041 36075 10107 36078
rect 11094 36076 11100 36078
rect 11164 36076 11211 36080
rect 11145 36075 11211 36076
rect 13169 36138 13235 36141
rect 17125 36138 17191 36141
rect 13169 36136 17191 36138
rect 13169 36080 13174 36136
rect 13230 36080 17130 36136
rect 17186 36080 17191 36136
rect 13169 36078 17191 36080
rect 13169 36075 13235 36078
rect 17125 36075 17191 36078
rect 4797 36004 4863 36005
rect 7281 36004 7347 36005
rect 4797 36000 4844 36004
rect 4908 36002 4914 36004
rect 7230 36002 7236 36004
rect 4797 35944 4802 36000
rect 4797 35940 4844 35944
rect 4908 35942 4954 36002
rect 7190 35942 7236 36002
rect 7300 36000 7347 36004
rect 7342 35944 7347 36000
rect 4908 35940 4914 35942
rect 7230 35940 7236 35942
rect 7300 35940 7347 35944
rect 4797 35939 4863 35940
rect 7281 35939 7347 35940
rect 8937 36002 9003 36005
rect 11789 36002 11855 36005
rect 8937 36000 11855 36002
rect 8937 35944 8942 36000
rect 8998 35944 11794 36000
rect 11850 35944 11855 36000
rect 8937 35942 11855 35944
rect 8937 35939 9003 35942
rect 11789 35939 11855 35942
rect 12249 36002 12315 36005
rect 13077 36002 13143 36005
rect 12249 36000 13143 36002
rect 12249 35944 12254 36000
rect 12310 35944 13082 36000
rect 13138 35944 13143 36000
rect 12249 35942 13143 35944
rect 12249 35939 12315 35942
rect 13077 35939 13143 35942
rect 15561 36002 15627 36005
rect 15694 36002 15700 36004
rect 15561 36000 15700 36002
rect 15561 35944 15566 36000
rect 15622 35944 15700 36000
rect 15561 35942 15700 35944
rect 15561 35939 15627 35942
rect 15694 35940 15700 35942
rect 15764 35940 15770 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 1301 35866 1367 35869
rect 19241 35866 19307 35869
rect 1301 35864 19307 35866
rect 1301 35808 1306 35864
rect 1362 35808 19246 35864
rect 19302 35808 19307 35864
rect 1301 35806 19307 35808
rect 1301 35803 1367 35806
rect 19241 35803 19307 35806
rect 7005 35730 7071 35733
rect 8569 35730 8635 35733
rect 9581 35730 9647 35733
rect 7005 35728 9647 35730
rect 7005 35672 7010 35728
rect 7066 35672 8574 35728
rect 8630 35672 9586 35728
rect 9642 35672 9647 35728
rect 7005 35670 9647 35672
rect 7005 35667 7071 35670
rect 8569 35667 8635 35670
rect 9581 35667 9647 35670
rect 12249 35730 12315 35733
rect 12617 35730 12683 35733
rect 12249 35728 12683 35730
rect 12249 35672 12254 35728
rect 12310 35672 12622 35728
rect 12678 35672 12683 35728
rect 12249 35670 12683 35672
rect 12249 35667 12315 35670
rect 12617 35667 12683 35670
rect 3325 35594 3391 35597
rect 12433 35594 12499 35597
rect 13670 35594 13676 35596
rect 3325 35592 13676 35594
rect 3325 35536 3330 35592
rect 3386 35536 12438 35592
rect 12494 35536 13676 35592
rect 3325 35534 13676 35536
rect 3325 35531 3391 35534
rect 12433 35531 12499 35534
rect 13670 35532 13676 35534
rect 13740 35532 13746 35596
rect 200 35368 800 35488
rect 9806 35396 9812 35460
rect 9876 35458 9882 35460
rect 9949 35458 10015 35461
rect 10869 35458 10935 35461
rect 9876 35456 10935 35458
rect 9876 35400 9954 35456
rect 10010 35400 10874 35456
rect 10930 35400 10935 35456
rect 9876 35398 10935 35400
rect 9876 35396 9882 35398
rect 9949 35395 10015 35398
rect 10869 35395 10935 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 8385 35322 8451 35325
rect 11145 35322 11211 35325
rect 8385 35320 11211 35322
rect 8385 35264 8390 35320
rect 8446 35264 11150 35320
rect 11206 35264 11211 35320
rect 8385 35262 11211 35264
rect 8385 35259 8451 35262
rect 11145 35259 11211 35262
rect 10501 35186 10567 35189
rect 17585 35186 17651 35189
rect 10501 35184 17651 35186
rect 10501 35128 10506 35184
rect 10562 35128 17590 35184
rect 17646 35128 17651 35184
rect 10501 35126 17651 35128
rect 10501 35123 10567 35126
rect 17585 35123 17651 35126
rect 3233 35050 3299 35053
rect 3366 35050 3372 35052
rect 3233 35048 3372 35050
rect 3233 34992 3238 35048
rect 3294 34992 3372 35048
rect 3233 34990 3372 34992
rect 3233 34987 3299 34990
rect 3366 34988 3372 34990
rect 3436 34988 3442 35052
rect 10593 35050 10659 35053
rect 14273 35050 14339 35053
rect 10593 35048 14339 35050
rect 10593 34992 10598 35048
rect 10654 34992 14278 35048
rect 14334 34992 14339 35048
rect 10593 34990 14339 34992
rect 10593 34987 10659 34990
rect 14273 34987 14339 34990
rect 3325 34914 3391 34917
rect 3550 34914 3556 34916
rect 3325 34912 3556 34914
rect 3325 34856 3330 34912
rect 3386 34856 3556 34912
rect 3325 34854 3556 34856
rect 3325 34851 3391 34854
rect 3550 34852 3556 34854
rect 3620 34852 3626 34916
rect 9489 34914 9555 34917
rect 11145 34914 11211 34917
rect 13261 34916 13327 34917
rect 13261 34914 13308 34916
rect 9489 34912 11211 34914
rect 9489 34856 9494 34912
rect 9550 34856 11150 34912
rect 11206 34856 11211 34912
rect 9489 34854 11211 34856
rect 13216 34912 13308 34914
rect 13216 34856 13266 34912
rect 13216 34854 13308 34856
rect 9489 34851 9555 34854
rect 11145 34851 11211 34854
rect 13261 34852 13308 34854
rect 13372 34852 13378 34916
rect 13261 34851 13327 34852
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 11145 34778 11211 34781
rect 13721 34778 13787 34781
rect 11145 34776 13787 34778
rect 11145 34720 11150 34776
rect 11206 34720 13726 34776
rect 13782 34720 13787 34776
rect 11145 34718 13787 34720
rect 11145 34715 11211 34718
rect 13721 34715 13787 34718
rect 13997 34778 14063 34781
rect 15009 34778 15075 34781
rect 13997 34776 15075 34778
rect 13997 34720 14002 34776
rect 14058 34720 15014 34776
rect 15070 34720 15075 34776
rect 13997 34718 15075 34720
rect 13997 34715 14063 34718
rect 15009 34715 15075 34718
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 12525 34644 12591 34645
rect 12525 34640 12572 34644
rect 12636 34642 12642 34644
rect 12525 34584 12530 34640
rect 12525 34580 12572 34584
rect 12636 34582 12682 34642
rect 12636 34580 12642 34582
rect 12525 34579 12591 34580
rect 5533 34506 5599 34509
rect 11697 34506 11763 34509
rect 5533 34504 11763 34506
rect 5533 34448 5538 34504
rect 5594 34448 11702 34504
rect 11758 34448 11763 34504
rect 5533 34446 11763 34448
rect 5533 34443 5599 34446
rect 11697 34443 11763 34446
rect 11237 34370 11303 34373
rect 13169 34370 13235 34373
rect 11237 34368 13235 34370
rect 11237 34312 11242 34368
rect 11298 34312 13174 34368
rect 13230 34312 13235 34368
rect 11237 34310 13235 34312
rect 11237 34307 11303 34310
rect 13169 34307 13235 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 6729 34234 6795 34237
rect 11421 34234 11487 34237
rect 6729 34232 11487 34234
rect 6729 34176 6734 34232
rect 6790 34176 11426 34232
rect 11482 34176 11487 34232
rect 6729 34174 11487 34176
rect 6729 34171 6795 34174
rect 11421 34171 11487 34174
rect 11605 34234 11671 34237
rect 12433 34234 12499 34237
rect 11605 34232 12499 34234
rect 11605 34176 11610 34232
rect 11666 34176 12438 34232
rect 12494 34176 12499 34232
rect 11605 34174 12499 34176
rect 11605 34171 11671 34174
rect 12433 34171 12499 34174
rect 3918 34036 3924 34100
rect 3988 34098 3994 34100
rect 8293 34098 8359 34101
rect 3988 34096 8359 34098
rect 3988 34040 8298 34096
rect 8354 34040 8359 34096
rect 3988 34038 8359 34040
rect 3988 34036 3994 34038
rect 8293 34035 8359 34038
rect 8201 33962 8267 33965
rect 15653 33962 15719 33965
rect 8201 33960 15719 33962
rect 8201 33904 8206 33960
rect 8262 33904 15658 33960
rect 15714 33904 15719 33960
rect 8201 33902 15719 33904
rect 8201 33899 8267 33902
rect 15653 33899 15719 33902
rect 11881 33826 11947 33829
rect 15193 33826 15259 33829
rect 11881 33824 15259 33826
rect 11881 33768 11886 33824
rect 11942 33768 15198 33824
rect 15254 33768 15259 33824
rect 11881 33766 15259 33768
rect 11881 33763 11947 33766
rect 15193 33763 15259 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 9765 33690 9831 33693
rect 10593 33690 10659 33693
rect 9765 33688 10659 33690
rect 9765 33632 9770 33688
rect 9826 33632 10598 33688
rect 10654 33632 10659 33688
rect 9765 33630 10659 33632
rect 9765 33627 9831 33630
rect 10593 33627 10659 33630
rect 11605 33690 11671 33693
rect 15929 33690 15995 33693
rect 11605 33688 15995 33690
rect 11605 33632 11610 33688
rect 11666 33632 15934 33688
rect 15990 33632 15995 33688
rect 11605 33630 15995 33632
rect 11605 33627 11671 33630
rect 15929 33627 15995 33630
rect 2313 33554 2379 33557
rect 11094 33554 11100 33556
rect 2313 33552 11100 33554
rect 2313 33496 2318 33552
rect 2374 33496 11100 33552
rect 2313 33494 11100 33496
rect 2313 33491 2379 33494
rect 11094 33492 11100 33494
rect 11164 33492 11170 33556
rect 11513 33554 11579 33557
rect 12617 33554 12683 33557
rect 11513 33552 12683 33554
rect 11513 33496 11518 33552
rect 11574 33496 12622 33552
rect 12678 33496 12683 33552
rect 11513 33494 12683 33496
rect 11513 33491 11579 33494
rect 12617 33491 12683 33494
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 4521 33418 4587 33421
rect 4981 33418 5047 33421
rect 6126 33418 6132 33420
rect 4521 33416 6132 33418
rect 4521 33360 4526 33416
rect 4582 33360 4986 33416
rect 5042 33360 6132 33416
rect 4521 33358 6132 33360
rect 4521 33355 4587 33358
rect 4981 33355 5047 33358
rect 6126 33356 6132 33358
rect 6196 33356 6202 33420
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 6318 33358 12220 33418
rect 4613 33282 4679 33285
rect 6318 33282 6378 33358
rect 4613 33280 6378 33282
rect 4613 33224 4618 33280
rect 4674 33224 6378 33280
rect 4613 33222 6378 33224
rect 6545 33282 6611 33285
rect 9949 33282 10015 33285
rect 10409 33282 10475 33285
rect 6545 33280 10475 33282
rect 6545 33224 6550 33280
rect 6606 33224 9954 33280
rect 10010 33224 10414 33280
rect 10470 33224 10475 33280
rect 6545 33222 10475 33224
rect 12160 33282 12220 33358
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 13537 33282 13603 33285
rect 12160 33280 13603 33282
rect 12160 33224 13542 33280
rect 13598 33224 13603 33280
rect 12160 33222 13603 33224
rect 4613 33219 4679 33222
rect 6545 33219 6611 33222
rect 9949 33219 10015 33222
rect 10409 33219 10475 33222
rect 13537 33219 13603 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 8385 33148 8451 33149
rect 8334 33146 8340 33148
rect 8294 33086 8340 33146
rect 8404 33144 8451 33148
rect 8446 33088 8451 33144
rect 8334 33084 8340 33086
rect 8404 33084 8451 33088
rect 14590 33084 14596 33148
rect 14660 33146 14666 33148
rect 19333 33146 19399 33149
rect 14660 33144 19399 33146
rect 14660 33088 19338 33144
rect 19394 33088 19399 33144
rect 14660 33086 19399 33088
rect 14660 33084 14666 33086
rect 8385 33083 8451 33084
rect 19333 33083 19399 33086
rect 9438 32948 9444 33012
rect 9508 33010 9514 33012
rect 9581 33010 9647 33013
rect 13997 33010 14063 33013
rect 9508 33008 9647 33010
rect 9508 32952 9586 33008
rect 9642 32952 9647 33008
rect 9508 32950 9647 32952
rect 9508 32948 9514 32950
rect 9581 32947 9647 32950
rect 12390 33008 14063 33010
rect 12390 32952 14002 33008
rect 14058 32952 14063 33008
rect 12390 32950 14063 32952
rect 9397 32874 9463 32877
rect 12390 32874 12450 32950
rect 13997 32947 14063 32950
rect 9397 32872 12450 32874
rect 9397 32816 9402 32872
rect 9458 32816 12450 32872
rect 9397 32814 12450 32816
rect 9397 32811 9463 32814
rect 5257 32738 5323 32741
rect 9397 32738 9463 32741
rect 5257 32736 9463 32738
rect 5257 32680 5262 32736
rect 5318 32680 9402 32736
rect 9458 32680 9463 32736
rect 5257 32678 9463 32680
rect 5257 32675 5323 32678
rect 9397 32675 9463 32678
rect 11789 32738 11855 32741
rect 13721 32738 13787 32741
rect 11789 32736 13787 32738
rect 11789 32680 11794 32736
rect 11850 32680 13726 32736
rect 13782 32680 13787 32736
rect 11789 32678 13787 32680
rect 11789 32675 11855 32678
rect 13721 32675 13787 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 10777 32602 10843 32605
rect 15653 32602 15719 32605
rect 10777 32600 15719 32602
rect 10777 32544 10782 32600
rect 10838 32544 15658 32600
rect 15714 32544 15719 32600
rect 10777 32542 15719 32544
rect 10777 32539 10843 32542
rect 15653 32539 15719 32542
rect 12341 32466 12407 32469
rect 2730 32464 12407 32466
rect 2730 32408 12346 32464
rect 12402 32408 12407 32464
rect 2730 32406 12407 32408
rect 200 32058 800 32088
rect 2730 32058 2790 32406
rect 12341 32403 12407 32406
rect 2865 32330 2931 32333
rect 4061 32330 4127 32333
rect 6821 32330 6887 32333
rect 8661 32330 8727 32333
rect 2865 32328 8727 32330
rect 2865 32272 2870 32328
rect 2926 32272 4066 32328
rect 4122 32272 6826 32328
rect 6882 32272 8666 32328
rect 8722 32272 8727 32328
rect 2865 32270 8727 32272
rect 2865 32267 2931 32270
rect 4061 32267 4127 32270
rect 6821 32267 6887 32270
rect 8661 32267 8727 32270
rect 9213 32332 9279 32333
rect 9213 32328 9260 32332
rect 9324 32330 9330 32332
rect 11697 32330 11763 32333
rect 14365 32330 14431 32333
rect 9213 32272 9218 32328
rect 9213 32268 9260 32272
rect 9324 32270 9370 32330
rect 11697 32328 14431 32330
rect 11697 32272 11702 32328
rect 11758 32272 14370 32328
rect 14426 32272 14431 32328
rect 11697 32270 14431 32272
rect 9324 32268 9330 32270
rect 9213 32267 9279 32268
rect 11697 32267 11763 32270
rect 14365 32267 14431 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 200 31998 2790 32058
rect 4797 32058 4863 32061
rect 8109 32058 8175 32061
rect 4797 32056 8175 32058
rect 4797 32000 4802 32056
rect 4858 32000 8114 32056
rect 8170 32000 8175 32056
rect 4797 31998 8175 32000
rect 200 31968 800 31998
rect 4797 31995 4863 31998
rect 8109 31995 8175 31998
rect 9857 32058 9923 32061
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 9857 32056 22110 32058
rect 9857 32000 9862 32056
rect 9918 32000 22110 32056
rect 9857 31998 22110 32000
rect 9857 31995 9923 31998
rect 3734 31860 3740 31924
rect 3804 31922 3810 31924
rect 3969 31922 4035 31925
rect 3804 31920 4035 31922
rect 3804 31864 3974 31920
rect 4030 31864 4035 31920
rect 3804 31862 4035 31864
rect 3804 31860 3810 31862
rect 3969 31859 4035 31862
rect 4521 31922 4587 31925
rect 14365 31922 14431 31925
rect 4521 31920 14431 31922
rect 4521 31864 4526 31920
rect 4582 31864 14370 31920
rect 14426 31864 14431 31920
rect 4521 31862 14431 31864
rect 22050 31922 22110 31998
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 25129 31922 25195 31925
rect 22050 31920 25195 31922
rect 22050 31864 25134 31920
rect 25190 31864 25195 31920
rect 22050 31862 25195 31864
rect 4521 31859 4587 31862
rect 14365 31859 14431 31862
rect 25129 31859 25195 31862
rect 1853 31786 1919 31789
rect 2630 31786 2636 31788
rect 1853 31784 2636 31786
rect 1853 31728 1858 31784
rect 1914 31728 2636 31784
rect 1853 31726 2636 31728
rect 1853 31723 1919 31726
rect 2630 31724 2636 31726
rect 2700 31724 2706 31788
rect 9673 31786 9739 31789
rect 12065 31786 12131 31789
rect 9673 31784 12131 31786
rect 9673 31728 9678 31784
rect 9734 31728 12070 31784
rect 12126 31728 12131 31784
rect 9673 31726 12131 31728
rect 9673 31723 9739 31726
rect 12065 31723 12131 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 10501 31514 10567 31517
rect 12525 31514 12591 31517
rect 10501 31512 12591 31514
rect 10501 31456 10506 31512
rect 10562 31456 12530 31512
rect 12586 31456 12591 31512
rect 10501 31454 12591 31456
rect 10501 31451 10567 31454
rect 12525 31451 12591 31454
rect 9121 31378 9187 31381
rect 10593 31378 10659 31381
rect 13445 31378 13511 31381
rect 9121 31376 10659 31378
rect 9121 31320 9126 31376
rect 9182 31320 10598 31376
rect 10654 31320 10659 31376
rect 9121 31318 10659 31320
rect 9121 31315 9187 31318
rect 10593 31315 10659 31318
rect 12390 31376 13511 31378
rect 12390 31320 13450 31376
rect 13506 31320 13511 31376
rect 12390 31318 13511 31320
rect 4981 31242 5047 31245
rect 12390 31242 12450 31318
rect 13445 31315 13511 31318
rect 4981 31240 12450 31242
rect 4981 31184 4986 31240
rect 5042 31184 12450 31240
rect 4981 31182 12450 31184
rect 4981 31179 5047 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 10409 30836 10475 30837
rect 10358 30834 10364 30836
rect 10318 30774 10364 30834
rect 10428 30832 10475 30836
rect 10470 30776 10475 30832
rect 10358 30772 10364 30774
rect 10428 30772 10475 30776
rect 10409 30771 10475 30772
rect 10685 30834 10751 30837
rect 15561 30834 15627 30837
rect 10685 30832 15627 30834
rect 10685 30776 10690 30832
rect 10746 30776 15566 30832
rect 15622 30776 15627 30832
rect 10685 30774 15627 30776
rect 10685 30771 10751 30774
rect 15561 30771 15627 30774
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 4654 30636 4660 30700
rect 4724 30698 4730 30700
rect 5165 30698 5231 30701
rect 24393 30698 24459 30701
rect 4724 30696 24459 30698
rect 4724 30640 5170 30696
rect 5226 30640 24398 30696
rect 24454 30640 24459 30696
rect 4724 30638 24459 30640
rect 4724 30636 4730 30638
rect 5165 30635 5231 30638
rect 24393 30635 24459 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 2446 30364 2452 30428
rect 2516 30426 2522 30428
rect 4521 30426 4587 30429
rect 5022 30426 5028 30428
rect 2516 30424 5028 30426
rect 2516 30368 4526 30424
rect 4582 30368 5028 30424
rect 2516 30366 5028 30368
rect 2516 30364 2522 30366
rect 4521 30363 4587 30366
rect 5022 30364 5028 30366
rect 5092 30364 5098 30428
rect 10869 30426 10935 30429
rect 13445 30426 13511 30429
rect 10869 30424 13511 30426
rect 10869 30368 10874 30424
rect 10930 30368 13450 30424
rect 13506 30368 13511 30424
rect 10869 30366 13511 30368
rect 10869 30363 10935 30366
rect 13445 30363 13511 30366
rect 5441 30290 5507 30293
rect 15009 30290 15075 30293
rect 5441 30288 15075 30290
rect 5441 30232 5446 30288
rect 5502 30232 15014 30288
rect 15070 30232 15075 30288
rect 5441 30230 15075 30232
rect 5441 30227 5507 30230
rect 15009 30227 15075 30230
rect 5073 30154 5139 30157
rect 5390 30154 5396 30156
rect 5073 30152 5396 30154
rect 5073 30096 5078 30152
rect 5134 30096 5396 30152
rect 5073 30094 5396 30096
rect 5073 30091 5139 30094
rect 5390 30092 5396 30094
rect 5460 30092 5466 30156
rect 10133 30154 10199 30157
rect 16941 30154 17007 30157
rect 10133 30152 17007 30154
rect 10133 30096 10138 30152
rect 10194 30096 16946 30152
rect 17002 30096 17007 30152
rect 10133 30094 17007 30096
rect 10133 30091 10199 30094
rect 16941 30091 17007 30094
rect 8201 30018 8267 30021
rect 10358 30018 10364 30020
rect 8201 30016 10364 30018
rect 8201 29960 8206 30016
rect 8262 29960 10364 30016
rect 8201 29958 10364 29960
rect 8201 29955 8267 29958
rect 10358 29956 10364 29958
rect 10428 30018 10434 30020
rect 12065 30018 12131 30021
rect 10428 30016 12131 30018
rect 10428 29960 12070 30016
rect 12126 29960 12131 30016
rect 10428 29958 12131 29960
rect 10428 29956 10434 29958
rect 12065 29955 12131 29958
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 7465 29746 7531 29749
rect 17769 29746 17835 29749
rect 7465 29744 17835 29746
rect 7465 29688 7470 29744
rect 7526 29688 17774 29744
rect 17830 29688 17835 29744
rect 7465 29686 17835 29688
rect 7465 29683 7531 29686
rect 17769 29683 17835 29686
rect 19517 29746 19583 29749
rect 21633 29746 21699 29749
rect 19517 29744 21699 29746
rect 19517 29688 19522 29744
rect 19578 29688 21638 29744
rect 21694 29688 21699 29744
rect 19517 29686 21699 29688
rect 19517 29683 19583 29686
rect 21633 29683 21699 29686
rect 1853 29612 1919 29613
rect 1853 29610 1900 29612
rect 1808 29608 1900 29610
rect 1808 29552 1858 29608
rect 1808 29550 1900 29552
rect 1853 29548 1900 29550
rect 1964 29548 1970 29612
rect 4521 29610 4587 29613
rect 4654 29610 4660 29612
rect 4521 29608 4660 29610
rect 4521 29552 4526 29608
rect 4582 29552 4660 29608
rect 4521 29550 4660 29552
rect 1853 29547 1919 29548
rect 4521 29547 4587 29550
rect 4654 29548 4660 29550
rect 4724 29548 4730 29612
rect 9121 29610 9187 29613
rect 9765 29610 9831 29613
rect 19609 29610 19675 29613
rect 9121 29608 9831 29610
rect 9121 29552 9126 29608
rect 9182 29552 9770 29608
rect 9826 29552 9831 29608
rect 9121 29550 9831 29552
rect 9121 29547 9187 29550
rect 9765 29547 9831 29550
rect 19382 29608 19675 29610
rect 19382 29552 19614 29608
rect 19670 29552 19675 29608
rect 19382 29550 19675 29552
rect 9397 29338 9463 29341
rect 9949 29338 10015 29341
rect 9397 29336 10015 29338
rect 9397 29280 9402 29336
rect 9458 29280 9954 29336
rect 10010 29280 10015 29336
rect 9397 29278 10015 29280
rect 9397 29275 9463 29278
rect 9949 29275 10015 29278
rect 10593 29338 10659 29341
rect 11646 29338 11652 29340
rect 10593 29336 11652 29338
rect 10593 29280 10598 29336
rect 10654 29280 11652 29336
rect 10593 29278 11652 29280
rect 10593 29275 10659 29278
rect 11646 29276 11652 29278
rect 11716 29276 11722 29340
rect 7741 29202 7807 29205
rect 12893 29202 12959 29205
rect 7741 29200 12959 29202
rect 7741 29144 7746 29200
rect 7802 29144 12898 29200
rect 12954 29144 12959 29200
rect 7741 29142 12959 29144
rect 19382 29202 19442 29550
rect 19609 29547 19675 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 19517 29202 19583 29205
rect 19382 29200 19583 29202
rect 19382 29144 19522 29200
rect 19578 29144 19583 29200
rect 19382 29142 19583 29144
rect 7741 29139 7807 29142
rect 12893 29139 12959 29142
rect 19517 29139 19583 29142
rect 3785 29066 3851 29069
rect 5574 29066 5580 29068
rect 3785 29064 5580 29066
rect 3785 29008 3790 29064
rect 3846 29008 5580 29064
rect 3785 29006 5580 29008
rect 3785 29003 3851 29006
rect 5574 29004 5580 29006
rect 5644 29004 5650 29068
rect 8753 29066 8819 29069
rect 11973 29066 12039 29069
rect 8753 29064 12039 29066
rect 8753 29008 8758 29064
rect 8814 29008 11978 29064
rect 12034 29008 12039 29064
rect 8753 29006 12039 29008
rect 8753 29003 8819 29006
rect 11973 29003 12039 29006
rect 12249 29066 12315 29069
rect 13169 29066 13235 29069
rect 12249 29064 13235 29066
rect 12249 29008 12254 29064
rect 12310 29008 13174 29064
rect 13230 29008 13235 29064
rect 12249 29006 13235 29008
rect 12249 29003 12315 29006
rect 13169 29003 13235 29006
rect 2313 28930 2379 28933
rect 2446 28930 2452 28932
rect 2313 28928 2452 28930
rect 2313 28872 2318 28928
rect 2374 28872 2452 28928
rect 2313 28870 2452 28872
rect 2313 28867 2379 28870
rect 2446 28868 2452 28870
rect 2516 28868 2522 28932
rect 10777 28930 10843 28933
rect 10910 28930 10916 28932
rect 10777 28928 10916 28930
rect 10777 28872 10782 28928
rect 10838 28872 10916 28928
rect 10777 28870 10916 28872
rect 10777 28867 10843 28870
rect 10910 28868 10916 28870
rect 10980 28868 10986 28932
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 9857 28794 9923 28797
rect 10961 28794 11027 28797
rect 11421 28794 11487 28797
rect 9857 28792 11027 28794
rect 9857 28736 9862 28792
rect 9918 28736 10966 28792
rect 11022 28736 11027 28792
rect 9857 28734 11027 28736
rect 9857 28731 9923 28734
rect 10961 28731 11027 28734
rect 11286 28792 11487 28794
rect 11286 28736 11426 28792
rect 11482 28736 11487 28792
rect 11286 28734 11487 28736
rect 200 28658 800 28688
rect 3141 28658 3207 28661
rect 200 28656 3207 28658
rect 200 28600 3146 28656
rect 3202 28600 3207 28656
rect 200 28598 3207 28600
rect 200 28568 800 28598
rect 3141 28595 3207 28598
rect 4429 28658 4495 28661
rect 11286 28658 11346 28734
rect 11421 28731 11487 28734
rect 4429 28656 11346 28658
rect 4429 28600 4434 28656
rect 4490 28600 11346 28656
rect 4429 28598 11346 28600
rect 4429 28595 4495 28598
rect 11462 28596 11468 28660
rect 11532 28658 11538 28660
rect 21909 28658 21975 28661
rect 11532 28656 21975 28658
rect 11532 28600 21914 28656
rect 21970 28600 21975 28656
rect 11532 28598 21975 28600
rect 11532 28596 11538 28598
rect 21909 28595 21975 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 10041 28522 10107 28525
rect 11697 28522 11763 28525
rect 10041 28520 11763 28522
rect 10041 28464 10046 28520
rect 10102 28464 11702 28520
rect 11758 28464 11763 28520
rect 10041 28462 11763 28464
rect 10041 28459 10107 28462
rect 11697 28459 11763 28462
rect 4337 28386 4403 28389
rect 8334 28386 8340 28388
rect 4337 28384 8340 28386
rect 4337 28328 4342 28384
rect 4398 28328 8340 28384
rect 4337 28326 8340 28328
rect 4337 28323 4403 28326
rect 8334 28324 8340 28326
rect 8404 28386 8410 28388
rect 9622 28386 9628 28388
rect 8404 28326 9628 28386
rect 8404 28324 8410 28326
rect 9622 28324 9628 28326
rect 9692 28324 9698 28388
rect 10317 28386 10383 28389
rect 10593 28386 10659 28389
rect 10317 28384 10659 28386
rect 10317 28328 10322 28384
rect 10378 28328 10598 28384
rect 10654 28328 10659 28384
rect 10317 28326 10659 28328
rect 10317 28323 10383 28326
rect 10593 28323 10659 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 2630 28188 2636 28252
rect 2700 28250 2706 28252
rect 3785 28250 3851 28253
rect 2700 28248 3851 28250
rect 2700 28192 3790 28248
rect 3846 28192 3851 28248
rect 2700 28190 3851 28192
rect 2700 28188 2706 28190
rect 3785 28187 3851 28190
rect 3969 28250 4035 28253
rect 10685 28250 10751 28253
rect 11421 28250 11487 28253
rect 3969 28248 11487 28250
rect 3969 28192 3974 28248
rect 4030 28192 10690 28248
rect 10746 28192 11426 28248
rect 11482 28192 11487 28248
rect 3969 28190 11487 28192
rect 3969 28187 4035 28190
rect 10685 28187 10751 28190
rect 11421 28187 11487 28190
rect 1853 28114 1919 28117
rect 2681 28114 2747 28117
rect 16849 28114 16915 28117
rect 1853 28112 16915 28114
rect 1853 28056 1858 28112
rect 1914 28056 2686 28112
rect 2742 28056 16854 28112
rect 16910 28056 16915 28112
rect 1853 28054 16915 28056
rect 1853 28051 1919 28054
rect 2681 28051 2747 28054
rect 16849 28051 16915 28054
rect 2405 27978 2471 27981
rect 8334 27978 8340 27980
rect 2405 27976 8340 27978
rect 2405 27920 2410 27976
rect 2466 27920 8340 27976
rect 2405 27918 8340 27920
rect 2405 27915 2471 27918
rect 8334 27916 8340 27918
rect 8404 27916 8410 27980
rect 8937 27978 9003 27981
rect 13445 27978 13511 27981
rect 8937 27976 13511 27978
rect 8937 27920 8942 27976
rect 8998 27920 13450 27976
rect 13506 27920 13511 27976
rect 8937 27918 13511 27920
rect 8937 27915 9003 27918
rect 13445 27915 13511 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 1853 27706 1919 27709
rect 2078 27706 2084 27708
rect 1853 27704 2084 27706
rect 1853 27648 1858 27704
rect 1914 27648 2084 27704
rect 1853 27646 2084 27648
rect 1853 27643 1919 27646
rect 2078 27644 2084 27646
rect 2148 27644 2154 27708
rect 7414 27644 7420 27708
rect 7484 27706 7490 27708
rect 7649 27706 7715 27709
rect 7484 27704 7715 27706
rect 7484 27648 7654 27704
rect 7710 27648 7715 27704
rect 7484 27646 7715 27648
rect 7484 27644 7490 27646
rect 7649 27643 7715 27646
rect 3601 27570 3667 27573
rect 3918 27570 3924 27572
rect 3601 27568 3924 27570
rect 3601 27512 3606 27568
rect 3662 27512 3924 27568
rect 3601 27510 3924 27512
rect 3601 27507 3667 27510
rect 3918 27508 3924 27510
rect 3988 27508 3994 27572
rect 7230 27508 7236 27572
rect 7300 27570 7306 27572
rect 11462 27570 11468 27572
rect 7300 27510 11468 27570
rect 7300 27508 7306 27510
rect 11462 27508 11468 27510
rect 11532 27508 11538 27572
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 3417 27026 3483 27029
rect 4613 27026 4679 27029
rect 17953 27026 18019 27029
rect 3417 27024 18019 27026
rect 3417 26968 3422 27024
rect 3478 26968 4618 27024
rect 4674 26968 17958 27024
rect 18014 26968 18019 27024
rect 3417 26966 18019 26968
rect 3417 26963 3483 26966
rect 4613 26963 4679 26966
rect 17953 26963 18019 26966
rect 3601 26890 3667 26893
rect 7230 26890 7236 26892
rect 3601 26888 7236 26890
rect 3601 26832 3606 26888
rect 3662 26832 7236 26888
rect 3601 26830 7236 26832
rect 3601 26827 3667 26830
rect 7230 26828 7236 26830
rect 7300 26828 7306 26892
rect 8845 26890 8911 26893
rect 11145 26890 11211 26893
rect 8845 26888 11211 26890
rect 8845 26832 8850 26888
rect 8906 26832 11150 26888
rect 11206 26832 11211 26888
rect 8845 26830 11211 26832
rect 8845 26827 8911 26830
rect 11145 26827 11211 26830
rect 15469 26890 15535 26893
rect 17585 26890 17651 26893
rect 15469 26888 17651 26890
rect 15469 26832 15474 26888
rect 15530 26832 17590 26888
rect 17646 26832 17651 26888
rect 15469 26830 17651 26832
rect 15469 26827 15535 26830
rect 17585 26827 17651 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 6545 26618 6611 26621
rect 9581 26618 9647 26621
rect 6545 26616 9647 26618
rect 6545 26560 6550 26616
rect 6606 26560 9586 26616
rect 9642 26560 9647 26616
rect 6545 26558 9647 26560
rect 6545 26555 6611 26558
rect 9581 26555 9647 26558
rect 12157 26618 12223 26621
rect 12433 26618 12499 26621
rect 12157 26616 12499 26618
rect 12157 26560 12162 26616
rect 12218 26560 12438 26616
rect 12494 26560 12499 26616
rect 12157 26558 12499 26560
rect 12157 26555 12223 26558
rect 12433 26555 12499 26558
rect 13905 26618 13971 26621
rect 16757 26618 16823 26621
rect 13905 26616 16823 26618
rect 13905 26560 13910 26616
rect 13966 26560 16762 26616
rect 16818 26560 16823 26616
rect 13905 26558 16823 26560
rect 13905 26555 13971 26558
rect 16757 26555 16823 26558
rect 6177 26482 6243 26485
rect 15009 26482 15075 26485
rect 6177 26480 15075 26482
rect 6177 26424 6182 26480
rect 6238 26424 15014 26480
rect 15070 26424 15075 26480
rect 6177 26422 15075 26424
rect 6177 26419 6243 26422
rect 15009 26419 15075 26422
rect 7925 26346 7991 26349
rect 11278 26346 11284 26348
rect 7925 26344 11284 26346
rect 7925 26288 7930 26344
rect 7986 26288 11284 26344
rect 7925 26286 11284 26288
rect 7925 26283 7991 26286
rect 11278 26284 11284 26286
rect 11348 26284 11354 26348
rect 12157 26346 12223 26349
rect 14733 26346 14799 26349
rect 12157 26344 14799 26346
rect 12157 26288 12162 26344
rect 12218 26288 14738 26344
rect 14794 26288 14799 26344
rect 12157 26286 14799 26288
rect 12157 26283 12223 26286
rect 14733 26283 14799 26286
rect 8334 26148 8340 26212
rect 8404 26210 8410 26212
rect 8937 26210 9003 26213
rect 8404 26208 9003 26210
rect 8404 26152 8942 26208
rect 8998 26152 9003 26208
rect 8404 26150 9003 26152
rect 8404 26148 8410 26150
rect 8937 26147 9003 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 10317 26074 10383 26077
rect 15561 26074 15627 26077
rect 17585 26074 17651 26077
rect 10317 26072 17651 26074
rect 10317 26016 10322 26072
rect 10378 26016 15566 26072
rect 15622 26016 17590 26072
rect 17646 26016 17651 26072
rect 10317 26014 17651 26016
rect 10317 26011 10383 26014
rect 15561 26011 15627 26014
rect 17585 26011 17651 26014
rect 9121 25938 9187 25941
rect 13353 25938 13419 25941
rect 9121 25936 13419 25938
rect 9121 25880 9126 25936
rect 9182 25880 13358 25936
rect 13414 25880 13419 25936
rect 9121 25878 13419 25880
rect 9121 25875 9187 25878
rect 13353 25875 13419 25878
rect 3734 25740 3740 25804
rect 3804 25802 3810 25804
rect 10961 25802 11027 25805
rect 3804 25800 11027 25802
rect 3804 25744 10966 25800
rect 11022 25744 11027 25800
rect 3804 25742 11027 25744
rect 3804 25740 3810 25742
rect 10961 25739 11027 25742
rect 7281 25666 7347 25669
rect 13077 25666 13143 25669
rect 7281 25664 13143 25666
rect 7281 25608 7286 25664
rect 7342 25608 13082 25664
rect 13138 25608 13143 25664
rect 7281 25606 13143 25608
rect 7281 25603 7347 25606
rect 13077 25603 13143 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 5717 25530 5783 25533
rect 13813 25530 13879 25533
rect 5717 25528 13879 25530
rect 5717 25472 5722 25528
rect 5778 25472 13818 25528
rect 13874 25472 13879 25528
rect 5717 25470 13879 25472
rect 5717 25467 5783 25470
rect 13813 25467 13879 25470
rect 3969 25394 4035 25397
rect 9254 25394 9260 25396
rect 3969 25392 9260 25394
rect 3969 25336 3974 25392
rect 4030 25336 9260 25392
rect 3969 25334 9260 25336
rect 3969 25331 4035 25334
rect 9254 25332 9260 25334
rect 9324 25332 9330 25396
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 9305 25258 9371 25261
rect 13486 25258 13492 25260
rect 9305 25256 13492 25258
rect 9305 25200 9310 25256
rect 9366 25200 13492 25256
rect 9305 25198 13492 25200
rect 9305 25195 9371 25198
rect 13486 25196 13492 25198
rect 13556 25196 13562 25260
rect 24577 25258 24643 25261
rect 17174 25256 24643 25258
rect 17174 25200 24582 25256
rect 24638 25200 24643 25256
rect 17174 25198 24643 25200
rect 5073 25122 5139 25125
rect 17174 25122 17234 25198
rect 24577 25195 24643 25198
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 5073 25120 17234 25122
rect 5073 25064 5078 25120
rect 5134 25064 17234 25120
rect 5073 25062 17234 25064
rect 5073 25059 5139 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 8293 24986 8359 24989
rect 15694 24986 15700 24988
rect 8293 24984 15700 24986
rect 8293 24928 8298 24984
rect 8354 24928 15700 24984
rect 8293 24926 15700 24928
rect 8293 24923 8359 24926
rect 15694 24924 15700 24926
rect 15764 24924 15770 24988
rect 5533 24850 5599 24853
rect 14590 24850 14596 24852
rect 5533 24848 14596 24850
rect 5533 24792 5538 24848
rect 5594 24792 14596 24848
rect 5533 24790 14596 24792
rect 5533 24787 5599 24790
rect 14590 24788 14596 24790
rect 14660 24788 14666 24852
rect 4061 24714 4127 24717
rect 4838 24714 4844 24716
rect 4061 24712 4844 24714
rect 4061 24656 4066 24712
rect 4122 24656 4844 24712
rect 4061 24654 4844 24656
rect 4061 24651 4127 24654
rect 4838 24652 4844 24654
rect 4908 24652 4914 24716
rect 5574 24652 5580 24716
rect 5644 24714 5650 24716
rect 7557 24714 7623 24717
rect 5644 24712 7623 24714
rect 5644 24656 7562 24712
rect 7618 24656 7623 24712
rect 5644 24654 7623 24656
rect 5644 24652 5650 24654
rect 7557 24651 7623 24654
rect 7741 24578 7807 24581
rect 9857 24578 9923 24581
rect 7741 24576 9923 24578
rect 7741 24520 7746 24576
rect 7802 24520 9862 24576
rect 9918 24520 9923 24576
rect 7741 24518 9923 24520
rect 7741 24515 7807 24518
rect 9857 24515 9923 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 8753 24442 8819 24445
rect 9581 24442 9647 24445
rect 8753 24440 9647 24442
rect 8753 24384 8758 24440
rect 8814 24384 9586 24440
rect 9642 24384 9647 24440
rect 8753 24382 9647 24384
rect 8753 24379 8819 24382
rect 9581 24379 9647 24382
rect 10961 24306 11027 24309
rect 12341 24306 12407 24309
rect 10961 24304 12407 24306
rect 10961 24248 10966 24304
rect 11022 24248 12346 24304
rect 12402 24248 12407 24304
rect 10961 24246 12407 24248
rect 10961 24243 11027 24246
rect 12341 24243 12407 24246
rect 19701 24306 19767 24309
rect 37917 24306 37983 24309
rect 19701 24304 37983 24306
rect 19701 24248 19706 24304
rect 19762 24248 37922 24304
rect 37978 24248 37983 24304
rect 19701 24246 37983 24248
rect 19701 24243 19767 24246
rect 37917 24243 37983 24246
rect 5758 24108 5764 24172
rect 5828 24170 5834 24172
rect 13445 24170 13511 24173
rect 5828 24168 13511 24170
rect 5828 24112 13450 24168
rect 13506 24112 13511 24168
rect 5828 24110 13511 24112
rect 5828 24108 5834 24110
rect 13445 24107 13511 24110
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 3601 23898 3667 23901
rect 5206 23898 5212 23900
rect 3601 23896 5212 23898
rect 3601 23840 3606 23896
rect 3662 23840 5212 23896
rect 3601 23838 5212 23840
rect 3601 23835 3667 23838
rect 5206 23836 5212 23838
rect 5276 23836 5282 23900
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 11646 23292 11652 23356
rect 11716 23354 11722 23356
rect 12157 23354 12223 23357
rect 11716 23352 12223 23354
rect 11716 23296 12162 23352
rect 12218 23296 12223 23352
rect 11716 23294 12223 23296
rect 11716 23292 11722 23294
rect 12157 23291 12223 23294
rect 11278 23156 11284 23220
rect 11348 23218 11354 23220
rect 14365 23218 14431 23221
rect 11348 23216 14431 23218
rect 11348 23160 14370 23216
rect 14426 23160 14431 23216
rect 11348 23158 14431 23160
rect 11348 23156 11354 23158
rect 14365 23155 14431 23158
rect 2313 23082 2379 23085
rect 12566 23082 12572 23084
rect 2313 23080 12572 23082
rect 2313 23024 2318 23080
rect 2374 23024 12572 23080
rect 2313 23022 12572 23024
rect 2313 23019 2379 23022
rect 12566 23020 12572 23022
rect 12636 23020 12642 23084
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 5022 22748 5028 22812
rect 5092 22810 5098 22812
rect 16481 22810 16547 22813
rect 5092 22808 16547 22810
rect 5092 22752 16486 22808
rect 16542 22752 16547 22808
rect 5092 22750 16547 22752
rect 5092 22748 5098 22750
rect 16481 22747 16547 22750
rect 9622 22612 9628 22676
rect 9692 22674 9698 22676
rect 15469 22674 15535 22677
rect 9692 22672 15535 22674
rect 9692 22616 15474 22672
rect 15530 22616 15535 22672
rect 9692 22614 15535 22616
rect 9692 22612 9698 22614
rect 15469 22611 15535 22614
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 10501 22538 10567 22541
rect 12249 22538 12315 22541
rect 10501 22536 12315 22538
rect 10501 22480 10506 22536
rect 10562 22480 12254 22536
rect 12310 22480 12315 22536
rect 10501 22478 12315 22480
rect 10501 22475 10567 22478
rect 12249 22475 12315 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 7649 22266 7715 22269
rect 13537 22266 13603 22269
rect 7649 22264 13603 22266
rect 7649 22208 7654 22264
rect 7710 22208 13542 22264
rect 13598 22208 13603 22264
rect 7649 22206 13603 22208
rect 7649 22203 7715 22206
rect 13537 22203 13603 22206
rect 10317 22130 10383 22133
rect 11053 22130 11119 22133
rect 10317 22128 11119 22130
rect 10317 22072 10322 22128
rect 10378 22072 11058 22128
rect 11114 22072 11119 22128
rect 10317 22070 11119 22072
rect 10317 22067 10383 22070
rect 11053 22067 11119 22070
rect 11646 22068 11652 22132
rect 11716 22130 11722 22132
rect 11716 22070 12266 22130
rect 11716 22068 11722 22070
rect 12206 21997 12266 22070
rect 9213 21994 9279 21997
rect 9857 21994 9923 21997
rect 9213 21992 9923 21994
rect 9213 21936 9218 21992
rect 9274 21936 9862 21992
rect 9918 21936 9923 21992
rect 9213 21934 9923 21936
rect 9213 21931 9279 21934
rect 9857 21931 9923 21934
rect 10501 21994 10567 21997
rect 11605 21994 11671 21997
rect 10501 21992 11671 21994
rect 10501 21936 10506 21992
rect 10562 21936 11610 21992
rect 11666 21936 11671 21992
rect 10501 21934 11671 21936
rect 12206 21992 12315 21997
rect 12206 21936 12254 21992
rect 12310 21936 12315 21992
rect 12206 21934 12315 21936
rect 10501 21931 10567 21934
rect 11605 21931 11671 21934
rect 12249 21931 12315 21934
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 11697 21450 11763 21453
rect 14549 21450 14615 21453
rect 11697 21448 14615 21450
rect 11697 21392 11702 21448
rect 11758 21392 14554 21448
rect 14610 21392 14615 21448
rect 11697 21390 14615 21392
rect 11697 21387 11763 21390
rect 14549 21387 14615 21390
rect 6126 21252 6132 21316
rect 6196 21314 6202 21316
rect 24577 21314 24643 21317
rect 6196 21312 24643 21314
rect 6196 21256 24582 21312
rect 24638 21256 24643 21312
rect 6196 21254 24643 21256
rect 6196 21252 6202 21254
rect 24577 21251 24643 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 9581 20906 9647 20909
rect 13353 20906 13419 20909
rect 9581 20904 13419 20906
rect 9581 20848 9586 20904
rect 9642 20848 13358 20904
rect 13414 20848 13419 20904
rect 9581 20846 13419 20848
rect 9581 20843 9647 20846
rect 13353 20843 13419 20846
rect 9397 20770 9463 20773
rect 11237 20770 11303 20773
rect 9397 20768 11303 20770
rect 9397 20712 9402 20768
rect 9458 20712 11242 20768
rect 11298 20712 11303 20768
rect 9397 20710 11303 20712
rect 9397 20707 9463 20710
rect 11237 20707 11303 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 11053 20498 11119 20501
rect 15469 20498 15535 20501
rect 11053 20496 15535 20498
rect 11053 20440 11058 20496
rect 11114 20440 15474 20496
rect 15530 20440 15535 20496
rect 11053 20438 15535 20440
rect 11053 20435 11119 20438
rect 15469 20435 15535 20438
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 9121 19410 9187 19413
rect 10961 19412 11027 19413
rect 10910 19410 10916 19412
rect 9121 19408 10916 19410
rect 10980 19410 11027 19412
rect 10980 19408 11072 19410
rect 9121 19352 9126 19408
rect 9182 19352 10916 19408
rect 11022 19352 11072 19408
rect 9121 19350 10916 19352
rect 9121 19347 9187 19350
rect 10910 19348 10916 19350
rect 10980 19350 11072 19352
rect 10980 19348 11027 19350
rect 10961 19347 11027 19348
rect 10133 19274 10199 19277
rect 11329 19274 11395 19277
rect 13302 19274 13308 19276
rect 10133 19272 10242 19274
rect 10133 19216 10138 19272
rect 10194 19216 10242 19272
rect 10133 19211 10242 19216
rect 11329 19272 13308 19274
rect 11329 19216 11334 19272
rect 11390 19216 13308 19272
rect 11329 19214 13308 19216
rect 11329 19211 11395 19214
rect 13302 19212 13308 19214
rect 13372 19212 13378 19276
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 9673 19138 9739 19141
rect 10182 19138 10242 19211
rect 14365 19138 14431 19141
rect 9673 19136 14431 19138
rect 9673 19080 9678 19136
rect 9734 19080 14370 19136
rect 14426 19080 14431 19136
rect 9673 19078 14431 19080
rect 9673 19075 9739 19078
rect 14365 19075 14431 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19168
rect 34930 19007 35246 19008
rect 8518 18940 8524 19004
rect 8588 19002 8594 19004
rect 13721 19002 13787 19005
rect 8588 19000 13787 19002
rect 8588 18944 13726 19000
rect 13782 18944 13787 19000
rect 8588 18942 13787 18944
rect 8588 18940 8594 18942
rect 13721 18939 13787 18942
rect 10041 18866 10107 18869
rect 11094 18866 11100 18868
rect 10041 18864 11100 18866
rect 10041 18808 10046 18864
rect 10102 18808 11100 18864
rect 10041 18806 11100 18808
rect 10041 18803 10107 18806
rect 11094 18804 11100 18806
rect 11164 18866 11170 18868
rect 12617 18866 12683 18869
rect 11164 18864 12683 18866
rect 11164 18808 12622 18864
rect 12678 18808 12683 18864
rect 11164 18806 12683 18808
rect 11164 18804 11170 18806
rect 12617 18803 12683 18806
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 8385 18050 8451 18053
rect 9806 18050 9812 18052
rect 8385 18048 9812 18050
rect 8385 17992 8390 18048
rect 8446 17992 9812 18048
rect 8385 17990 9812 17992
rect 8385 17987 8451 17990
rect 9806 17988 9812 17990
rect 9876 17988 9882 18052
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 3550 17716 3556 17780
rect 3620 17778 3626 17780
rect 18689 17778 18755 17781
rect 3620 17776 18755 17778
rect 3620 17720 18694 17776
rect 18750 17720 18755 17776
rect 3620 17718 18755 17720
rect 3620 17716 3626 17718
rect 18689 17715 18755 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 9438 16900 9444 16964
rect 9508 16962 9514 16964
rect 14365 16962 14431 16965
rect 9508 16960 14431 16962
rect 9508 16904 14370 16960
rect 14426 16904 14431 16960
rect 9508 16902 14431 16904
rect 9508 16900 9514 16902
rect 14365 16899 14431 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 3366 15948 3372 16012
rect 3436 16010 3442 16012
rect 12341 16010 12407 16013
rect 15142 16010 15148 16012
rect 3436 16008 15148 16010
rect 3436 15952 12346 16008
rect 12402 15952 15148 16008
rect 3436 15950 15148 15952
rect 3436 15948 3442 15950
rect 12341 15947 12407 15950
rect 15142 15948 15148 15950
rect 15212 15948 15218 16012
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 13721 14516 13787 14517
rect 13670 14452 13676 14516
rect 13740 14514 13787 14516
rect 13740 14512 13832 14514
rect 13782 14456 13832 14512
rect 13740 14454 13832 14456
rect 13740 14452 13787 14454
rect 13721 14451 13787 14452
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 5390 13908 5396 13972
rect 5460 13970 5466 13972
rect 17033 13970 17099 13973
rect 5460 13968 17099 13970
rect 5460 13912 17038 13968
rect 17094 13912 17099 13968
rect 5460 13910 17099 13912
rect 5460 13908 5466 13910
rect 17033 13907 17099 13910
rect 15193 13700 15259 13701
rect 15142 13698 15148 13700
rect 15102 13638 15148 13698
rect 15212 13696 15259 13700
rect 15254 13640 15259 13696
rect 15142 13636 15148 13638
rect 15212 13636 15259 13640
rect 15193 13635 15259 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 7414 6156 7420 6220
rect 7484 6218 7490 6220
rect 37273 6218 37339 6221
rect 7484 6216 37339 6218
rect 7484 6160 37278 6216
rect 37334 6160 37339 6216
rect 7484 6158 37339 6160
rect 7484 6156 7490 6158
rect 37273 6155 37339 6158
rect 38101 6218 38167 6221
rect 39200 6218 39800 6248
rect 38101 6216 39800 6218
rect 38101 6160 38106 6216
rect 38162 6160 39800 6216
rect 38101 6158 39800 6160
rect 38101 6155 38167 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 1853 5404 1919 5405
rect 1853 5402 1900 5404
rect 1808 5400 1900 5402
rect 1808 5344 1858 5400
rect 1808 5342 1900 5344
rect 1853 5340 1900 5342
rect 1964 5340 1970 5404
rect 1853 5339 1919 5340
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2848
rect 1761 2818 1827 2821
rect 200 2816 1827 2818
rect 200 2760 1766 2816
rect 1822 2760 1827 2816
rect 200 2758 1827 2760
rect 200 2728 800 2758
rect 1761 2755 1827 2758
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1761 1458 1827 1461
rect 200 1456 1827 1458
rect 200 1400 1766 1456
rect 1822 1400 1827 1456
rect 200 1398 1827 1400
rect 200 1368 800 1398
rect 1761 1395 1827 1398
rect 36905 1458 36971 1461
rect 39200 1458 39800 1488
rect 36905 1456 39800 1458
rect 36905 1400 36910 1456
rect 36966 1400 39800 1456
rect 36905 1398 39800 1400
rect 36905 1395 36971 1398
rect 39200 1368 39800 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 5764 37088 5828 37092
rect 5764 37032 5778 37088
rect 5778 37032 5828 37088
rect 5764 37028 5828 37032
rect 8524 37088 8588 37092
rect 8524 37032 8538 37088
rect 8538 37032 8588 37088
rect 8524 37028 8588 37032
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 8524 36484 8588 36548
rect 13492 36484 13556 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 2084 36212 2148 36276
rect 5212 36076 5276 36140
rect 11100 36136 11164 36140
rect 11100 36080 11150 36136
rect 11150 36080 11164 36136
rect 11100 36076 11164 36080
rect 4844 36000 4908 36004
rect 4844 35944 4858 36000
rect 4858 35944 4908 36000
rect 4844 35940 4908 35944
rect 7236 36000 7300 36004
rect 7236 35944 7286 36000
rect 7286 35944 7300 36000
rect 7236 35940 7300 35944
rect 15700 35940 15764 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 13676 35532 13740 35596
rect 9812 35396 9876 35460
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 3372 34988 3436 35052
rect 3556 34852 3620 34916
rect 13308 34912 13372 34916
rect 13308 34856 13322 34912
rect 13322 34856 13372 34912
rect 13308 34852 13372 34856
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 12572 34640 12636 34644
rect 12572 34584 12586 34640
rect 12586 34584 12636 34640
rect 12572 34580 12636 34584
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 3924 34036 3988 34100
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 11100 33492 11164 33556
rect 6132 33356 6196 33420
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 8340 33144 8404 33148
rect 8340 33088 8390 33144
rect 8390 33088 8404 33144
rect 8340 33084 8404 33088
rect 14596 33084 14660 33148
rect 9444 32948 9508 33012
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 9260 32328 9324 32332
rect 9260 32272 9274 32328
rect 9274 32272 9324 32328
rect 9260 32268 9324 32272
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 3740 31860 3804 31924
rect 2636 31724 2700 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 10364 30832 10428 30836
rect 10364 30776 10414 30832
rect 10414 30776 10428 30832
rect 10364 30772 10428 30776
rect 4660 30636 4724 30700
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 2452 30364 2516 30428
rect 5028 30364 5092 30428
rect 5396 30092 5460 30156
rect 10364 29956 10428 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 1900 29608 1964 29612
rect 1900 29552 1914 29608
rect 1914 29552 1964 29608
rect 1900 29548 1964 29552
rect 4660 29548 4724 29612
rect 11652 29276 11716 29340
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 5580 29004 5644 29068
rect 2452 28868 2516 28932
rect 10916 28868 10980 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 11468 28596 11532 28660
rect 8340 28324 8404 28388
rect 9628 28324 9692 28388
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 2636 28188 2700 28252
rect 8340 27916 8404 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 2084 27644 2148 27708
rect 7420 27644 7484 27708
rect 3924 27508 3988 27572
rect 7236 27508 7300 27572
rect 11468 27508 11532 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 7236 26828 7300 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 11284 26284 11348 26348
rect 8340 26148 8404 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 3740 25740 3804 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 9260 25332 9324 25396
rect 13492 25196 13556 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 15700 24924 15764 24988
rect 14596 24788 14660 24852
rect 4844 24652 4908 24716
rect 5580 24652 5644 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 5764 24108 5828 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 5212 23836 5276 23900
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 11652 23292 11716 23356
rect 11284 23156 11348 23220
rect 12572 23020 12636 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 5028 22748 5092 22812
rect 9628 22612 9692 22676
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 11652 22068 11716 22132
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 6132 21252 6196 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 10916 19408 10980 19412
rect 10916 19352 10966 19408
rect 10966 19352 10980 19408
rect 10916 19348 10980 19352
rect 13308 19212 13372 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 8524 18940 8588 19004
rect 11100 18804 11164 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 9812 17988 9876 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 3556 17716 3620 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 9444 16900 9508 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 3372 15948 3436 16012
rect 15148 15948 15212 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 13676 14512 13740 14516
rect 13676 14456 13726 14512
rect 13726 14456 13740 14512
rect 13676 14452 13740 14456
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 5396 13908 5460 13972
rect 15148 13696 15212 13700
rect 15148 13640 15198 13696
rect 15198 13640 15212 13696
rect 15148 13636 15212 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 7420 6156 7484 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 1900 5400 1964 5404
rect 1900 5344 1914 5400
rect 1914 5344 1964 5400
rect 1900 5340 1964 5344
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 5763 37092 5829 37093
rect 5763 37028 5764 37092
rect 5828 37028 5829 37092
rect 5763 37027 5829 37028
rect 8523 37092 8589 37093
rect 8523 37028 8524 37092
rect 8588 37028 8589 37092
rect 8523 37027 8589 37028
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 2083 36276 2149 36277
rect 2083 36212 2084 36276
rect 2148 36212 2149 36276
rect 2083 36211 2149 36212
rect 1899 29612 1965 29613
rect 1899 29548 1900 29612
rect 1964 29548 1965 29612
rect 1899 29547 1965 29548
rect 1902 5405 1962 29547
rect 2086 27709 2146 36211
rect 4208 35392 4528 36416
rect 5211 36140 5277 36141
rect 5211 36076 5212 36140
rect 5276 36076 5277 36140
rect 5211 36075 5277 36076
rect 4843 36004 4909 36005
rect 4843 35940 4844 36004
rect 4908 35940 4909 36004
rect 4843 35939 4909 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 3371 35052 3437 35053
rect 3371 34988 3372 35052
rect 3436 34988 3437 35052
rect 3371 34987 3437 34988
rect 2635 31788 2701 31789
rect 2635 31724 2636 31788
rect 2700 31724 2701 31788
rect 2635 31723 2701 31724
rect 2451 30428 2517 30429
rect 2451 30364 2452 30428
rect 2516 30364 2517 30428
rect 2451 30363 2517 30364
rect 2454 28933 2514 30363
rect 2451 28932 2517 28933
rect 2451 28868 2452 28932
rect 2516 28868 2517 28932
rect 2451 28867 2517 28868
rect 2638 28253 2698 31723
rect 2635 28252 2701 28253
rect 2635 28188 2636 28252
rect 2700 28188 2701 28252
rect 2635 28187 2701 28188
rect 2083 27708 2149 27709
rect 2083 27644 2084 27708
rect 2148 27644 2149 27708
rect 2083 27643 2149 27644
rect 3374 16013 3434 34987
rect 3555 34916 3621 34917
rect 3555 34852 3556 34916
rect 3620 34852 3621 34916
rect 3555 34851 3621 34852
rect 3558 17781 3618 34851
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 3923 34100 3989 34101
rect 3923 34036 3924 34100
rect 3988 34036 3989 34100
rect 3923 34035 3989 34036
rect 3739 31924 3805 31925
rect 3739 31860 3740 31924
rect 3804 31860 3805 31924
rect 3739 31859 3805 31860
rect 3742 25805 3802 31859
rect 3926 27573 3986 34035
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4659 30700 4725 30701
rect 4659 30636 4660 30700
rect 4724 30636 4725 30700
rect 4659 30635 4725 30636
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4662 29613 4722 30635
rect 4659 29612 4725 29613
rect 4659 29548 4660 29612
rect 4724 29548 4725 29612
rect 4659 29547 4725 29548
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 3923 27572 3989 27573
rect 3923 27508 3924 27572
rect 3988 27508 3989 27572
rect 3923 27507 3989 27508
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 3739 25804 3805 25805
rect 3739 25740 3740 25804
rect 3804 25740 3805 25804
rect 3739 25739 3805 25740
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4846 24717 4906 35939
rect 5027 30428 5093 30429
rect 5027 30364 5028 30428
rect 5092 30364 5093 30428
rect 5027 30363 5093 30364
rect 4843 24716 4909 24717
rect 4843 24652 4844 24716
rect 4908 24652 4909 24716
rect 4843 24651 4909 24652
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 5030 22813 5090 30363
rect 5214 23901 5274 36075
rect 5395 30156 5461 30157
rect 5395 30092 5396 30156
rect 5460 30092 5461 30156
rect 5395 30091 5461 30092
rect 5211 23900 5277 23901
rect 5211 23836 5212 23900
rect 5276 23836 5277 23900
rect 5211 23835 5277 23836
rect 5027 22812 5093 22813
rect 5027 22748 5028 22812
rect 5092 22748 5093 22812
rect 5027 22747 5093 22748
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 3555 17780 3621 17781
rect 3555 17716 3556 17780
rect 3620 17716 3621 17780
rect 3555 17715 3621 17716
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 3371 16012 3437 16013
rect 3371 15948 3372 16012
rect 3436 15948 3437 16012
rect 3371 15947 3437 15948
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 5398 13973 5458 30091
rect 5579 29068 5645 29069
rect 5579 29004 5580 29068
rect 5644 29004 5645 29068
rect 5579 29003 5645 29004
rect 5582 24717 5642 29003
rect 5579 24716 5645 24717
rect 5579 24652 5580 24716
rect 5644 24652 5645 24716
rect 5579 24651 5645 24652
rect 5766 24173 5826 37027
rect 8526 36549 8586 37027
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 8523 36548 8589 36549
rect 8523 36484 8524 36548
rect 8588 36484 8589 36548
rect 8523 36483 8589 36484
rect 13491 36548 13557 36549
rect 13491 36484 13492 36548
rect 13556 36484 13557 36548
rect 13491 36483 13557 36484
rect 7235 36004 7301 36005
rect 7235 35940 7236 36004
rect 7300 35940 7301 36004
rect 7235 35939 7301 35940
rect 6131 33420 6197 33421
rect 6131 33356 6132 33420
rect 6196 33356 6197 33420
rect 6131 33355 6197 33356
rect 5763 24172 5829 24173
rect 5763 24108 5764 24172
rect 5828 24108 5829 24172
rect 5763 24107 5829 24108
rect 6134 21317 6194 33355
rect 7238 27573 7298 35939
rect 8339 33148 8405 33149
rect 8339 33084 8340 33148
rect 8404 33084 8405 33148
rect 8339 33083 8405 33084
rect 8342 28389 8402 33083
rect 8339 28388 8405 28389
rect 8339 28324 8340 28388
rect 8404 28324 8405 28388
rect 8339 28323 8405 28324
rect 8339 27980 8405 27981
rect 8339 27916 8340 27980
rect 8404 27916 8405 27980
rect 8339 27915 8405 27916
rect 7419 27708 7485 27709
rect 7419 27644 7420 27708
rect 7484 27644 7485 27708
rect 7419 27643 7485 27644
rect 7235 27572 7301 27573
rect 7235 27508 7236 27572
rect 7300 27508 7301 27572
rect 7235 27507 7301 27508
rect 7238 26893 7298 27507
rect 7235 26892 7301 26893
rect 7235 26828 7236 26892
rect 7300 26828 7301 26892
rect 7235 26827 7301 26828
rect 6131 21316 6197 21317
rect 6131 21252 6132 21316
rect 6196 21252 6197 21316
rect 6131 21251 6197 21252
rect 5395 13972 5461 13973
rect 5395 13908 5396 13972
rect 5460 13908 5461 13972
rect 5395 13907 5461 13908
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 7422 6221 7482 27643
rect 8342 26213 8402 27915
rect 8339 26212 8405 26213
rect 8339 26148 8340 26212
rect 8404 26148 8405 26212
rect 8339 26147 8405 26148
rect 8526 19005 8586 36483
rect 11099 36140 11165 36141
rect 11099 36076 11100 36140
rect 11164 36076 11165 36140
rect 11099 36075 11165 36076
rect 9811 35460 9877 35461
rect 9811 35396 9812 35460
rect 9876 35396 9877 35460
rect 9811 35395 9877 35396
rect 9443 33012 9509 33013
rect 9443 32948 9444 33012
rect 9508 32948 9509 33012
rect 9443 32947 9509 32948
rect 9259 32332 9325 32333
rect 9259 32268 9260 32332
rect 9324 32268 9325 32332
rect 9259 32267 9325 32268
rect 9262 25397 9322 32267
rect 9259 25396 9325 25397
rect 9259 25332 9260 25396
rect 9324 25332 9325 25396
rect 9259 25331 9325 25332
rect 8523 19004 8589 19005
rect 8523 18940 8524 19004
rect 8588 18940 8589 19004
rect 8523 18939 8589 18940
rect 9446 16965 9506 32947
rect 9627 28388 9693 28389
rect 9627 28324 9628 28388
rect 9692 28324 9693 28388
rect 9627 28323 9693 28324
rect 9630 22677 9690 28323
rect 9627 22676 9693 22677
rect 9627 22612 9628 22676
rect 9692 22612 9693 22676
rect 9627 22611 9693 22612
rect 9814 18053 9874 35395
rect 11102 33557 11162 36075
rect 13307 34916 13373 34917
rect 13307 34852 13308 34916
rect 13372 34852 13373 34916
rect 13307 34851 13373 34852
rect 12571 34644 12637 34645
rect 12571 34580 12572 34644
rect 12636 34580 12637 34644
rect 12571 34579 12637 34580
rect 11099 33556 11165 33557
rect 11099 33492 11100 33556
rect 11164 33492 11165 33556
rect 11099 33491 11165 33492
rect 10363 30836 10429 30837
rect 10363 30772 10364 30836
rect 10428 30772 10429 30836
rect 10363 30771 10429 30772
rect 10366 30021 10426 30771
rect 10363 30020 10429 30021
rect 10363 29956 10364 30020
rect 10428 29956 10429 30020
rect 10363 29955 10429 29956
rect 10915 28932 10981 28933
rect 10915 28868 10916 28932
rect 10980 28868 10981 28932
rect 10915 28867 10981 28868
rect 10918 19413 10978 28867
rect 10915 19412 10981 19413
rect 10915 19348 10916 19412
rect 10980 19348 10981 19412
rect 10915 19347 10981 19348
rect 11102 18869 11162 33491
rect 11651 29340 11717 29341
rect 11651 29276 11652 29340
rect 11716 29276 11717 29340
rect 11651 29275 11717 29276
rect 11467 28660 11533 28661
rect 11467 28596 11468 28660
rect 11532 28596 11533 28660
rect 11467 28595 11533 28596
rect 11470 27573 11530 28595
rect 11467 27572 11533 27573
rect 11467 27508 11468 27572
rect 11532 27508 11533 27572
rect 11467 27507 11533 27508
rect 11283 26348 11349 26349
rect 11283 26284 11284 26348
rect 11348 26284 11349 26348
rect 11283 26283 11349 26284
rect 11286 23221 11346 26283
rect 11654 23357 11714 29275
rect 11651 23356 11717 23357
rect 11651 23292 11652 23356
rect 11716 23292 11717 23356
rect 11651 23291 11717 23292
rect 11283 23220 11349 23221
rect 11283 23156 11284 23220
rect 11348 23156 11349 23220
rect 11283 23155 11349 23156
rect 11654 22133 11714 23291
rect 12574 23085 12634 34579
rect 12571 23084 12637 23085
rect 12571 23020 12572 23084
rect 12636 23020 12637 23084
rect 12571 23019 12637 23020
rect 11651 22132 11717 22133
rect 11651 22068 11652 22132
rect 11716 22068 11717 22132
rect 11651 22067 11717 22068
rect 13310 19277 13370 34851
rect 13494 25261 13554 36483
rect 15699 36004 15765 36005
rect 15699 35940 15700 36004
rect 15764 35940 15765 36004
rect 15699 35939 15765 35940
rect 13675 35596 13741 35597
rect 13675 35532 13676 35596
rect 13740 35532 13741 35596
rect 13675 35531 13741 35532
rect 13491 25260 13557 25261
rect 13491 25196 13492 25260
rect 13556 25196 13557 25260
rect 13491 25195 13557 25196
rect 13307 19276 13373 19277
rect 13307 19212 13308 19276
rect 13372 19212 13373 19276
rect 13307 19211 13373 19212
rect 11099 18868 11165 18869
rect 11099 18804 11100 18868
rect 11164 18804 11165 18868
rect 11099 18803 11165 18804
rect 9811 18052 9877 18053
rect 9811 17988 9812 18052
rect 9876 17988 9877 18052
rect 9811 17987 9877 17988
rect 9443 16964 9509 16965
rect 9443 16900 9444 16964
rect 9508 16900 9509 16964
rect 9443 16899 9509 16900
rect 13678 14517 13738 35531
rect 14595 33148 14661 33149
rect 14595 33084 14596 33148
rect 14660 33084 14661 33148
rect 14595 33083 14661 33084
rect 14598 24853 14658 33083
rect 15702 24989 15762 35939
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 15699 24988 15765 24989
rect 15699 24924 15700 24988
rect 15764 24924 15765 24988
rect 15699 24923 15765 24924
rect 14595 24852 14661 24853
rect 14595 24788 14596 24852
rect 14660 24788 14661 24852
rect 14595 24787 14661 24788
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 15147 16012 15213 16013
rect 15147 15948 15148 16012
rect 15212 15948 15213 16012
rect 15147 15947 15213 15948
rect 13675 14516 13741 14517
rect 13675 14452 13676 14516
rect 13740 14452 13741 14516
rect 13675 14451 13741 14452
rect 15150 13701 15210 15947
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 15147 13700 15213 13701
rect 15147 13636 15148 13700
rect 15212 13636 15213 13700
rect 15147 13635 15213 13636
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 7419 6220 7485 6221
rect 7419 6156 7420 6220
rect 7484 6156 7485 6220
rect 7419 6155 7485 6156
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 1899 5404 1965 5405
rect 1899 5340 1900 5404
rect 1964 5340 1965 5404
rect 1899 5339 1965 5340
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17940 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 14352 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 19872 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1667941163
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1667941163
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1667941163
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1667941163
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1667941163
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1667941163
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1667941163
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_20
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_24
timestamp 1667941163
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1667941163
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1667941163
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1667941163
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_396
timestamp 1667941163
transform 1 0 37536 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_21
timestamp 1667941163
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_25
timestamp 1667941163
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_37
timestamp 1667941163
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1667941163
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_329
timestamp 1667941163
transform 1 0 31372 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1667941163
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_118
timestamp 1667941163
transform 1 0 11960 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_130
timestamp 1667941163
transform 1 0 13064 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_142
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_150
timestamp 1667941163
transform 1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1667941163
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_182
timestamp 1667941163
transform 1 0 17848 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_194
timestamp 1667941163
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_209
timestamp 1667941163
transform 1 0 20332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1667941163
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_292
timestamp 1667941163
transform 1 0 27968 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_304
timestamp 1667941163
transform 1 0 29072 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_316
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1667941163
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_42
timestamp 1667941163
transform 1 0 4968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_54
timestamp 1667941163
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_60
timestamp 1667941163
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_72
timestamp 1667941163
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_94
timestamp 1667941163
transform 1 0 9752 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_106
timestamp 1667941163
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_118
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1667941163
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1667941163
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_215
timestamp 1667941163
transform 1 0 20884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_219
timestamp 1667941163
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_231
timestamp 1667941163
transform 1 0 22356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1667941163
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_258
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_270
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1667941163
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_317
timestamp 1667941163
transform 1 0 30268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_341
timestamp 1667941163
transform 1 0 32476 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_346
timestamp 1667941163
transform 1 0 32936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1667941163
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_392
timestamp 1667941163
transform 1 0 37168 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_404
timestamp 1667941163
transform 1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1667941163
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1667941163
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1667941163
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_85
timestamp 1667941163
transform 1 0 8924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_97
timestamp 1667941163
transform 1 0 10028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1667941163
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_118
timestamp 1667941163
transform 1 0 11960 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_130
timestamp 1667941163
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_142
timestamp 1667941163
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_154
timestamp 1667941163
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_304
timestamp 1667941163
transform 1 0 29072 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_316
timestamp 1667941163
transform 1 0 30176 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1667941163
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_259
timestamp 1667941163
transform 1 0 24932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_271
timestamp 1667941163
transform 1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_283
timestamp 1667941163
transform 1 0 27140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_295
timestamp 1667941163
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_357
timestamp 1667941163
transform 1 0 33948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_363
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1667941163
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1667941163
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1667941163
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1667941163
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_90
timestamp 1667941163
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_102
timestamp 1667941163
transform 1 0 10488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_114
timestamp 1667941163
transform 1 0 11592 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1667941163
transform 1 0 12696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1667941163
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_283
timestamp 1667941163
transform 1 0 27140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_295
timestamp 1667941163
transform 1 0 28244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_374
timestamp 1667941163
transform 1 0 35512 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_386
timestamp 1667941163
transform 1 0 36616 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_398
timestamp 1667941163
transform 1 0 37720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1667941163
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_94
timestamp 1667941163
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1667941163
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_118
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_130
timestamp 1667941163
transform 1 0 13064 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_142
timestamp 1667941163
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1667941163
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_200
timestamp 1667941163
transform 1 0 19504 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_212
timestamp 1667941163
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_233
timestamp 1667941163
transform 1 0 22540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_245
timestamp 1667941163
transform 1 0 23644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_257
timestamp 1667941163
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1667941163
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1667941163
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1667941163
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_188
timestamp 1667941163
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1667941163
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1667941163
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_46
timestamp 1667941163
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_70
timestamp 1667941163
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_103
timestamp 1667941163
transform 1 0 10580 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_107
timestamp 1667941163
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_119
timestamp 1667941163
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_118
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_130
timestamp 1667941163
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_142
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_154
timestamp 1667941163
transform 1 0 15272 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1667941163
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_188
timestamp 1667941163
transform 1 0 18400 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_200
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_247
timestamp 1667941163
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_259
timestamp 1667941163
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_271
timestamp 1667941163
transform 1 0 26036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1667941163
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_214
timestamp 1667941163
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_226
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_238
timestamp 1667941163
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_342
timestamp 1667941163
transform 1 0 32568 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_354
timestamp 1667941163
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_366
timestamp 1667941163
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_378
timestamp 1667941163
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_60
timestamp 1667941163
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_72
timestamp 1667941163
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1667941163
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_354
timestamp 1667941163
transform 1 0 33672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1667941163
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1667941163
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1667941163
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1667941163
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1667941163
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp 1667941163
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1667941163
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1667941163
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_248
timestamp 1667941163
transform 1 0 23920 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_260
timestamp 1667941163
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1667941163
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_369
timestamp 1667941163
transform 1 0 35052 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_375
timestamp 1667941163
transform 1 0 35604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1667941163
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1667941163
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_161
timestamp 1667941163
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_145
timestamp 1667941163
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1667941163
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_176
timestamp 1667941163
transform 1 0 17296 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_200
timestamp 1667941163
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_212
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1667941163
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1667941163
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1667941163
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1667941163
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_167
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_185
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1667941163
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_370
timestamp 1667941163
transform 1 0 35144 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_382
timestamp 1667941163
transform 1 0 36248 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_394
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_400
timestamp 1667941163
transform 1 0 37904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1667941163
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1667941163
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_85
timestamp 1667941163
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1667941163
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1667941163
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1667941163
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_191
timestamp 1667941163
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_203
timestamp 1667941163
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_95
timestamp 1667941163
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_104
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1667941163
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1667941163
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_160
timestamp 1667941163
transform 1 0 15824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1667941163
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_202
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_214
timestamp 1667941163
transform 1 0 20792 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_226
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_238
timestamp 1667941163
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_370
timestamp 1667941163
transform 1 0 35144 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_382
timestamp 1667941163
transform 1 0 36248 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_394
timestamp 1667941163
transform 1 0 37352 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1667941163
transform 1 0 38456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1667941163
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_94
timestamp 1667941163
transform 1 0 9752 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1667941163
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1667941163
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_136
timestamp 1667941163
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1667941163
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_174
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_354
timestamp 1667941163
transform 1 0 33672 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_366
timestamp 1667941163
transform 1 0 34776 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_378
timestamp 1667941163
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1667941163
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_92
timestamp 1667941163
transform 1 0 9568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1667941163
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1667941163
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_118
timestamp 1667941163
transform 1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_126
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_168
timestamp 1667941163
transform 1 0 16560 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1667941163
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1667941163
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1667941163
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1667941163
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_216
timestamp 1667941163
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_240
timestamp 1667941163
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1667941163
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 1667941163
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1667941163
transform 1 0 8188 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_86
timestamp 1667941163
transform 1 0 9016 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1667941163
transform 1 0 9568 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1667941163
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1667941163
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1667941163
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1667941163
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_156
timestamp 1667941163
transform 1 0 15456 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_162
timestamp 1667941163
transform 1 0 16008 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1667941163
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1667941163
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_230
timestamp 1667941163
transform 1 0 22264 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_242
timestamp 1667941163
transform 1 0 23368 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_254
timestamp 1667941163
transform 1 0 24472 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_266
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_71
timestamp 1667941163
transform 1 0 7636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1667941163
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_156
timestamp 1667941163
transform 1 0 15456 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_183
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1667941163
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_223
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1667941163
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1667941163
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1667941163
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1667941163
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_70
timestamp 1667941163
transform 1 0 7544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_77
timestamp 1667941163
transform 1 0 8188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_84
timestamp 1667941163
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1667941163
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1667941163
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_124
timestamp 1667941163
transform 1 0 12512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_136
timestamp 1667941163
transform 1 0 13616 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1667941163
transform 1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1667941163
transform 1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_252
timestamp 1667941163
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_264
timestamp 1667941163
transform 1 0 25392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1667941163
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1667941163
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_98
timestamp 1667941163
transform 1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1667941163
transform 1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1667941163
transform 1 0 12328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_126
timestamp 1667941163
transform 1 0 12696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_156
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_214
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1667941163
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1667941163
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1667941163
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_314
timestamp 1667941163
transform 1 0 29992 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_326
timestamp 1667941163
transform 1 0 31096 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_338
timestamp 1667941163
transform 1 0 32200 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_350
timestamp 1667941163
transform 1 0 33304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1667941163
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_370
timestamp 1667941163
transform 1 0 35144 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_382
timestamp 1667941163
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1667941163
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1667941163
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_8
timestamp 1667941163
transform 1 0 1840 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_20
timestamp 1667941163
transform 1 0 2944 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_32
timestamp 1667941163
transform 1 0 4048 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1667941163
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1667941163
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1667941163
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_89
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_126
timestamp 1667941163
transform 1 0 12696 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_134
timestamp 1667941163
transform 1 0 13432 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1667941163
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_155
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_180
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_203
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1667941163
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_250
timestamp 1667941163
transform 1 0 24104 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_262
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1667941163
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_304
timestamp 1667941163
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1667941163
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_49
timestamp 1667941163
transform 1 0 5612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1667941163
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1667941163
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1667941163
transform 1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1667941163
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_110
timestamp 1667941163
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_118
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1667941163
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1667941163
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_171
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_183
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1667941163
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1667941163
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1667941163
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1667941163
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_282
timestamp 1667941163
transform 1 0 27048 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_294
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1667941163
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1667941163
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1667941163
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1667941163
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1667941163
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1667941163
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_124
timestamp 1667941163
transform 1 0 12512 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_130
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1667941163
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1667941163
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1667941163
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_201
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1667941163
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_256
timestamp 1667941163
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_263
timestamp 1667941163
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1667941163
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_57
timestamp 1667941163
transform 1 0 6348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_61
timestamp 1667941163
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_68
timestamp 1667941163
transform 1 0 7360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_94
timestamp 1667941163
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_106
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_114
timestamp 1667941163
transform 1 0 11592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_146
timestamp 1667941163
transform 1 0 14536 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_172
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1667941163
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1667941163
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_207
timestamp 1667941163
transform 1 0 20148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1667941163
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_223
timestamp 1667941163
transform 1 0 21620 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_240
timestamp 1667941163
transform 1 0 23184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1667941163
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_258
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_270
timestamp 1667941163
transform 1 0 25944 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_282
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_294
timestamp 1667941163
transform 1 0 28152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1667941163
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1667941163
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_94
timestamp 1667941163
transform 1 0 9752 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_123
timestamp 1667941163
transform 1 0 12420 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_143
timestamp 1667941163
transform 1 0 14260 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1667941163
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_235
timestamp 1667941163
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_59
timestamp 1667941163
transform 1 0 6532 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1667941163
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1667941163
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_95
timestamp 1667941163
transform 1 0 9844 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_103
timestamp 1667941163
transform 1 0 10580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_114
timestamp 1667941163
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1667941163
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1667941163
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_178
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_207
timestamp 1667941163
transform 1 0 20148 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1667941163
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_228
timestamp 1667941163
transform 1 0 22080 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_236
timestamp 1667941163
transform 1 0 22816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1667941163
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_330
timestamp 1667941163
transform 1 0 31464 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_342
timestamp 1667941163
transform 1 0 32568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1667941163
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1667941163
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp 1667941163
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_82
timestamp 1667941163
transform 1 0 8648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_89
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_96
timestamp 1667941163
transform 1 0 9936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_103
timestamp 1667941163
transform 1 0 10580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1667941163
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1667941163
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_133
timestamp 1667941163
transform 1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_140
timestamp 1667941163
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_159
timestamp 1667941163
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_176
timestamp 1667941163
transform 1 0 17296 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_183
timestamp 1667941163
transform 1 0 17940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1667941163
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_209
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1667941163
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1667941163
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1667941163
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_320
timestamp 1667941163
transform 1 0 30544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1667941163
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 1667941163
transform 1 0 34684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_369
timestamp 1667941163
transform 1 0 35052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1667941163
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1667941163
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_8
timestamp 1667941163
transform 1 0 1840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1667941163
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1667941163
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_98
timestamp 1667941163
transform 1 0 10120 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_114
timestamp 1667941163
transform 1 0 11592 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1667941163
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_156
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_167
timestamp 1667941163
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_180
timestamp 1667941163
transform 1 0 17664 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_224
timestamp 1667941163
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1667941163
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_258
timestamp 1667941163
transform 1 0 24840 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_270
timestamp 1667941163
transform 1 0 25944 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_282
timestamp 1667941163
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_294
timestamp 1667941163
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1667941163
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_8
timestamp 1667941163
transform 1 0 1840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_22
timestamp 1667941163
transform 1 0 3128 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1667941163
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1667941163
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_64
timestamp 1667941163
transform 1 0 6992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_72
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_77
timestamp 1667941163
transform 1 0 8188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1667941163
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_97
timestamp 1667941163
transform 1 0 10028 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_123
timestamp 1667941163
transform 1 0 12420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_131
timestamp 1667941163
transform 1 0 13156 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_143
timestamp 1667941163
transform 1 0 14260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1667941163
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1667941163
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1667941163
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_201
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_215
timestamp 1667941163
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_263
timestamp 1667941163
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_16
timestamp 1667941163
transform 1 0 2576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1667941163
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 1667941163
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_64
timestamp 1667941163
transform 1 0 6992 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_73
timestamp 1667941163
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1667941163
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1667941163
transform 1 0 9476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_100
timestamp 1667941163
transform 1 0 10304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_115
timestamp 1667941163
transform 1 0 11684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1667941163
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_131
timestamp 1667941163
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1667941163
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1667941163
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_169
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1667941163
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_212
timestamp 1667941163
transform 1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_219
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_236
timestamp 1667941163
transform 1 0 22816 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_270
timestamp 1667941163
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1667941163
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_14
timestamp 1667941163
transform 1 0 2392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_35
timestamp 1667941163
transform 1 0 4324 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_44
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_62
timestamp 1667941163
transform 1 0 6808 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 7544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_74
timestamp 1667941163
transform 1 0 7912 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_82
timestamp 1667941163
transform 1 0 8648 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_86
timestamp 1667941163
transform 1 0 9016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_99
timestamp 1667941163
transform 1 0 10212 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1667941163
transform 1 0 10580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_122
timestamp 1667941163
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_129
timestamp 1667941163
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_136
timestamp 1667941163
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1667941163
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_175
timestamp 1667941163
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_188
timestamp 1667941163
transform 1 0 18400 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1667941163
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_212
timestamp 1667941163
transform 1 0 20608 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1667941163
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_229
timestamp 1667941163
transform 1 0 22172 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_233
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_248
timestamp 1667941163
transform 1 0 23920 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_255
timestamp 1667941163
transform 1 0 24564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1667941163
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1667941163
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1667941163
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_290
timestamp 1667941163
transform 1 0 27784 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_302
timestamp 1667941163
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_314
timestamp 1667941163
transform 1 0 29992 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_326
timestamp 1667941163
transform 1 0 31096 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1667941163
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1667941163
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_34
timestamp 1667941163
transform 1 0 4232 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_40
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_44
timestamp 1667941163
transform 1 0 5152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_52
timestamp 1667941163
transform 1 0 5888 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1667941163
transform 1 0 6624 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1667941163
transform 1 0 6992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_71
timestamp 1667941163
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1667941163
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_92
timestamp 1667941163
transform 1 0 9568 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_101
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_111
timestamp 1667941163
transform 1 0 11316 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_118
timestamp 1667941163
transform 1 0 11960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1667941163
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_152
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_160
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_169
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1667941163
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_185
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_216
timestamp 1667941163
transform 1 0 20976 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_222
timestamp 1667941163
transform 1 0 21528 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_231
timestamp 1667941163
transform 1 0 22356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_235
timestamp 1667941163
transform 1 0 22724 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1667941163
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_258
timestamp 1667941163
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_270
timestamp 1667941163
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_282
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_28
timestamp 1667941163
transform 1 0 3680 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_73
timestamp 1667941163
transform 1 0 7820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_97
timestamp 1667941163
transform 1 0 10028 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1667941163
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_132
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_142
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1667941163
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1667941163
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_209
timestamp 1667941163
transform 1 0 20332 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_242
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1667941163
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_263
timestamp 1667941163
transform 1 0 25300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1667941163
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_285
timestamp 1667941163
transform 1 0 27324 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_289
timestamp 1667941163
transform 1 0 27692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_301
timestamp 1667941163
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_313
timestamp 1667941163
transform 1 0 29900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_325
timestamp 1667941163
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1667941163
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_365
timestamp 1667941163
transform 1 0 34684 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_377
timestamp 1667941163
transform 1 0 35788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1667941163
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1667941163
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_51
timestamp 1667941163
transform 1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1667941163
transform 1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1667941163
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_99
timestamp 1667941163
transform 1 0 10212 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_110
timestamp 1667941163
transform 1 0 11224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_124
timestamp 1667941163
transform 1 0 12512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1667941163
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_161
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_173
timestamp 1667941163
transform 1 0 17020 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1667941163
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_208
timestamp 1667941163
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1667941163
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_229
timestamp 1667941163
transform 1 0 22172 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_236
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1667941163
transform 1 0 24840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_272
timestamp 1667941163
transform 1 0 26128 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_284
timestamp 1667941163
transform 1 0 27232 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_296
timestamp 1667941163
transform 1 0 28336 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_370
timestamp 1667941163
transform 1 0 35144 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_382
timestamp 1667941163
transform 1 0 36248 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_394
timestamp 1667941163
transform 1 0 37352 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1667941163
transform 1 0 38456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_20
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1667941163
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1667941163
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1667941163
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1667941163
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_150
timestamp 1667941163
transform 1 0 14904 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1667941163
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_192
timestamp 1667941163
transform 1 0 18768 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_200
timestamp 1667941163
transform 1 0 19504 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_204
timestamp 1667941163
transform 1 0 19872 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1667941163
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_247
timestamp 1667941163
transform 1 0 23828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_253
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_262
timestamp 1667941163
transform 1 0 25208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1667941163
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_301
timestamp 1667941163
transform 1 0 28796 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_307
timestamp 1667941163
transform 1 0 29348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_319
timestamp 1667941163
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1667941163
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_344
timestamp 1667941163
transform 1 0 32752 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_356
timestamp 1667941163
transform 1 0 33856 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_368
timestamp 1667941163
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_380
timestamp 1667941163
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_40
timestamp 1667941163
transform 1 0 4784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_67
timestamp 1667941163
transform 1 0 7268 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_73
timestamp 1667941163
transform 1 0 7820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1667941163
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1667941163
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1667941163
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_159
timestamp 1667941163
transform 1 0 15732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_171
timestamp 1667941163
transform 1 0 16836 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_182
timestamp 1667941163
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1667941163
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_227
timestamp 1667941163
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_239
timestamp 1667941163
transform 1 0 23092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1667941163
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_270
timestamp 1667941163
transform 1 0 25944 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_282
timestamp 1667941163
transform 1 0 27048 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_294
timestamp 1667941163
transform 1 0 28152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1667941163
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_329
timestamp 1667941163
transform 1 0 31372 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_335
timestamp 1667941163
transform 1 0 31924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_347
timestamp 1667941163
transform 1 0 33028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1667941163
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_28
timestamp 1667941163
transform 1 0 3680 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1667941163
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_63
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_87
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_103
timestamp 1667941163
transform 1 0 10580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1667941163
transform 1 0 13524 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_143
timestamp 1667941163
transform 1 0 14260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_147
timestamp 1667941163
transform 1 0 14628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_154
timestamp 1667941163
transform 1 0 15272 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_183
timestamp 1667941163
transform 1 0 17940 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_192
timestamp 1667941163
transform 1 0 18768 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1667941163
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1667941163
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1667941163
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_242
timestamp 1667941163
transform 1 0 23368 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1667941163
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_36
timestamp 1667941163
transform 1 0 4416 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_48
timestamp 1667941163
transform 1 0 5520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_72
timestamp 1667941163
transform 1 0 7728 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_78
timestamp 1667941163
transform 1 0 8280 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1667941163
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1667941163
transform 1 0 9660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_120
timestamp 1667941163
transform 1 0 12144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1667941163
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_147
timestamp 1667941163
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_151
timestamp 1667941163
transform 1 0 14996 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_162
timestamp 1667941163
transform 1 0 16008 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_168
timestamp 1667941163
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_172
timestamp 1667941163
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1667941163
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_186
timestamp 1667941163
transform 1 0 18216 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1667941163
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1667941163
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1667941163
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_227
timestamp 1667941163
transform 1 0 21988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1667941163
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_38
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_42
timestamp 1667941163
transform 1 0 4968 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1667941163
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_97
timestamp 1667941163
transform 1 0 10028 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1667941163
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_152
timestamp 1667941163
transform 1 0 15088 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1667941163
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_180
timestamp 1667941163
transform 1 0 17664 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 1667941163
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_196
timestamp 1667941163
transform 1 0 19136 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_204
timestamp 1667941163
transform 1 0 19872 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_213
timestamp 1667941163
transform 1 0 20700 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_234
timestamp 1667941163
transform 1 0 22632 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1667941163
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_245
timestamp 1667941163
transform 1 0 23644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_257
timestamp 1667941163
transform 1 0 24748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_265
timestamp 1667941163
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1667941163
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 1667941163
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_14
timestamp 1667941163
transform 1 0 2392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1667941163
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_34
timestamp 1667941163
transform 1 0 4232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_61
timestamp 1667941163
transform 1 0 6716 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1667941163
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_108
timestamp 1667941163
transform 1 0 11040 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_120
timestamp 1667941163
transform 1 0 12144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_124
timestamp 1667941163
transform 1 0 12512 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_128
timestamp 1667941163
transform 1 0 12880 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_134
timestamp 1667941163
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_148
timestamp 1667941163
transform 1 0 14720 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_155
timestamp 1667941163
transform 1 0 15364 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_167
timestamp 1667941163
transform 1 0 16468 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_173
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_182
timestamp 1667941163
transform 1 0 17848 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_190
timestamp 1667941163
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_204
timestamp 1667941163
transform 1 0 19872 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_211
timestamp 1667941163
transform 1 0 20516 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1667941163
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_225
timestamp 1667941163
transform 1 0 21804 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_237
timestamp 1667941163
transform 1 0 22908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_258
timestamp 1667941163
transform 1 0 24840 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_270
timestamp 1667941163
transform 1 0 25944 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_282
timestamp 1667941163
transform 1 0 27048 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_294
timestamp 1667941163
transform 1 0 28152 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1667941163
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_7
timestamp 1667941163
transform 1 0 1748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_31
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_38
timestamp 1667941163
transform 1 0 4600 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_45
timestamp 1667941163
transform 1 0 5244 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_80
timestamp 1667941163
transform 1 0 8464 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_104
timestamp 1667941163
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_118
timestamp 1667941163
transform 1 0 11960 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_126
timestamp 1667941163
transform 1 0 12696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_130
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_142
timestamp 1667941163
transform 1 0 14168 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_146
timestamp 1667941163
transform 1 0 14536 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_151
timestamp 1667941163
transform 1 0 14996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_155
timestamp 1667941163
transform 1 0 15364 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1667941163
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_177
timestamp 1667941163
transform 1 0 17388 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_182
timestamp 1667941163
transform 1 0 17848 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_210
timestamp 1667941163
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1667941163
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_259
timestamp 1667941163
transform 1 0 24932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_263
timestamp 1667941163
transform 1 0 25300 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_296
timestamp 1667941163
transform 1 0 28336 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_308
timestamp 1667941163
transform 1 0 29440 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_320
timestamp 1667941163
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1667941163
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_357
timestamp 1667941163
transform 1 0 33948 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_363
timestamp 1667941163
transform 1 0 34500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_375
timestamp 1667941163
transform 1 0 35604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_387
timestamp 1667941163
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1667941163
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_14
timestamp 1667941163
transform 1 0 2392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_34
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_49
timestamp 1667941163
transform 1 0 5612 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_54
timestamp 1667941163
transform 1 0 6072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_61
timestamp 1667941163
transform 1 0 6716 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_68
timestamp 1667941163
transform 1 0 7360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_75
timestamp 1667941163
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1667941163
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_104
timestamp 1667941163
transform 1 0 10672 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_111
timestamp 1667941163
transform 1 0 11316 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_120
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_127
timestamp 1667941163
transform 1 0 12788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1667941163
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_160
timestamp 1667941163
transform 1 0 15824 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_164
timestamp 1667941163
transform 1 0 16192 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_168
timestamp 1667941163
transform 1 0 16560 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1667941163
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_184
timestamp 1667941163
transform 1 0 18032 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_202
timestamp 1667941163
transform 1 0 19688 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_214
timestamp 1667941163
transform 1 0 20792 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_226
timestamp 1667941163
transform 1 0 21896 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_238
timestamp 1667941163
transform 1 0 23000 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1667941163
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_280
timestamp 1667941163
transform 1 0 26864 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_287
timestamp 1667941163
transform 1 0 27508 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1667941163
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_13
timestamp 1667941163
transform 1 0 2300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_38
timestamp 1667941163
transform 1 0 4600 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_45
timestamp 1667941163
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1667941163
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_79
timestamp 1667941163
transform 1 0 8372 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_119
timestamp 1667941163
transform 1 0 12052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_123
timestamp 1667941163
transform 1 0 12420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_130
timestamp 1667941163
transform 1 0 13064 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_144
timestamp 1667941163
transform 1 0 14352 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_151
timestamp 1667941163
transform 1 0 14996 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_158
timestamp 1667941163
transform 1 0 15640 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1667941163
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_174
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_182
timestamp 1667941163
transform 1 0 17848 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1667941163
transform 1 0 18308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_200
timestamp 1667941163
transform 1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1667941163
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_257
timestamp 1667941163
transform 1 0 24748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_342
timestamp 1667941163
transform 1 0 32568 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_354
timestamp 1667941163
transform 1 0 33672 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_366
timestamp 1667941163
transform 1 0 34776 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_378
timestamp 1667941163
transform 1 0 35880 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1667941163
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1667941163
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_40
timestamp 1667941163
transform 1 0 4784 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_64
timestamp 1667941163
transform 1 0 6992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_71
timestamp 1667941163
transform 1 0 7636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1667941163
transform 1 0 9476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_95
timestamp 1667941163
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_102
timestamp 1667941163
transform 1 0 10488 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_110
timestamp 1667941163
transform 1 0 11224 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_131
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1667941163
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_160
timestamp 1667941163
transform 1 0 15824 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1667941163
transform 1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_174
timestamp 1667941163
transform 1 0 17112 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_186
timestamp 1667941163
transform 1 0 18216 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_190
timestamp 1667941163
transform 1 0 18584 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_203
timestamp 1667941163
transform 1 0 19780 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_216
timestamp 1667941163
transform 1 0 20976 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_224
timestamp 1667941163
transform 1 0 21712 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_235
timestamp 1667941163
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1667941163
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_264
timestamp 1667941163
transform 1 0 25392 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_271
timestamp 1667941163
transform 1 0 26036 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_283
timestamp 1667941163
transform 1 0 27140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_295
timestamp 1667941163
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_13
timestamp 1667941163
transform 1 0 2300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_38
timestamp 1667941163
transform 1 0 4600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1667941163
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_62
timestamp 1667941163
transform 1 0 6808 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_70
timestamp 1667941163
transform 1 0 7544 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_95
timestamp 1667941163
transform 1 0 9844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_102
timestamp 1667941163
transform 1 0 10488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1667941163
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_135
timestamp 1667941163
transform 1 0 13524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_142
timestamp 1667941163
transform 1 0 14168 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_156
timestamp 1667941163
transform 1 0 15456 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1667941163
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_174
timestamp 1667941163
transform 1 0 17112 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_189
timestamp 1667941163
transform 1 0 18492 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_194
timestamp 1667941163
transform 1 0 18952 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_203
timestamp 1667941163
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_215
timestamp 1667941163
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_239
timestamp 1667941163
transform 1 0 23092 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_247
timestamp 1667941163
transform 1 0 23828 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_251
timestamp 1667941163
transform 1 0 24196 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_263
timestamp 1667941163
transform 1 0 25300 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1667941163
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_300
timestamp 1667941163
transform 1 0 28704 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_312
timestamp 1667941163
transform 1 0 29808 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_324
timestamp 1667941163
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_342
timestamp 1667941163
transform 1 0 32568 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_350
timestamp 1667941163
transform 1 0 33304 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_356
timestamp 1667941163
transform 1 0 33856 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_363
timestamp 1667941163
transform 1 0 34500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_375
timestamp 1667941163
transform 1 0 35604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1667941163
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_401
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_16
timestamp 1667941163
transform 1 0 2576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1667941163
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_34
timestamp 1667941163
transform 1 0 4232 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_48
timestamp 1667941163
transform 1 0 5520 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_55
timestamp 1667941163
transform 1 0 6164 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_90
timestamp 1667941163
transform 1 0 9384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_104
timestamp 1667941163
transform 1 0 10672 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_130
timestamp 1667941163
transform 1 0 13064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1667941163
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1667941163
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_154
timestamp 1667941163
transform 1 0 15272 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_162
timestamp 1667941163
transform 1 0 16008 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1667941163
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1667941163
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_181
timestamp 1667941163
transform 1 0 17756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 1667941163
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_217
timestamp 1667941163
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1667941163
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_230
timestamp 1667941163
transform 1 0 22264 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_237
timestamp 1667941163
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1667941163
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_260
timestamp 1667941163
transform 1 0 25024 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_272
timestamp 1667941163
transform 1 0 26128 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_284
timestamp 1667941163
transform 1 0 27232 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_296
timestamp 1667941163
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1667941163
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1667941163
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1667941163
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_30
timestamp 1667941163
transform 1 0 3864 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1667941163
transform 1 0 6808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_96
timestamp 1667941163
transform 1 0 9936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_103
timestamp 1667941163
transform 1 0 10580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1667941163
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_135
timestamp 1667941163
transform 1 0 13524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_142
timestamp 1667941163
transform 1 0 14168 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_156
timestamp 1667941163
transform 1 0 15456 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_174
timestamp 1667941163
transform 1 0 17112 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_189
timestamp 1667941163
transform 1 0 18492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_201
timestamp 1667941163
transform 1 0 19596 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_210
timestamp 1667941163
transform 1 0 20424 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1667941163
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1667941163
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_7
timestamp 1667941163
transform 1 0 1748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_14
timestamp 1667941163
transform 1 0 2392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1667941163
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_54
timestamp 1667941163
transform 1 0 6072 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_107
timestamp 1667941163
transform 1 0 10948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1667941163
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_152
timestamp 1667941163
transform 1 0 15088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_159
timestamp 1667941163
transform 1 0 15732 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_172
timestamp 1667941163
transform 1 0 16928 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_179
timestamp 1667941163
transform 1 0 17572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_186
timestamp 1667941163
transform 1 0 18216 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1667941163
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_381
timestamp 1667941163
transform 1 0 36156 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_393
timestamp 1667941163
transform 1 0 37260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1667941163
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_7
timestamp 1667941163
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_14
timestamp 1667941163
transform 1 0 2392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_24
timestamp 1667941163
transform 1 0 3312 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_32
timestamp 1667941163
transform 1 0 4048 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1667941163
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_63
timestamp 1667941163
transform 1 0 6900 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_71
timestamp 1667941163
transform 1 0 7636 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_94
timestamp 1667941163
transform 1 0 9752 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_101
timestamp 1667941163
transform 1 0 10396 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1667941163
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_136
timestamp 1667941163
transform 1 0 13616 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_144
timestamp 1667941163
transform 1 0 14352 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_151
timestamp 1667941163
transform 1 0 14996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_158
timestamp 1667941163
transform 1 0 15640 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_174
timestamp 1667941163
transform 1 0 17112 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_188
timestamp 1667941163
transform 1 0 18400 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_200
timestamp 1667941163
transform 1 0 19504 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_212
timestamp 1667941163
transform 1 0 20608 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1667941163
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_35
timestamp 1667941163
transform 1 0 4324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_56
timestamp 1667941163
transform 1 0 6256 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_81
timestamp 1667941163
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_108
timestamp 1667941163
transform 1 0 11040 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_112
timestamp 1667941163
transform 1 0 11408 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_134
timestamp 1667941163
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_163
timestamp 1667941163
transform 1 0 16100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_170
timestamp 1667941163
transform 1 0 16744 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_176
timestamp 1667941163
transform 1 0 17296 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_180
timestamp 1667941163
transform 1 0 17664 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1667941163
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_238
timestamp 1667941163
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1667941163
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1667941163
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_14
timestamp 1667941163
transform 1 0 2392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_20
timestamp 1667941163
transform 1 0 2944 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_42
timestamp 1667941163
transform 1 0 4968 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_61
timestamp 1667941163
transform 1 0 6716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_83
timestamp 1667941163
transform 1 0 8740 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1667941163
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_142
timestamp 1667941163
transform 1 0 14168 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_156
timestamp 1667941163
transform 1 0 15456 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1667941163
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_35
timestamp 1667941163
transform 1 0 4324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_57
timestamp 1667941163
transform 1 0 6348 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_91
timestamp 1667941163
transform 1 0 9476 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_95
timestamp 1667941163
transform 1 0 9844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_100
timestamp 1667941163
transform 1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_125
timestamp 1667941163
transform 1 0 12604 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1667941163
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_148
timestamp 1667941163
transform 1 0 14720 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1667941163
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_162
timestamp 1667941163
transform 1 0 16008 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_169
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_176
timestamp 1667941163
transform 1 0 17296 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_181
timestamp 1667941163
transform 1 0 17756 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_185
timestamp 1667941163
transform 1 0 18124 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1667941163
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_28
timestamp 1667941163
transform 1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_32
timestamp 1667941163
transform 1 0 4048 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_63
timestamp 1667941163
transform 1 0 6900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1667941163
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1667941163
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1667941163
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_188
timestamp 1667941163
transform 1 0 18400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_195
timestamp 1667941163
transform 1 0 19044 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_202
timestamp 1667941163
transform 1 0 19688 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1667941163
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_398
timestamp 1667941163
transform 1 0 37720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1667941163
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_135
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1667941163
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1667941163
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1667941163
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_386
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0410_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 24748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 24656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 17296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 22632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 21344 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 21988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 16008 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 15456 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 19504 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 23092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 13892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 14352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 21712 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 24380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 19504 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 18032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 15272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 10396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 13524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 15640 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 14352 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 15088 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 19596 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 12420 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 5704 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 4876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 7176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 9384 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 14536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 8372 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 18584 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 18676 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 18676 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 11868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 7268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 9568 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 25024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 7268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 7728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 4140 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 6716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 10212 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 19596 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 15548 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 18216 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0532_
timestamp 1667941163
transform 1 0 9844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 21804 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 26312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0541_
timestamp 1667941163
transform 1 0 25576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 20976 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 17296 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 25024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 16652 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 23736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 14904 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1667941163
transform 1 0 14536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 15548 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 21528 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 22724 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 23460 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 25668 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 20700 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 23736 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 12604 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1667941163
transform 1 0 12788 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 18124 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 24932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1667941163
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1667941163
transform 1 0 24288 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 18216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 16192 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 12144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1667941163
transform 1 0 13524 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 6440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1667941163
transform 1 0 13064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1667941163
transform 1 0 9292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1667941163
transform 1 0 14444 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 15824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 20240 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 18952 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 11316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 11684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 10304 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1667941163
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1667941163
transform 1 0 10672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 8372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 8372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 10304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1667941163
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 13524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1667941163
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 12696 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 14720 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 17940 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1667941163
transform 1 0 18584 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 14996 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 20056 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 17480 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 9292 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1667941163
transform 1 0 12880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 11040 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 14904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 16008 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1667941163
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0677_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 13984 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 7728 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 12880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform 1 0 12880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 7360 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1667941163
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1667941163
transform 1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform 1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 13432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 5520 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 23552 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 27508 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 6624 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 13524 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 31648 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 17112 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 7636 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 25208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 16192 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 10212 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 28796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0719_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 17572 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 32292 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 31188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 32476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 29072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 33396 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 14536 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 6716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 31556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 9108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 15824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 32292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 28428 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 12512 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 18584 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 20148 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 13892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0755_
timestamp 1667941163
transform 1 0 5520 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 26404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 28796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 27784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 6164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 27232 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 32292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 6532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0771_
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 27416 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 19504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 32660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 35788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 24748 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0787_
timestamp 1667941163
transform 1 0 13984 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 34224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 15088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 34224 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 33580 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 31464 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0794_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0795_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2760 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 16836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 4968 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 17940 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 16468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 16836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 16008 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 15364 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 15180 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 2852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 13432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_
timestamp 1667941163
transform 1 0 1840 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 17480 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 18124 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 15824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 18584 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 15180 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 17480 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 15364 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 13892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 14904 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 2852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 5244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 10304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 6532 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 12788 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 9752 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0828_
timestamp 1667941163
transform 1 0 1840 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 4968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 14720 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 7360 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 14536 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 17480 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 14720 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 5888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 2760 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 14076 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 10396 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 10948 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 2024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0850_
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 15548 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 16192 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 3496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 1564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 2300 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 2208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 14996 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 14536 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 16836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0861_
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 2760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 7176 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 3956 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 5612 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 5612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 4968 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 17480 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1667941163
transform 1 0 18768 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 17020 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 18124 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 17480 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 17480 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0878_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11224 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0879_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6992 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0880_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7820 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0881_
timestamp 1667941163
transform 1 0 11500 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0882_
timestamp 1667941163
transform 1 0 6624 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0883_
timestamp 1667941163
transform 1 0 6532 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0885_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 6808 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 9200 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0888_
timestamp 1667941163
transform 1 0 8188 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0891_
timestamp 1667941163
transform 1 0 7820 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0893_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 8832 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 7728 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 9108 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0900_
timestamp 1667941163
transform 1 0 2668 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 6992 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 4600 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 2668 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 5152 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0906_
timestamp 1667941163
transform 1 0 1564 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 1840 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 1564 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0912_
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 3956 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0916_
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 3312 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 9292 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0921_
timestamp 1667941163
transform 1 0 9108 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0922_
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0923_
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0924_
timestamp 1667941163
transform 1 0 6624 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 4232 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 5888 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0930_
timestamp 1667941163
transform 1 0 9292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 14168 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 8188 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 2024 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 6716 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0935_
timestamp 1667941163
transform 1 0 11500 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0936_
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0937_
timestamp 1667941163
transform 1 0 4416 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0938_
timestamp 1667941163
transform 1 0 10672 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0939_
timestamp 1667941163
transform 1 0 11868 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0940_
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0941_
timestamp 1667941163
transform 1 0 3036 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0942_
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0943_
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 4048 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0948_
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0949_
timestamp 1667941163
transform 1 0 6992 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 4416 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 6808 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1667941163
transform 1 0 6716 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0953_
timestamp 1667941163
transform 1 0 6808 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 35880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 15180 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 34776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 14444 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 35328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 15732 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 34224 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 4324 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 34408 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 33396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 12144 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 13432 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 13156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 27692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1030_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1031__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10120 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1032_
timestamp 1667941163
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1033_
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1034_
timestamp 1667941163
transform 1 0 12880 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1035_
timestamp 1667941163
transform 1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1036_
timestamp 1667941163
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1037_
timestamp 1667941163
transform 1 0 14444 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1037__101
timestamp 1667941163
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1038_
timestamp 1667941163
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1039_
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1040_
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1041_
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1042_
timestamp 1667941163
transform 1 0 16836 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1043__102
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1043_
timestamp 1667941163
transform 1 0 16192 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 17848 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 11684 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 17664 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 9752 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1049__103
timestamp 1667941163
transform 1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1050_
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 11408 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 13984 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1054_
timestamp 1667941163
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1055__104
timestamp 1667941163
transform 1 0 20884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1057_
timestamp 1667941163
transform 1 0 16100 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 18032 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 15824 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1061__105
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 12512 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 15088 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 15180 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 12604 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 17020 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1067__106
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 11684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 10856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1073__107
timestamp 1667941163
transform 1 0 9016 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 11960 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 14352 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 9384 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1078_
timestamp 1667941163
transform 1 0 17204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1079__108
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 11500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1081_
timestamp 1667941163
transform 1 0 14168 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1084_
timestamp 1667941163
transform 1 0 10948 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1085__109
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 14904 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 14352 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 9568 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 13156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 9016 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1091__110
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 22080 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 20516 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1097__111
timestamp 1667941163
transform 1 0 20148 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 19320 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 22080 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 19872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 14904 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1103__112
timestamp 1667941163
transform 1 0 18492 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 12788 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 12788 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 18216 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1107_
timestamp 1667941163
transform 1 0 9200 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 21712 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1109__113
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1110_
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1113_
timestamp 1667941163
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 22908 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1115__114
timestamp 1667941163
transform 1 0 22632 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 23092 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 21344 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 22724 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 17112 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1121__115
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 21252 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 17296 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 15456 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 12512 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1127__116
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 23092 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 23000 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform 1 0 23276 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1133__117
timestamp 1667941163
transform 1 0 20332 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1139__118
timestamp 1667941163
transform 1 0 7728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1140_
timestamp 1667941163
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 10396 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1145__119
timestamp 1667941163
transform 1 0 17204 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 20148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 19504 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 20608 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1150_
timestamp 1667941163
transform 1 0 9936 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1150__120
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 4784 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 11408 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1153_
timestamp 1667941163
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1154__121
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 8280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 14628 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 9292 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 23828 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1158__122
timestamp 1667941163
transform 1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1159_
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 22632 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 22080 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1162__123
timestamp 1667941163
transform 1 0 17480 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 9384 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 16652 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 12972 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1166__124
timestamp 1667941163
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1167_
timestamp 1667941163
transform 1 0 19872 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 12972 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 18124 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1170__125
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 10396 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1174_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17296 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1174__126
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1176_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1178__127
timestamp 1667941163
transform 1 0 8372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 4048 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1180_
timestamp 1667941163
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1182__128
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1186__129
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 14444 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1190__130
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 13984 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1194__131
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 17296 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1196_
timestamp 1667941163
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1198_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1198__132
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 19228 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1200_
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1202__133
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1202_
timestamp 1667941163
transform 1 0 14168 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1203_
timestamp 1667941163
transform 1 0 19596 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1204_
timestamp 1667941163
transform 1 0 14628 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1205_
timestamp 1667941163
transform 1 0 20148 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1206__134
timestamp 1667941163
transform 1 0 25024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 22540 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1207_
timestamp 1667941163
transform 1 0 18676 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 20700 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1209_
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1210__135
timestamp 1667941163
transform 1 0 23736 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 22356 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 20976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 21620 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 16100 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1214__136
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 17664 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 22356 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1218__137
timestamp 1667941163
transform 1 0 25760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 24472 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 25392 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 25484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 18308 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 38088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 1564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 14720 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 2944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 16376 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 10120 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 5704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 2 nsew signal input
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 3 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 4 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 5 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 6 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 7 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 8 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 9 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 10 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 11 nsew signal input
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 12 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 13 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 14 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 15 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 16 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 17 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 18 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 19 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 20 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 21 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 22 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 23 nsew signal tristate
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 24 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 26 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 27 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 28 nsew signal tristate
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 29 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 30 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 32 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 33 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 34 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 35 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 36 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 37 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 38 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 pReset
port 78 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 prog_clk
port 79 nsew signal input
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 80 nsew signal input
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 81 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 82 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 83 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 84 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 85 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 86 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 87 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 88 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 89 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 90 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 91 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 96 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 97 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 98 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 99 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 vssd1
port 101 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 10120 33286 10120 33286 0 _0000_
rlabel via2 14398 31875 14398 31875 0 _0001_
rlabel metal1 6716 33286 6716 33286 0 _0002_
rlabel metal2 12926 30141 12926 30141 0 _0003_
rlabel metal3 7360 32708 7360 32708 0 _0004_
rlabel metal1 4324 32198 4324 32198 0 _0005_
rlabel metal1 13294 30260 13294 30260 0 _0006_
rlabel via3 9269 32300 9269 32300 0 _0007_
rlabel metal1 7406 31858 7406 31858 0 _0008_
rlabel metal1 3871 31722 3871 31722 0 _0009_
rlabel metal2 3082 25959 3082 25959 0 _0010_
rlabel metal1 17158 33014 17158 33014 0 _0011_
rlabel metal1 6079 33898 6079 33898 0 _0012_
rlabel metal1 6072 32742 6072 32742 0 _0013_
rlabel metal2 4738 29852 4738 29852 0 _0014_
rlabel metal2 9706 31977 9706 31977 0 _0015_
rlabel metal2 2438 24650 2438 24650 0 _0016_
rlabel metal1 14260 31450 14260 31450 0 _0017_
rlabel metal1 10856 32538 10856 32538 0 _0018_
rlabel metal2 8970 36108 8970 36108 0 _0019_
rlabel via3 4853 35972 4853 35972 0 _0020_
rlabel metal1 9752 32810 9752 32810 0 _0021_
rlabel metal1 10373 33354 10373 33354 0 _0022_
rlabel metal1 2392 32198 2392 32198 0 _0023_
rlabel metal1 4462 31790 4462 31790 0 _0024_
rlabel metal2 15686 32283 15686 32283 0 _0025_
rlabel metal1 16146 31994 16146 31994 0 _0026_
rlabel metal3 7659 36108 7659 36108 0 _0027_
rlabel metal3 15663 35972 15663 35972 0 _0028_
rlabel metal2 2438 30345 2438 30345 0 _0029_
rlabel metal1 2254 23834 2254 23834 0 _0030_
rlabel metal1 14812 32742 14812 32742 0 _0031_
rlabel via2 2346 23035 2346 23035 0 _0032_
rlabel via2 14398 32317 14398 32317 0 _0033_
rlabel metal1 16928 31994 16928 31994 0 _0034_
rlabel metal1 4830 34170 4830 34170 0 _0035_
rlabel metal2 12650 36601 12650 36601 0 _0036_
rlabel metal1 3634 33082 3634 33082 0 _0037_
rlabel metal1 5796 32266 5796 32266 0 _0038_
rlabel via2 4462 36805 4462 36805 0 _0039_
rlabel metal1 5888 32402 5888 32402 0 _0040_
rlabel metal2 5106 27982 5106 27982 0 _0041_
rlabel metal1 3871 27370 3871 27370 0 _0042_
rlabel metal2 2898 27319 2898 27319 0 _0043_
rlabel metal1 4002 30566 4002 30566 0 _0044_
rlabel metal2 10534 35105 10534 35105 0 _0045_
rlabel metal2 15502 36482 15502 36482 0 _0046_
rlabel metal2 13202 35513 13202 35513 0 _0047_
rlabel metal2 15686 35309 15686 35309 0 _0048_
rlabel metal2 17618 36380 17618 36380 0 _0049_
rlabel metal1 14582 35768 14582 35768 0 _0050_
rlabel metal1 12650 32919 12650 32919 0 _0051_
rlabel metal1 7353 28118 7353 28118 0 _0052_
rlabel metal1 17986 34170 17986 34170 0 _0053_
rlabel metal1 16238 34986 16238 34986 0 _0054_
rlabel metal1 8970 30056 8970 30056 0 _0055_
rlabel metal2 13754 33796 13754 33796 0 _0056_
rlabel metal1 14582 31178 14582 31178 0 _0057_
rlabel metal1 10534 29655 10534 29655 0 _0058_
rlabel metal1 4324 23834 4324 23834 0 _0059_
rlabel metal1 11139 27030 11139 27030 0 _0060_
rlabel metal1 14490 32266 14490 32266 0 _0061_
rlabel metal1 14858 27608 14858 27608 0 _0062_
rlabel metal2 18262 35156 18262 35156 0 _0063_
rlabel metal1 9460 33490 9460 33490 0 _0064_
rlabel metal2 18722 33456 18722 33456 0 _0065_
rlabel metal2 16974 35054 16974 35054 0 _0066_
rlabel metal1 7406 24106 7406 24106 0 _0067_
rlabel metal1 14720 33286 14720 33286 0 _0068_
rlabel metal2 17618 33898 17618 33898 0 _0069_
rlabel metal2 11546 32708 11546 32708 0 _0070_
rlabel metal1 10350 31450 10350 31450 0 _0071_
rlabel metal1 14030 30124 14030 30124 0 _0072_
rlabel via2 8142 32011 8142 32011 0 _0073_
rlabel metal1 4554 23290 4554 23290 0 _0074_
rlabel metal1 5566 32742 5566 32742 0 _0075_
rlabel metal2 24978 28764 24978 28764 0 _0076_
rlabel metal1 24886 30090 24886 30090 0 _0077_
rlabel metal1 22218 32844 22218 32844 0 _0078_
rlabel metal2 16054 33796 16054 33796 0 _0079_
rlabel metal1 21022 19380 21022 19380 0 _0080_
rlabel metal1 21597 29274 21597 29274 0 _0081_
rlabel metal1 17066 32436 17066 32436 0 _0082_
rlabel metal2 24610 27268 24610 27268 0 _0083_
rlabel metal2 19642 30906 19642 30906 0 _0084_
rlabel metal1 10994 23222 10994 23222 0 _0085_
rlabel metal1 18446 16762 18446 16762 0 _0086_
rlabel metal2 22862 17476 22862 17476 0 _0087_
rlabel metal2 19642 15674 19642 15674 0 _0088_
rlabel metal1 7314 19788 7314 19788 0 _0089_
rlabel metal2 13938 14892 13938 14892 0 _0090_
rlabel metal1 10304 15470 10304 15470 0 _0091_
rlabel metal2 13570 14790 13570 14790 0 _0092_
rlabel metal2 17066 29308 17066 29308 0 _0093_
rlabel metal1 19458 26962 19458 26962 0 _0094_
rlabel metal1 10948 16218 10948 16218 0 _0095_
rlabel metal1 18538 16116 18538 16116 0 _0096_
rlabel metal1 5428 24378 5428 24378 0 _0097_
rlabel metal1 6256 30362 6256 30362 0 _0098_
rlabel metal1 6624 22406 6624 22406 0 _0099_
rlabel metal1 10718 18768 10718 18768 0 _0100_
rlabel metal1 16744 22406 16744 22406 0 _0101_
rlabel metal1 8602 28560 8602 28560 0 _0102_
rlabel metal2 18906 31994 18906 31994 0 _0103_
rlabel metal2 10534 21590 10534 21590 0 _0104_
rlabel metal1 9844 31790 9844 31790 0 _0105_
rlabel metal1 16928 20434 16928 20434 0 _0106_
rlabel metal2 23690 19108 23690 19108 0 _0107_
rlabel metal2 25070 20740 25070 20740 0 _0108_
rlabel metal1 7636 17646 7636 17646 0 _0109_
rlabel metal1 17940 14858 17940 14858 0 _0110_
rlabel metal1 6394 24378 6394 24378 0 _0111_
rlabel metal1 10212 32402 10212 32402 0 _0112_
rlabel metal1 21022 24786 21022 24786 0 _0113_
rlabel metal2 17894 23052 17894 23052 0 _0114_
rlabel metal1 18446 25840 18446 25840 0 _0115_
rlabel metal2 10074 18428 10074 18428 0 _0116_
rlabel metal1 7958 19380 7958 19380 0 _0117_
rlabel metal1 8832 19482 8832 19482 0 _0118_
rlabel metal2 26358 24582 26358 24582 0 _0119_
rlabel metal2 21482 23868 21482 23868 0 _0120_
rlabel metal2 20562 24378 20562 24378 0 _0121_
rlabel metal1 26082 26316 26082 26316 0 _0122_
rlabel metal1 17802 28730 17802 28730 0 _0123_
rlabel metal2 24610 23494 24610 23494 0 _0124_
rlabel metal1 14444 24174 14444 24174 0 _0125_
rlabel metal1 16514 30668 16514 30668 0 _0126_
rlabel metal2 19642 27642 19642 27642 0 _0127_
rlabel metal1 24150 26350 24150 26350 0 _0128_
rlabel metal1 24610 22644 24610 22644 0 _0129_
rlabel metal1 23966 21488 23966 21488 0 _0130_
rlabel metal1 18630 19482 18630 19482 0 _0131_
rlabel metal2 22862 21267 22862 21267 0 _0132_
rlabel metal1 23138 20978 23138 20978 0 _0133_
rlabel metal1 9798 22406 9798 22406 0 _0134_
rlabel metal2 13754 29818 13754 29818 0 _0135_
rlabel metal1 17664 26010 17664 26010 0 _0136_
rlabel metal1 20286 16524 20286 16524 0 _0137_
rlabel metal1 22770 24786 22770 24786 0 _0138_
rlabel metal1 21758 18768 21758 18768 0 _0139_
rlabel metal2 12466 19482 12466 19482 0 _0140_
rlabel metal1 10488 19346 10488 19346 0 _0141_
rlabel metal1 18446 15470 18446 15470 0 _0142_
rlabel metal1 12282 20774 12282 20774 0 _0143_
rlabel metal1 10350 25296 10350 25296 0 _0144_
rlabel metal1 10534 20400 10534 20400 0 _0145_
rlabel metal2 8602 18938 8602 18938 0 _0146_
rlabel metal1 16054 29172 16054 29172 0 _0147_
rlabel metal1 19688 26010 19688 26010 0 _0148_
rlabel metal2 13570 23358 13570 23358 0 _0149_
rlabel metal1 11316 20910 11316 20910 0 _0150_
rlabel metal1 8648 21522 8648 21522 0 _0151_
rlabel metal2 9614 24531 9614 24531 0 _0152_
rlabel metal1 9016 18258 9016 18258 0 _0153_
rlabel metal2 18078 14586 18078 14586 0 _0154_
rlabel metal1 12098 26554 12098 26554 0 _0155_
rlabel metal1 12558 24786 12558 24786 0 _0156_
rlabel metal1 12558 25296 12558 25296 0 _0157_
rlabel metal1 18814 28560 18814 28560 0 _0158_
rlabel metal2 15226 28526 15226 28526 0 _0159_
rlabel metal1 17526 26452 17526 26452 0 _0160_
rlabel metal1 13156 26350 13156 26350 0 _0161_
rlabel metal1 6072 26962 6072 26962 0 _0162_
rlabel metal1 9752 23290 9752 23290 0 _0163_
rlabel metal2 16054 21692 16054 21692 0 _0164_
rlabel metal2 14214 23868 14214 23868 0 _0165_
rlabel metal1 15870 19482 15870 19482 0 _0166_
rlabel metal2 15502 14790 15502 14790 0 _0167_
rlabel metal1 12696 15130 12696 15130 0 _0168_
rlabel metal2 16330 15708 16330 15708 0 _0169_
rlabel metal2 8142 18428 8142 18428 0 _0170_
rlabel metal1 7820 20434 7820 20434 0 _0171_
rlabel metal1 1932 33966 1932 33966 0 _0172_
rlabel metal1 15318 32402 15318 32402 0 _0173_
rlabel metal1 1794 33898 1794 33898 0 _0174_
rlabel metal1 14628 31790 14628 31790 0 _0175_
rlabel metal1 14306 33490 14306 33490 0 _0176_
rlabel metal1 2346 24140 2346 24140 0 _0177_
rlabel metal1 2116 23698 2116 23698 0 _0178_
rlabel metal2 13110 31076 13110 31076 0 _0179_
rlabel metal1 9476 19754 9476 19754 0 _0180_
rlabel metal1 8050 20570 8050 20570 0 _0181_
rlabel metal1 10718 18156 10718 18156 0 _0182_
rlabel metal1 11362 18632 11362 18632 0 _0183_
rlabel metal2 13110 17748 13110 17748 0 _0184_
rlabel metal2 7498 25636 7498 25636 0 _0185_
rlabel metal2 16146 17170 16146 17170 0 _0186_
rlabel metal2 13570 16184 13570 16184 0 _0187_
rlabel metal1 15134 14858 15134 14858 0 _0188_
rlabel metal1 15042 15674 15042 15674 0 _0189_
rlabel metal1 13110 15980 13110 15980 0 _0190_
rlabel metal1 14628 15130 14628 15130 0 _0191_
rlabel metal2 17066 23256 17066 23256 0 _0192_
rlabel metal1 16422 21012 16422 21012 0 _0193_
rlabel metal1 17986 21420 17986 21420 0 _0194_
rlabel metal1 16698 23834 16698 23834 0 _0195_
rlabel metal1 10902 21454 10902 21454 0 _0196_
rlabel metal1 17894 20876 17894 20876 0 _0197_
rlabel metal1 7774 27098 7774 27098 0 _0198_
rlabel metal1 11868 22610 11868 22610 0 _0199_
rlabel metal1 16460 26418 16460 26418 0 _0200_
rlabel metal1 11362 27370 11362 27370 0 _0201_
rlabel metal1 7682 23018 7682 23018 0 _0202_
rlabel metal1 13616 24378 13616 24378 0 _0203_
rlabel metal1 15824 26894 15824 26894 0 _0204_
rlabel metal1 20884 25806 20884 25806 0 _0205_
rlabel metal1 18538 27506 18538 27506 0 _0206_
rlabel metal1 16008 27506 16008 27506 0 _0207_
rlabel metal2 22218 27370 22218 27370 0 _0208_
rlabel metal2 18262 27948 18262 27948 0 _0209_
rlabel metal2 16054 24344 16054 24344 0 _0210_
rlabel metal1 16146 25398 16146 25398 0 _0211_
rlabel metal1 12834 25874 12834 25874 0 _0212_
rlabel metal1 12650 24684 12650 24684 0 _0213_
rlabel metal2 15870 28220 15870 28220 0 _0214_
rlabel metal1 15410 25908 15410 25908 0 _0215_
rlabel metal1 11086 18088 11086 18088 0 _0216_
rlabel metal2 17894 15844 17894 15844 0 _0217_
rlabel metal1 11868 23698 11868 23698 0 _0218_
rlabel metal2 11914 20434 11914 20434 0 _0219_
rlabel metal1 17526 14586 17526 14586 0 _0220_
rlabel metal1 9798 22746 9798 22746 0 _0221_
rlabel metal2 11730 21267 11730 21267 0 _0222_
rlabel metal1 8924 21658 8924 21658 0 _0223_
rlabel metal1 13984 23154 13984 23154 0 _0224_
rlabel metal1 13248 21930 13248 21930 0 _0225_
rlabel metal1 9568 23154 9568 23154 0 _0226_
rlabel metal2 11822 24140 11822 24140 0 _0227_
rlabel metal1 17112 28050 17112 28050 0 _0228_
rlabel metal1 20562 25330 20562 25330 0 _0229_
rlabel metal1 10718 17714 10718 17714 0 _0230_
rlabel metal1 14352 26962 14352 26962 0 _0231_
rlabel metal2 20194 29308 20194 29308 0 _0232_
rlabel metal1 13110 20400 13110 20400 0 _0233_
rlabel metal2 11178 24820 11178 24820 0 _0234_
rlabel metal2 10902 20060 10902 20060 0 _0235_
rlabel metal1 14582 22644 14582 22644 0 _0236_
rlabel metal1 9338 24242 9338 24242 0 _0237_
rlabel metal2 13386 20196 13386 20196 0 _0238_
rlabel metal1 7912 21114 7912 21114 0 _0239_
rlabel metal1 11040 19414 11040 19414 0 _0240_
rlabel metal1 18308 15674 18308 15674 0 _0241_
rlabel metal2 13570 19414 13570 19414 0 _0242_
rlabel metal1 15548 20434 15548 20434 0 _0243_
rlabel metal1 16100 14586 16100 14586 0 _0244_
rlabel metal1 16468 23290 16468 23290 0 _0245_
rlabel metal2 22310 23800 22310 23800 0 _0246_
rlabel metal1 21160 18938 21160 18938 0 _0247_
rlabel metal1 19826 16762 19826 16762 0 _0248_
rlabel metal1 22310 23800 22310 23800 0 _0249_
rlabel metal2 20930 19210 20930 19210 0 _0250_
rlabel metal1 20838 17306 20838 17306 0 _0251_
rlabel metal2 15134 28560 15134 28560 0 _0252_
rlabel metal2 18722 25636 18722 25636 0 _0253_
rlabel metal1 12650 19720 12650 19720 0 _0254_
rlabel metal2 13018 28424 13018 28424 0 _0255_
rlabel metal1 17986 25330 17986 25330 0 _0256_
rlabel metal1 8740 23766 8740 23766 0 _0257_
rlabel metal1 22011 20842 22011 20842 0 _0258_
rlabel metal2 21022 21284 21022 21284 0 _0259_
rlabel metal1 18768 20298 18768 20298 0 _0260_
rlabel metal1 19596 20026 19596 20026 0 _0261_
rlabel metal2 21206 22916 21206 22916 0 _0262_
rlabel metal1 17434 19924 17434 19924 0 _0263_
rlabel metal1 23322 21930 23322 21930 0 _0264_
rlabel metal1 22586 21454 22586 21454 0 _0265_
rlabel metal1 23598 25330 23598 25330 0 _0266_
rlabel metal1 24012 24854 24012 24854 0 _0267_
rlabel metal1 21206 22066 21206 22066 0 _0268_
rlabel metal1 22908 28594 22908 28594 0 _0269_
rlabel metal1 16836 29682 16836 29682 0 _0270_
rlabel metal1 21482 27370 21482 27370 0 _0271_
rlabel metal1 16054 24378 16054 24378 0 _0272_
rlabel metal1 15548 30226 15548 30226 0 _0273_
rlabel metal2 22218 28764 22218 28764 0 _0274_
rlabel metal2 12742 28356 12742 28356 0 _0275_
rlabel metal1 19780 27370 19780 27370 0 _0276_
rlabel metal1 23966 23630 23966 23630 0 _0277_
rlabel metal1 24610 26554 24610 26554 0 _0278_
rlabel metal1 19642 28424 19642 28424 0 _0279_
rlabel metal1 23552 24242 23552 24242 0 _0280_
rlabel metal1 24334 22542 24334 22542 0 _0281_
rlabel metal2 20930 23086 20930 23086 0 _0282_
rlabel metal1 20240 23154 20240 23154 0 _0283_
rlabel metal1 25208 24242 25208 24242 0 _0284_
rlabel metal2 22770 23494 22770 23494 0 _0285_
rlabel metal1 17802 22678 17802 22678 0 _0286_
rlabel metal2 23598 26860 23598 26860 0 _0287_
rlabel metal1 11960 19414 11960 19414 0 _0288_
rlabel metal2 13202 21216 13202 21216 0 _0289_
rlabel metal1 10350 18394 10350 18394 0 _0290_
rlabel metal1 10534 16490 10534 16490 0 _0291_
rlabel metal1 12857 21998 12857 21998 0 _0292_
rlabel metal1 10534 16218 10534 16218 0 _0293_
rlabel metal1 18538 22712 18538 22712 0 _0294_
rlabel metal1 18124 23698 18124 23698 0 _0295_
rlabel metal1 20700 23698 20700 23698 0 _0296_
rlabel metal1 19872 22678 19872 22678 0 _0297_
rlabel metal1 16192 23222 16192 23222 0 _0298_
rlabel metal2 20838 29070 20838 29070 0 _0299_
rlabel metal1 10212 30770 10212 30770 0 _0300_
rlabel metal2 5014 29580 5014 29580 0 _0301_
rlabel metal2 11638 30226 11638 30226 0 _0302_
rlabel metal2 8142 27812 8142 27812 0 _0303_
rlabel metal1 20332 16422 20332 16422 0 _0304_
rlabel metal2 8510 17340 8510 17340 0 _0305_
rlabel metal1 14904 14586 14904 14586 0 _0306_
rlabel metal1 9016 17714 9016 17714 0 _0307_
rlabel metal2 24058 20638 24058 20638 0 _0308_
rlabel metal2 23506 19380 23506 19380 0 _0309_
rlabel metal1 23782 20026 23782 20026 0 _0310_
rlabel metal2 22954 19108 22954 19108 0 _0311_
rlabel metal1 18998 20536 18998 20536 0 _0312_
rlabel metal1 9568 31926 9568 31926 0 _0313_
rlabel metal1 16238 22474 16238 22474 0 _0314_
rlabel metal1 14490 26248 14490 26248 0 _0315_
rlabel metal1 13202 20808 13202 20808 0 _0316_
rlabel metal1 19412 31926 19412 31926 0 _0317_
rlabel metal2 13202 25704 13202 25704 0 _0318_
rlabel metal1 18538 30362 18538 30362 0 _0319_
rlabel metal1 9016 28730 9016 28730 0 _0320_
rlabel metal2 17158 21760 17158 21760 0 _0321_
rlabel metal2 11914 27710 11914 27710 0 _0322_
rlabel metal2 17250 25534 17250 25534 0 _0323_
rlabel metal1 15226 18802 15226 18802 0 _0324_
rlabel metal1 7544 19890 7544 19890 0 _0325_
rlabel metal1 13754 15674 13754 15674 0 _0326_
rlabel metal1 9338 22100 9338 22100 0 _0327_
rlabel metal1 7636 29682 7636 29682 0 _0328_
rlabel metal2 4922 26044 4922 26044 0 _0329_
rlabel metal1 5566 29172 5566 29172 0 _0330_
rlabel metal1 7038 25466 7038 25466 0 _0331_
rlabel metal2 18354 17544 18354 17544 0 _0332_
rlabel metal1 12466 17068 12466 17068 0 _0333_
rlabel metal1 16514 18326 16514 18326 0 _0334_
rlabel metal1 10902 16558 10902 16558 0 _0335_
rlabel metal2 20930 26350 20930 26350 0 _0336_
rlabel metal1 17986 29036 17986 29036 0 _0337_
rlabel metal1 19642 26248 19642 26248 0 _0338_
rlabel metal2 14674 27132 14674 27132 0 _0339_
rlabel metal1 13570 15096 13570 15096 0 _0340_
rlabel metal1 10948 15674 10948 15674 0 _0341_
rlabel metal2 13294 15504 13294 15504 0 _0342_
rlabel metal2 9338 15708 9338 15708 0 _0343_
rlabel metal2 15318 14756 15318 14756 0 _0344_
rlabel metal1 17526 15572 17526 15572 0 _0345_
rlabel metal1 16284 13498 16284 13498 0 _0346_
rlabel metal1 17342 14042 17342 14042 0 _0347_
rlabel metal1 22448 17850 22448 17850 0 _0348_
rlabel metal1 18768 17850 18768 17850 0 _0349_
rlabel metal1 21114 17238 21114 17238 0 _0350_
rlabel metal1 19412 17714 19412 17714 0 _0351_
rlabel metal1 13754 19448 13754 19448 0 _0352_
rlabel metal1 19642 30294 19642 30294 0 _0353_
rlabel metal2 12374 23902 12374 23902 0 _0354_
rlabel metal1 20010 32198 20010 32198 0 _0355_
rlabel metal1 22770 25976 22770 25976 0 _0356_
rlabel metal1 17756 32266 17756 32266 0 _0357_
rlabel metal1 22080 28118 22080 28118 0 _0358_
rlabel metal2 14030 33762 14030 33762 0 _0359_
rlabel metal2 22034 28254 22034 28254 0 _0360_
rlabel metal1 21022 19482 21022 19482 0 _0361_
rlabel metal2 22678 25772 22678 25772 0 _0362_
rlabel metal2 22310 19346 22310 19346 0 _0363_
rlabel metal1 16330 33864 16330 33864 0 _0364_
rlabel metal2 22218 32300 22218 32300 0 _0365_
rlabel metal2 17894 33694 17894 33694 0 _0366_
rlabel metal2 22586 32572 22586 32572 0 _0367_
rlabel metal2 25622 30702 25622 30702 0 _0368_
rlabel metal1 24748 26962 24748 26962 0 _0369_
rlabel metal1 25622 30600 25622 30600 0 _0370_
rlabel metal1 25484 31314 25484 31314 0 _0371_
rlabel metal2 38134 6239 38134 6239 0 ccff_head
rlabel via2 38226 33371 38226 33371 0 ccff_tail
rlabel metal1 22724 37230 22724 37230 0 chanx_right_in[0]
rlabel metal1 37766 36142 37766 36142 0 chanx_right_in[10]
rlabel metal3 1234 12308 1234 12308 0 chanx_right_in[11]
rlabel metal2 34822 1588 34822 1588 0 chanx_right_in[12]
rlabel metal1 17388 36346 17388 36346 0 chanx_right_in[13]
rlabel metal1 38180 36754 38180 36754 0 chanx_right_in[14]
rlabel metal2 29026 1588 29026 1588 0 chanx_right_in[15]
rlabel metal3 1234 7548 1234 7548 0 chanx_right_in[16]
rlabel metal1 1748 23086 1748 23086 0 chanx_right_in[17]
rlabel metal2 10350 1588 10350 1588 0 chanx_right_in[18]
rlabel metal2 19366 37196 19366 37196 0 chanx_right_in[1]
rlabel metal2 4554 1588 4554 1588 0 chanx_right_in[2]
rlabel metal3 1234 20468 1234 20468 0 chanx_right_in[3]
rlabel metal3 1234 17748 1234 17748 0 chanx_right_in[4]
rlabel metal2 38318 28883 38318 28883 0 chanx_right_in[5]
rlabel metal1 18216 37230 18216 37230 0 chanx_right_in[6]
rlabel metal2 33534 1588 33534 1588 0 chanx_right_in[7]
rlabel metal3 1234 25228 1234 25228 0 chanx_right_in[8]
rlabel metal1 14398 30328 14398 30328 0 chanx_right_in[9]
rlabel metal2 1794 27183 1794 27183 0 chanx_right_out[0]
rlabel metal2 22586 1520 22586 1520 0 chanx_right_out[10]
rlabel metal2 14858 1520 14858 1520 0 chanx_right_out[11]
rlabel metal2 39330 1520 39330 1520 0 chanx_right_out[12]
rlabel metal3 1234 1428 1234 1428 0 chanx_right_out[13]
rlabel metal2 38226 20621 38226 20621 0 chanx_right_out[14]
rlabel metal1 24656 37094 24656 37094 0 chanx_right_out[15]
rlabel metal1 14030 37094 14030 37094 0 chanx_right_out[16]
rlabel metal2 38226 36941 38226 36941 0 chanx_right_out[17]
rlabel metal2 16790 1520 16790 1520 0 chanx_right_out[18]
rlabel metal3 1234 15708 1234 15708 0 chanx_right_out[1]
rlabel metal2 38226 34833 38226 34833 0 chanx_right_out[2]
rlabel metal1 15640 37094 15640 37094 0 chanx_right_out[3]
rlabel metal2 38226 8857 38226 8857 0 chanx_right_out[4]
rlabel metal2 38226 12461 38226 12461 0 chanx_right_out[5]
rlabel metal1 16928 37094 16928 37094 0 chanx_right_out[6]
rlabel metal1 10258 36346 10258 36346 0 chanx_right_out[7]
rlabel metal2 25806 1520 25806 1520 0 chanx_right_out[8]
rlabel metal2 9062 1520 9062 1520 0 chanx_right_out[9]
rlabel metal2 38318 30107 38318 30107 0 chany_top_in[0]
rlabel metal2 38042 1367 38042 1367 0 chany_top_in[10]
rlabel metal2 38318 15895 38318 15895 0 chany_top_in[11]
rlabel metal1 29486 37230 29486 37230 0 chany_top_in[12]
rlabel metal2 12558 37213 12558 37213 0 chany_top_in[13]
rlabel metal2 36938 2227 36938 2227 0 chany_top_in[14]
rlabel metal2 38318 32215 38318 32215 0 chany_top_in[15]
rlabel metal1 36846 37230 36846 37230 0 chany_top_in[16]
rlabel metal2 21298 38226 21298 38226 0 chany_top_in[17]
rlabel metal3 1234 19108 1234 19108 0 chany_top_in[18]
rlabel metal2 38318 7701 38318 7701 0 chany_top_in[1]
rlabel metal3 1234 22508 1234 22508 0 chany_top_in[2]
rlabel metal3 1234 2788 1234 2788 0 chany_top_in[3]
rlabel metal1 25944 37230 25944 37230 0 chany_top_in[4]
rlabel metal3 1924 28628 1924 28628 0 chany_top_in[5]
rlabel metal2 30314 1588 30314 1588 0 chany_top_in[6]
rlabel metal1 33672 37230 33672 37230 0 chany_top_in[7]
rlabel metal3 1234 9588 1234 9588 0 chany_top_in[8]
rlabel metal2 2622 1588 2622 1588 0 chany_top_in[9]
rlabel metal2 11638 1520 11638 1520 0 chany_top_out[0]
rlabel metal2 36110 1520 36110 1520 0 chany_top_out[10]
rlabel via2 38226 17051 38226 17051 0 chany_top_out[11]
rlabel metal2 38226 11101 38226 11101 0 chany_top_out[12]
rlabel metal3 1234 6188 1234 6188 0 chany_top_out[13]
rlabel metal2 1794 33235 1794 33235 0 chany_top_out[14]
rlabel via2 38226 2805 38226 2805 0 chany_top_out[15]
rlabel metal1 6670 34442 6670 34442 0 chany_top_out[16]
rlabel metal2 38226 14297 38226 14297 0 chany_top_out[17]
rlabel metal2 38226 25177 38226 25177 0 chany_top_out[18]
rlabel metal2 31602 1520 31602 1520 0 chany_top_out[1]
rlabel via2 38226 27285 38226 27285 0 chany_top_out[2]
rlabel metal1 5888 35802 5888 35802 0 chany_top_out[3]
rlabel metal3 1234 23868 1234 23868 0 chany_top_out[4]
rlabel metal2 19366 1520 19366 1520 0 chany_top_out[5]
rlabel metal2 46 1792 46 1792 0 chany_top_out[6]
rlabel metal2 23874 1520 23874 1520 0 chany_top_out[7]
rlabel metal1 9338 36040 9338 36040 0 chany_top_out[8]
rlabel metal1 20148 37094 20148 37094 0 chany_top_out[9]
rlabel metal1 15640 26350 15640 26350 0 mem_right_track_0.DFFR_0_.D
rlabel metal1 12489 20910 12489 20910 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 12972 33422 12972 33422 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 2293 28934 2293 28934 0 mem_right_track_10.DFFR_0_.D
rlabel metal2 1886 28934 1886 28934 0 mem_right_track_10.DFFR_0_.Q
rlabel metal3 17204 25160 17204 25160 0 mem_right_track_10.DFFR_1_.Q
rlabel metal1 19642 28016 19642 28016 0 mem_right_track_12.DFFR_0_.Q
rlabel metal1 14858 30702 14858 30702 0 mem_right_track_12.DFFR_1_.Q
rlabel metal1 16054 25330 16054 25330 0 mem_right_track_14.DFFR_0_.Q
rlabel via2 1886 28101 1886 28101 0 mem_right_track_14.DFFR_1_.Q
rlabel metal3 2277 31756 2277 31756 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 21206 24208 21206 24208 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 9246 19312 9246 19312 0 mem_right_track_18.DFFR_0_.Q
rlabel metal1 13432 37094 13432 37094 0 mem_right_track_18.DFFR_1_.Q
rlabel metal1 16882 16082 16882 16082 0 mem_right_track_2.DFFR_0_.Q
rlabel metal2 10994 21420 10994 21420 0 mem_right_track_2.DFFR_1_.Q
rlabel via2 13662 36533 13662 36533 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 13754 14433 13754 14433 0 mem_right_track_20.DFFR_1_.Q
rlabel via2 17066 13923 17066 13923 0 mem_right_track_22.DFFR_0_.Q
rlabel metal4 15180 14824 15180 14824 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 18722 17697 18722 17697 0 mem_right_track_24.DFFR_0_.Q
rlabel via1 1879 27642 1879 27642 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 18814 32334 18814 32334 0 mem_right_track_26.DFFR_0_.Q
rlabel metal2 5842 26112 5842 26112 0 mem_right_track_26.DFFR_1_.Q
rlabel metal1 14582 32844 14582 32844 0 mem_right_track_28.DFFR_0_.Q
rlabel metal2 21942 28577 21942 28577 0 mem_right_track_28.DFFR_1_.Q
rlabel metal1 19918 19346 19918 19346 0 mem_right_track_30.DFFR_0_.Q
rlabel metal2 14122 34000 14122 34000 0 mem_right_track_30.DFFR_1_.Q
rlabel metal1 22678 32912 22678 32912 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 16238 33524 16238 33524 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 25162 31841 25162 31841 0 mem_right_track_34.DFFR_0_.Q
rlabel metal2 13110 34612 13110 34612 0 mem_right_track_34.DFFR_1_.Q
rlabel metal1 19550 25262 19550 25262 0 mem_right_track_36.DFFR_0_.Q
rlabel metal2 18446 19550 18446 19550 0 mem_right_track_4.DFFR_0_.Q
rlabel metal1 4830 32266 4830 32266 0 mem_right_track_4.DFFR_1_.Q
rlabel metal1 6854 29546 6854 29546 0 mem_right_track_6.DFFR_0_.Q
rlabel metal2 8786 27897 8786 27897 0 mem_right_track_6.DFFR_1_.Q
rlabel metal1 13938 19822 13938 19822 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 7958 18020 7958 18020 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 6946 19822 6946 19822 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 14582 28526 14582 28526 0 mem_top_track_10.DFFR_0_.D
rlabel metal1 10948 27642 10948 27642 0 mem_top_track_10.DFFR_0_.Q
rlabel metal1 8740 33422 8740 33422 0 mem_top_track_10.DFFR_1_.Q
rlabel metal1 10350 24786 10350 24786 0 mem_top_track_12.DFFR_0_.Q
rlabel metal1 7130 20400 7130 20400 0 mem_top_track_12.DFFR_1_.Q
rlabel metal1 11776 25262 11776 25262 0 mem_top_track_14.DFFR_0_.Q
rlabel metal1 14030 32198 14030 32198 0 mem_top_track_14.DFFR_1_.Q
rlabel metal1 4324 28526 4324 28526 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 8142 30702 8142 30702 0 mem_top_track_16.DFFR_1_.Q
rlabel metal1 15088 29070 15088 29070 0 mem_top_track_18.DFFR_0_.Q
rlabel metal1 14674 29648 14674 29648 0 mem_top_track_18.DFFR_1_.Q
rlabel metal1 12788 16558 12788 16558 0 mem_top_track_2.DFFR_0_.Q
rlabel metal1 14444 15470 14444 15470 0 mem_top_track_2.DFFR_1_.Q
rlabel metal2 8418 17833 8418 17833 0 mem_top_track_20.DFFR_0_.Q
rlabel metal1 14812 14382 14812 14382 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 13570 21386 13570 21386 0 mem_top_track_22.DFFR_0_.Q
rlabel via2 4554 33405 4554 33405 0 mem_top_track_22.DFFR_1_.Q
rlabel metal1 6900 33626 6900 33626 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 15640 20910 15640 20910 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 18354 32402 18354 32402 0 mem_top_track_26.DFFR_0_.Q
rlabel metal1 7314 36210 7314 36210 0 mem_top_track_26.DFFR_1_.Q
rlabel metal1 14950 25874 14950 25874 0 mem_top_track_28.DFFR_0_.Q
rlabel metal1 10626 28934 10626 28934 0 mem_top_track_28.DFFR_1_.Q
rlabel metal2 12558 36839 12558 36839 0 mem_top_track_30.DFFR_0_.Q
rlabel via2 2346 33541 2346 33541 0 mem_top_track_30.DFFR_1_.Q
rlabel metal1 4646 33626 4646 33626 0 mem_top_track_32.DFFR_0_.Q
rlabel metal2 9568 32878 9568 32878 0 mem_top_track_32.DFFR_1_.Q
rlabel via2 13294 34901 13294 34901 0 mem_top_track_34.DFFR_0_.Q
rlabel metal1 12466 18700 12466 18700 0 mem_top_track_34.DFFR_1_.Q
rlabel metal1 15180 29614 15180 29614 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 14950 20842 14950 20842 0 mem_top_track_4.DFFR_0_.Q
rlabel metal1 9200 29546 9200 29546 0 mem_top_track_4.DFFR_1_.Q
rlabel metal1 12926 24276 12926 24276 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 13202 28186 13202 28186 0 mem_top_track_6.DFFR_1_.Q
rlabel metal1 17526 26350 17526 26350 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 5428 20570 5428 20570 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 13662 18734 13662 18734 0 mux_right_track_0.INVTX1_1_.out
rlabel metal1 11132 8534 11132 8534 0 mux_right_track_0.INVTX1_2_.out
rlabel metal1 10074 21658 10074 21658 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14582 20026 14582 20026 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 9982 24786 9982 24786 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6670 25330 6670 25330 0 mux_right_track_0.out
rlabel metal1 23414 32266 23414 32266 0 mux_right_track_10.INVTX1_0_.out
rlabel metal2 18814 31076 18814 31076 0 mux_right_track_10.INVTX1_1_.out
rlabel metal1 19826 9146 19826 9146 0 mux_right_track_10.INVTX1_2_.out
rlabel metal1 23598 25466 23598 25466 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22678 21794 22678 21794 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23736 21930 23736 21930 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 34086 15470 34086 15470 0 mux_right_track_10.out
rlabel metal1 9614 24038 9614 24038 0 mux_right_track_12.INVTX1_0_.out
rlabel metal1 23322 31824 23322 31824 0 mux_right_track_12.INVTX1_2_.out
rlabel metal1 16606 30158 16606 30158 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18722 29648 18722 29648 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16698 29750 16698 29750 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 15318 32538 15318 32538 0 mux_right_track_12.out
rlabel metal1 25576 8058 25576 8058 0 mux_right_track_14.INVTX1_0_.out
rlabel metal1 28428 11526 28428 11526 0 mux_right_track_14.INVTX1_2_.out
rlabel metal1 19550 28662 19550 28662 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21574 27472 21574 27472 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20010 30022 20010 30022 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16238 35802 16238 35802 0 mux_right_track_14.out
rlabel metal1 27462 32198 27462 32198 0 mux_right_track_16.INVTX1_0_.out
rlabel metal1 12972 22066 12972 22066 0 mux_right_track_16.INVTX1_2_.out
rlabel metal2 24978 25330 24978 25330 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19596 23222 19596 23222 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23782 12818 23782 12818 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 24748 5678 24748 5678 0 mux_right_track_16.out
rlabel metal2 8050 15538 8050 15538 0 mux_right_track_18.INVTX1_0_.out
rlabel metal2 11822 18598 11822 18598 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13386 21454 13386 21454 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11408 10030 11408 10030 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 10258 9894 10258 9894 0 mux_right_track_18.out
rlabel metal2 32614 25126 32614 25126 0 mux_right_track_2.INVTX1_0_.out
rlabel metal1 15134 9146 15134 9146 0 mux_right_track_2.INVTX1_2_.out
rlabel metal1 17020 20026 17020 20026 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16330 18496 16330 18496 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 15226 17408 15226 17408 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 8924 17238 8924 17238 0 mux_right_track_2.out
rlabel metal1 7820 5882 7820 5882 0 mux_right_track_20.INVTX1_0_.out
rlabel metal2 12834 16320 12834 16320 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17802 10642 17802 10642 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19274 10438 19274 10438 0 mux_right_track_20.out
rlabel metal1 25070 5746 25070 5746 0 mux_right_track_22.INVTX1_0_.out
rlabel metal1 17112 15402 17112 15402 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15916 15334 15916 15334 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15732 10438 15732 10438 0 mux_right_track_22.out
rlabel metal2 33718 16320 33718 16320 0 mux_right_track_24.INVTX1_0_.out
rlabel metal1 12328 8602 12328 8602 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 20194 18190 20194 18190 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29486 4114 29486 4114 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 37490 3706 37490 3706 0 mux_right_track_24.out
rlabel metal1 20148 31858 20148 31858 0 mux_right_track_26.INVTX1_0_.out
rlabel metal1 19504 21522 19504 21522 0 mux_right_track_26.INVTX1_1_.out
rlabel metal2 20562 31799 20562 31799 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 4738 5712 4738 5712 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4094 4114 4094 4114 0 mux_right_track_26.out
rlabel metal2 14398 34204 14398 34204 0 mux_right_track_28.INVTX1_0_.out
rlabel metal1 18492 34102 18492 34102 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 21758 26860 21758 26860 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35006 22576 35006 22576 0 mux_right_track_28.out
rlabel metal1 28428 7174 28428 7174 0 mux_right_track_30.INVTX1_0_.out
rlabel metal1 21620 25262 21620 25262 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22770 26520 22770 26520 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23230 29274 23230 29274 0 mux_right_track_30.out
rlabel metal1 24311 32334 24311 32334 0 mux_right_track_32.INVTX1_0_.out
rlabel metal2 22862 32096 22862 32096 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16330 34102 16330 34102 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 15410 35836 15410 35836 0 mux_right_track_32.out
rlabel metal1 30314 33286 30314 33286 0 mux_right_track_34.INVTX1_0_.out
rlabel metal1 25438 30634 25438 30634 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28382 32368 28382 32368 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34132 32470 34132 32470 0 mux_right_track_34.out
rlabel metal1 20470 28594 20470 28594 0 mux_right_track_36.INVTX1_0_.out
rlabel metal1 20976 23834 20976 23834 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18492 23834 18492 23834 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18860 12818 18860 12818 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 18262 5202 18262 5202 0 mux_right_track_36.out
rlabel metal1 27738 12070 27738 12070 0 mux_right_track_4.INVTX1_0_.out
rlabel metal2 22402 17408 22402 17408 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21252 20978 21252 20978 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 22862 25398 22862 25398 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 34454 28662 34454 28662 0 mux_right_track_4.out
rlabel metal1 8096 23630 8096 23630 0 mux_right_track_6.INVTX1_0_.out
rlabel metal1 10764 23766 10764 23766 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18400 25466 18400 25466 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14766 35666 14766 35666 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14720 35802 14720 35802 0 mux_right_track_6.out
rlabel metal1 16859 7718 16859 7718 0 mux_right_track_8.INVTX1_0_.out
rlabel metal2 20286 20162 20286 20162 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21574 21658 21574 21658 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 22540 20910 22540 20910 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 34454 12818 34454 12818 0 mux_right_track_8.out
rlabel metal1 13616 8058 13616 8058 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 14766 17034 14766 17034 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 6394 24718 6394 24718 0 mux_top_track_0.INVTX1_2_.out
rlabel metal1 12857 18122 12857 18122 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10534 19924 10534 19924 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11638 10642 11638 10642 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 11868 10438 11868 10438 0 mux_top_track_0.out
rlabel metal1 18538 27438 18538 27438 0 mux_top_track_10.INVTX1_0_.out
rlabel metal1 12489 25806 12489 25806 0 mux_top_track_10.INVTX1_1_.out
rlabel metal1 16192 32742 16192 32742 0 mux_top_track_10.INVTX1_2_.out
rlabel metal1 14536 26010 14536 26010 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16606 26656 16606 26656 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16882 12206 16882 12206 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17802 12070 17802 12070 0 mux_top_track_10.out
rlabel metal2 8234 29767 8234 29767 0 mux_top_track_12.INVTX1_1_.out
rlabel metal2 19274 15572 19274 15572 0 mux_top_track_12.INVTX1_2_.out
rlabel metal1 11684 20502 11684 20502 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16284 16966 16284 16966 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 5658 8466 5658 8466 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 3956 3026 3956 3026 0 mux_top_track_12.out
rlabel metal2 22402 10200 22402 10200 0 mux_top_track_14.INVTX1_1_.out
rlabel metal1 7222 23154 7222 23154 0 mux_top_track_14.INVTX1_2_.out
rlabel metal1 14030 23222 14030 23222 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12374 22542 12374 22542 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 20010 11118 20010 11118 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 20378 11050 20378 11050 0 mux_top_track_14.out
rlabel metal2 5566 26996 5566 26996 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 8648 27574 8648 27574 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13938 32470 13938 32470 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 14030 32708 14030 32708 0 mux_top_track_16.out
rlabel metal1 9430 15130 9430 15130 0 mux_top_track_18.INVTX1_1_.out
rlabel metal2 32430 30158 32430 30158 0 mux_top_track_18.INVTX1_2_.out
rlabel metal1 13616 17782 13616 17782 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20838 29002 20838 29002 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17572 27846 17572 27846 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17664 35054 17664 35054 0 mux_top_track_18.out
rlabel metal2 16974 19482 16974 19482 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 10856 6358 10856 6358 0 mux_top_track_2.INVTX1_2_.out
rlabel metal2 16514 18530 16514 18530 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15134 16320 15134 16320 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16974 16626 16974 16626 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 24656 10438 24656 10438 0 mux_top_track_2.out
rlabel metal2 7038 16116 7038 16116 0 mux_top_track_20.INVTX1_1_.out
rlabel metal2 8970 17340 8970 17340 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24127 10710 24127 10710 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30038 4590 30038 4590 0 mux_top_track_20.out
rlabel metal1 23230 5644 23230 5644 0 mux_top_track_22.INVTX1_1_.out
rlabel metal2 22770 19924 22770 19924 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 24518 19822 24518 19822 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30314 19040 30314 19040 0 mux_top_track_22.out
rlabel metal1 17940 21522 17940 21522 0 mux_top_track_24.INVTX1_0_.out
rlabel metal1 8234 26418 8234 26418 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 16054 22066 16054 22066 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19458 20264 19458 20264 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34822 14382 34822 14382 0 mux_top_track_24.out
rlabel metal2 18262 30736 18262 30736 0 mux_top_track_26.INVTX1_0_.out
rlabel metal2 31786 32096 31786 32096 0 mux_top_track_26.INVTX1_1_.out
rlabel metal1 18952 30634 18952 30634 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13478 19499 13478 19499 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4830 10030 4830 10030 0 mux_top_track_26.out
rlabel metal1 23138 6970 23138 6970 0 mux_top_track_28.INVTX1_1_.out
rlabel metal1 19596 22134 19596 22134 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12328 26826 12328 26826 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 6670 24990 6670 24990 0 mux_top_track_28.out
rlabel metal1 7268 19958 7268 19958 0 mux_top_track_30.INVTX1_1_.out
rlabel metal1 9062 19686 9062 19686 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 35052 7854 35052 7854 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 37122 6698 37122 6698 0 mux_top_track_30.out
rlabel metal1 2990 27098 2990 27098 0 mux_top_track_32.INVTX1_1_.out
rlabel metal1 5382 29036 5382 29036 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9660 29478 9660 29478 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12006 31110 12006 31110 0 mux_top_track_32.out
rlabel metal1 12052 17102 12052 17102 0 mux_top_track_34.INVTX1_1_.out
rlabel metal2 14030 17714 14030 17714 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20194 18496 20194 18496 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33580 16082 33580 16082 0 mux_top_track_34.out
rlabel metal1 19504 31858 19504 31858 0 mux_top_track_36.INVTX1_1_.out
rlabel metal2 19550 26418 19550 26418 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 21482 26112 21482 26112 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 31096 25874 31096 25874 0 mux_top_track_36.out
rlabel metal2 6762 21726 6762 21726 0 mux_top_track_4.INVTX1_2_.out
rlabel metal1 18216 21658 18216 21658 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16790 21114 16790 21114 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17894 23154 17894 23154 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 34822 26350 34822 26350 0 mux_top_track_4.out
rlabel metal1 6946 20026 6946 20026 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 14168 24582 14168 24582 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 10626 21964 10626 21964 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13570 29716 13570 29716 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 13662 34034 13662 34034 0 mux_top_track_6.out
rlabel metal2 31786 27064 31786 27064 0 mux_top_track_8.INVTX1_2_.out
rlabel metal1 17526 27370 17526 27370 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20010 26282 20010 26282 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15042 26826 15042 26826 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 9384 25806 9384 25806 0 mux_top_track_8.out
rlabel metal2 37306 6137 37306 6137 0 net1
rlabel metal1 2116 23290 2116 23290 0 net10
rlabel metal1 8648 20978 8648 20978 0 net100
rlabel metal1 14536 14042 14536 14042 0 net101
rlabel metal1 14996 22746 14996 22746 0 net102
rlabel metal2 7774 22814 7774 22814 0 net103
rlabel metal1 20056 25874 20056 25874 0 net104
rlabel metal1 14674 24922 14674 24922 0 net105
rlabel metal1 19182 16150 19182 16150 0 net106
rlabel metal2 9522 22338 9522 22338 0 net107
rlabel metal2 20286 26112 20286 26112 0 net108
rlabel metal2 13662 19992 13662 19992 0 net109
rlabel metal1 10810 2618 10810 2618 0 net11
rlabel metal1 14444 16558 14444 16558 0 net110
rlabel metal1 20378 19482 20378 19482 0 net111
rlabel metal2 18538 26384 18538 26384 0 net112
rlabel metal1 21436 20570 21436 20570 0 net113
rlabel metal1 22080 21522 22080 21522 0 net114
rlabel metal2 21298 28458 21298 28458 0 net115
rlabel metal1 23322 23732 23322 23732 0 net116
rlabel metal1 20056 23086 20056 23086 0 net117
rlabel metal2 13110 21216 13110 21216 0 net118
rlabel metal2 17802 23868 17802 23868 0 net119
rlabel metal3 16997 33116 16997 33116 0 net12
rlabel metal2 13478 30345 13478 30345 0 net120
rlabel metal2 18998 16660 18998 16660 0 net121
rlabel metal1 23920 19482 23920 19482 0 net122
rlabel metal1 18216 20366 18216 20366 0 net123
rlabel metal2 13110 20706 13110 20706 0 net124
rlabel metal2 10534 29614 10534 29614 0 net125
rlabel metal1 16790 17306 16790 17306 0 net126
rlabel metal2 7958 30668 7958 30668 0 net127
rlabel metal2 18630 18530 18630 18530 0 net128
rlabel metal2 20838 26078 20838 26078 0 net129
rlabel metal1 4692 2550 4692 2550 0 net13
rlabel metal1 13064 15538 13064 15538 0 net130
rlabel metal2 15962 14790 15962 14790 0 net131
rlabel metal2 22126 17952 22126 17952 0 net132
rlabel metal2 13202 19618 13202 19618 0 net133
rlabel metal1 22954 25806 22954 25806 0 net134
rlabel metal1 22954 27438 22954 27438 0 net135
rlabel metal1 16560 33626 16560 33626 0 net136
rlabel metal1 25668 31790 25668 31790 0 net137
rlabel metal2 1610 21556 1610 21556 0 net14
rlabel metal2 5842 19108 5842 19108 0 net15
rlabel metal2 35466 28220 35466 28220 0 net16
rlabel metal1 16238 32844 16238 32844 0 net17
rlabel metal1 31970 2550 31970 2550 0 net18
rlabel metal1 3818 24616 3818 24616 0 net19
rlabel metal1 22678 37128 22678 37128 0 net2
rlabel metal2 13846 27761 13846 27761 0 net20
rlabel metal2 37030 28492 37030 28492 0 net21
rlabel metal2 34546 4692 34546 4692 0 net22
rlabel metal1 34730 16626 34730 16626 0 net23
rlabel metal1 27278 32878 27278 32878 0 net24
rlabel metal1 14214 34544 14214 34544 0 net25
rlabel metal1 36294 3162 36294 3162 0 net26
rlabel metal1 37007 32538 37007 32538 0 net27
rlabel metal1 36317 37094 36317 37094 0 net28
rlabel metal1 20286 33490 20286 33490 0 net29
rlabel metal1 37122 36006 37122 36006 0 net3
rlabel metal2 1610 19958 1610 19958 0 net30
rlabel metal2 38134 10132 38134 10132 0 net31
rlabel metal2 6762 23222 6762 23222 0 net32
rlabel metal1 4968 3706 4968 3706 0 net33
rlabel metal1 24932 37162 24932 37162 0 net34
rlabel metal1 3404 32742 3404 32742 0 net35
rlabel metal1 29532 2618 29532 2618 0 net36
rlabel metal1 33028 37094 33028 37094 0 net37
rlabel metal1 4784 10234 4784 10234 0 net38
rlabel metal1 4554 2618 4554 2618 0 net39
rlabel metal2 6946 13974 6946 13974 0 net4
rlabel metal2 1886 5321 1886 5321 0 net40
rlabel metal1 6739 2278 6739 2278 0 net41
rlabel metal2 2346 5780 2346 5780 0 net42
rlabel metal1 34730 37094 34730 37094 0 net43
rlabel metal2 27830 36992 27830 36992 0 net44
rlabel metal2 18170 5780 18170 5780 0 net45
rlabel metal1 36754 36550 36754 36550 0 net46
rlabel metal1 38042 4794 38042 4794 0 net47
rlabel metal2 19458 33932 19458 33932 0 net48
rlabel metal1 37007 21862 37007 21862 0 net49
rlabel metal1 33764 2618 33764 2618 0 net5
rlabel metal1 8372 2618 8372 2618 0 net50
rlabel metal1 13892 7854 13892 7854 0 net51
rlabel metal2 8878 15334 8878 15334 0 net52
rlabel metal2 38134 23358 38134 23358 0 net53
rlabel metal1 20654 8466 20654 8466 0 net54
rlabel metal1 31510 37094 31510 37094 0 net55
rlabel metal1 27830 29138 27830 29138 0 net56
rlabel metal1 16376 36006 16376 36006 0 net57
rlabel metal1 10212 31790 10212 31790 0 net58
rlabel metal1 23644 8466 23644 8466 0 net59
rlabel metal1 18400 36006 18400 36006 0 net6
rlabel metal1 4600 11322 4600 11322 0 net60
rlabel metal1 37996 33490 37996 33490 0 net61
rlabel metal1 1794 26962 1794 26962 0 net62
rlabel metal2 22678 3706 22678 3706 0 net63
rlabel metal2 14950 3706 14950 3706 0 net64
rlabel metal2 38042 2890 38042 2890 0 net65
rlabel metal1 1610 2448 1610 2448 0 net66
rlabel metal2 38042 21658 38042 21658 0 net67
rlabel metal1 23690 35258 23690 35258 0 net68
rlabel metal1 15180 35802 15180 35802 0 net69
rlabel metal1 37030 36618 37030 36618 0 net7
rlabel metal1 37674 37230 37674 37230 0 net70
rlabel metal2 16882 3706 16882 3706 0 net71
rlabel metal2 5750 17068 5750 17068 0 net72
rlabel metal2 34270 32572 34270 32572 0 net73
rlabel metal2 15778 36788 15778 36788 0 net74
rlabel metal2 35374 10778 35374 10778 0 net75
rlabel metal2 38042 14076 38042 14076 0 net76
rlabel metal1 15686 36278 15686 36278 0 net77
rlabel metal1 13478 35530 13478 35530 0 net78
rlabel metal2 25898 3978 25898 3978 0 net79
rlabel metal2 25438 4624 25438 4624 0 net8
rlabel metal2 9154 3978 9154 3978 0 net80
rlabel metal2 11730 3706 11730 3706 0 net81
rlabel metal1 36041 2414 36041 2414 0 net82
rlabel metal2 38042 17884 38042 17884 0 net83
rlabel metal2 37306 12682 37306 12682 0 net84
rlabel metal1 2806 6290 2806 6290 0 net85
rlabel metal1 1564 32878 1564 32878 0 net86
rlabel metal1 37950 3026 37950 3026 0 net87
rlabel metal1 6900 34578 6900 34578 0 net88
rlabel metal2 35374 15130 35374 15130 0 net89
rlabel metal1 4002 8058 4002 8058 0 net9
rlabel metal2 38042 25466 38042 25466 0 net90
rlabel metal1 32016 2414 32016 2414 0 net91
rlabel metal2 38042 26996 38042 26996 0 net92
rlabel metal2 12650 35853 12650 35853 0 net93
rlabel metal1 1610 24208 1610 24208 0 net94
rlabel metal2 19458 3978 19458 3978 0 net95
rlabel metal1 1610 3060 1610 3060 0 net96
rlabel metal1 23920 2414 23920 2414 0 net97
rlabel metal1 12926 32776 12926 32776 0 net98
rlabel metal1 18768 35190 18768 35190 0 net99
rlabel metal3 1188 4828 1188 4828 0 pReset
rlabel metal1 2070 25330 2070 25330 0 prog_clk
rlabel metal2 5842 1588 5842 1588 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 1334 1860 1334 1860 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 34960 37230 34960 37230 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 27876 37230 27876 37230 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 18078 1588 18078 1588 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 37674 36788 37674 36788 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 38318 4369 38318 4369 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 1334 37529 1334 37529 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 38318 21913 38318 21913 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 7130 1588 7130 1588 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 13570 1588 13570 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1234 14348 1234 14348 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 38318 24021 38318 24021 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 32384 37230 32384 37230 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 30498 37230 30498 37230 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 14490 35496 14490 35496 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 10350 34544 10350 34544 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 27094 1588 27094 1588 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal3 1234 10948 1234 10948 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
