// This is the unpowered netlist.
module cbx_1__1_ (bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_,
    top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_,
    vccd1,
    vssd1,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out);
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
 inout vccd1;
 inout vssd1;
 input [0:18] chanx_left_in;
 output [0:18] chanx_left_out;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire \mem_bottom_ipin_0.DFFR_0_.Q ;
 wire \mem_bottom_ipin_0.DFFR_1_.Q ;
 wire \mem_bottom_ipin_0.DFFR_2_.Q ;
 wire \mem_bottom_ipin_0.DFFR_3_.Q ;
 wire \mem_bottom_ipin_0.DFFR_4_.Q ;
 wire \mem_bottom_ipin_0.DFFR_5_.Q ;
 wire \mem_bottom_ipin_1.DFFR_0_.Q ;
 wire \mem_bottom_ipin_1.DFFR_1_.Q ;
 wire \mem_bottom_ipin_1.DFFR_2_.Q ;
 wire \mem_bottom_ipin_1.DFFR_3_.Q ;
 wire \mem_bottom_ipin_1.DFFR_4_.Q ;
 wire \mem_bottom_ipin_1.DFFR_5_.Q ;
 wire \mem_bottom_ipin_2.DFFR_0_.Q ;
 wire \mem_bottom_ipin_2.DFFR_1_.Q ;
 wire \mem_bottom_ipin_2.DFFR_2_.Q ;
 wire \mem_bottom_ipin_2.DFFR_3_.Q ;
 wire \mem_bottom_ipin_2.DFFR_4_.Q ;
 wire \mem_bottom_ipin_2.DFFR_5_.Q ;
 wire \mem_top_ipin_0.DFFR_0_.Q ;
 wire \mem_top_ipin_0.DFFR_1_.Q ;
 wire \mem_top_ipin_0.DFFR_2_.Q ;
 wire \mem_top_ipin_0.DFFR_3_.Q ;
 wire \mem_top_ipin_0.DFFR_4_.Q ;
 wire \mem_top_ipin_0.DFFR_5_.Q ;
 wire \mem_top_ipin_1.DFFR_0_.Q ;
 wire \mem_top_ipin_1.DFFR_1_.Q ;
 wire \mem_top_ipin_1.DFFR_2_.Q ;
 wire \mem_top_ipin_1.DFFR_3_.Q ;
 wire \mem_top_ipin_1.DFFR_4_.Q ;
 wire \mem_top_ipin_1.DFFR_5_.Q ;
 wire \mem_top_ipin_2.DFFR_0_.Q ;
 wire \mem_top_ipin_2.DFFR_1_.Q ;
 wire \mem_top_ipin_2.DFFR_2_.Q ;
 wire \mem_top_ipin_2.DFFR_3_.Q ;
 wire \mem_top_ipin_2.DFFR_4_.Q ;
 wire \mem_top_ipin_2.DFFR_5_.Q ;
 wire \mem_top_ipin_3.DFFR_0_.Q ;
 wire \mem_top_ipin_3.DFFR_1_.Q ;
 wire \mem_top_ipin_3.DFFR_2_.Q ;
 wire \mem_top_ipin_3.DFFR_3_.Q ;
 wire \mem_top_ipin_3.DFFR_4_.Q ;
 wire \mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \mux_bottom_ipin_0.INVTX1_2_.out ;
 wire \mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \mux_bottom_ipin_0.INVTX1_4_.out ;
 wire \mux_bottom_ipin_0.INVTX1_5_.out ;
 wire \mux_bottom_ipin_0.INVTX1_6_.out ;
 wire \mux_bottom_ipin_0.INVTX1_7_.out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_1.INVTX1_2_.out ;
 wire \mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \mux_bottom_ipin_1.INVTX1_4_.out ;
 wire \mux_bottom_ipin_1.INVTX1_5_.out ;
 wire \mux_bottom_ipin_1.INVTX1_6_.out ;
 wire \mux_bottom_ipin_1.INVTX1_7_.out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_0.INVTX1_2_.out ;
 wire \mux_top_ipin_0.INVTX1_3_.out ;
 wire \mux_top_ipin_0.INVTX1_4_.out ;
 wire \mux_top_ipin_0.INVTX1_5_.out ;
 wire \mux_top_ipin_0.INVTX1_6_.out ;
 wire \mux_top_ipin_0.INVTX1_7_.out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_1.INVTX1_2_.out ;
 wire \mux_top_ipin_1.INVTX1_3_.out ;
 wire \mux_top_ipin_1.INVTX1_4_.out ;
 wire \mux_top_ipin_1.INVTX1_5_.out ;
 wire \mux_top_ipin_1.INVTX1_6_.out ;
 wire \mux_top_ipin_1.INVTX1_7_.out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_2.INVTX1_2_.out ;
 wire \mux_top_ipin_2.INVTX1_3_.out ;
 wire \mux_top_ipin_2.INVTX1_6_.out ;
 wire \mux_top_ipin_2.INVTX1_7_.out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;

 sky130_fd_sc_hd__inv_2 _134_ (.A(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _136_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _137_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _138_ (.A(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _139_ (.A(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _140_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _141_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _142_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _143_ (.A(\mem_top_ipin_3.DFFR_3_.Q ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _146_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(net45),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _148_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _149_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _150_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _151_ (.A(\mem_top_ipin_3.DFFR_4_.Q ),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _152_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _153_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _154_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _155_ (.A(\mem_top_ipin_2.DFFR_3_.Q ),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _156_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _157_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _158_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _159_ (.A(\mem_top_ipin_2.DFFR_5_.Q ),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(\mem_top_ipin_2.DFFR_4_.Q ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(\mem_top_ipin_1.DFFR_3_.Q ),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _170_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(\mem_top_ipin_1.DFFR_5_.Q ),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(\mem_top_ipin_1.DFFR_4_.Q ),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(\mem_top_ipin_0.DFFR_3_.Q ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _181_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(\mem_top_ipin_0.DFFR_5_.Q ),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(\mem_top_ipin_0.DFFR_4_.Q ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _193_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _194_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _195_ (.A(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _196_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _197_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _202_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _210_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _211_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _212_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _213_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _215_ (.A(net24),
    .Y(\mux_bottom_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _216_ (.A(net11),
    .Y(\mux_bottom_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _217_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _218_ (.A(net30),
    .Y(\mux_bottom_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _219_ (.A(net2),
    .Y(\mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _220_ (.A(net21),
    .Y(\mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _221_ (.A(net17),
    .Y(\mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _222_ (.A(net36),
    .Y(\mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _223_ (.A(net5),
    .Y(\mux_bottom_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _224_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _225_ (.A(net6),
    .Y(\mux_bottom_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _226_ (.A(net37),
    .Y(\mux_bottom_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _227_ (.A(net18),
    .Y(\mux_bottom_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _228_ (.A(net31),
    .Y(\mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _229_ (.A(net12),
    .Y(\mux_bottom_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _230_ (.A(net25),
    .Y(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _231_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net41));
 sky130_fd_sc_hd__clkinv_2 _232_ (.A(net8),
    .Y(\mux_top_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _233_ (.A(net39),
    .Y(\mux_top_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _234_ (.A(net20),
    .Y(\mux_top_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _235_ (.A(net33),
    .Y(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net14),
    .Y(\mux_top_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _237_ (.A(net27),
    .Y(\mux_top_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _238_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _239_ (.A(net9),
    .Y(\mux_top_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net22),
    .Y(\mux_top_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _241_ (.A(net3),
    .Y(\mux_top_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _242_ (.A(net34),
    .Y(\mux_top_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _243_ (.A(net15),
    .Y(\mux_top_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _244_ (.A(net28),
    .Y(\mux_top_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _245_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _246_ (.A(net10),
    .Y(\mux_top_ipin_2.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _247_ (.A(net35),
    .Y(\mux_top_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _248_ (.A(net16),
    .Y(\mux_top_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _249_ (.A(net29),
    .Y(\mux_top_ipin_2.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _250_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _251_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _252_ (.A(net4),
    .Y(\mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _253_ (.A(net32),
    .Y(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _254_ (.A(net13),
    .Y(\mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _255_ (.A(net23),
    .Y(\mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__buf_4 _256_ (.A(net40),
    .X(_042_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(_042_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(_042_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(_042_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(_042_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(_042_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(_042_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(_042_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(_042_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(_042_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(_042_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_4 _267_ (.A(net40),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(_043_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(_043_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _270_ (.A(_043_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _271_ (.A(_043_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _272_ (.A(_043_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _273_ (.A(_043_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _274_ (.A(_043_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _275_ (.A(_043_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _276_ (.A(_043_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _277_ (.A(_043_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _278_ (.A(net40),
    .X(_044_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(_044_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(_044_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(_044_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(_044_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(_044_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(_044_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(_044_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _286_ (.A(_044_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(_044_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(_044_),
    .Y(_029_));
 sky130_fd_sc_hd__buf_4 _289_ (.A(net40),
    .X(_045_));
 sky130_fd_sc_hd__inv_2 _290_ (.A(_045_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(_045_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _292_ (.A(_045_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(_045_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(_045_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(_045_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(_045_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _297_ (.A(_045_),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(_045_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(_045_),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(net40),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(net40),
    .Y(_041_));
 sky130_fd_sc_hd__dfrtp_1 _302_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .RESET_B(_000_),
    .Q(\mem_bottom_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _303_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .RESET_B(_001_),
    .Q(\mem_bottom_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _304_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .RESET_B(_002_),
    .Q(\mem_bottom_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _305_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .RESET_B(_003_),
    .Q(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _306_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .RESET_B(_004_),
    .Q(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _307_ (.CLK(prog_clk),
    .D(net1),
    .RESET_B(_005_),
    .Q(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _308_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .RESET_B(_006_),
    .Q(\mem_bottom_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _309_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .RESET_B(_007_),
    .Q(\mem_bottom_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _310_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .RESET_B(_008_),
    .Q(\mem_bottom_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _311_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .RESET_B(_009_),
    .Q(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _312_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .RESET_B(_010_),
    .Q(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _313_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .RESET_B(_011_),
    .Q(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _314_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_4_.Q ),
    .RESET_B(_012_),
    .Q(\mem_top_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _315_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_3_.Q ),
    .RESET_B(_013_),
    .Q(\mem_top_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _316_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_2_.Q ),
    .RESET_B(_014_),
    .Q(\mem_top_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _317_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_1_.Q ),
    .RESET_B(_015_),
    .Q(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _318_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_0_.Q ),
    .RESET_B(_016_),
    .Q(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _319_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .RESET_B(_017_),
    .Q(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _320_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_4_.Q ),
    .RESET_B(_018_),
    .Q(\mem_top_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _321_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_3_.Q ),
    .RESET_B(_019_),
    .Q(\mem_top_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _322_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_2_.Q ),
    .RESET_B(_020_),
    .Q(\mem_top_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _323_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_1_.Q ),
    .RESET_B(_021_),
    .Q(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _324_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_0_.Q ),
    .RESET_B(_022_),
    .Q(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _325_ (.CLK(prog_clk),
    .D(\mem_top_ipin_0.DFFR_5_.Q ),
    .RESET_B(_023_),
    .Q(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _326_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_4_.Q ),
    .RESET_B(_024_),
    .Q(\mem_top_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _327_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_3_.Q ),
    .RESET_B(_025_),
    .Q(\mem_top_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _328_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_2_.Q ),
    .RESET_B(_026_),
    .Q(\mem_top_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _329_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_1_.Q ),
    .RESET_B(_027_),
    .Q(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _330_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_0_.Q ),
    .RESET_B(_028_),
    .Q(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _331_ (.CLK(prog_clk),
    .D(\mem_top_ipin_1.DFFR_5_.Q ),
    .RESET_B(_029_),
    .Q(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _332_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_4_.Q ),
    .RESET_B(_030_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _333_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_3_.Q ),
    .RESET_B(_031_),
    .Q(\mem_top_ipin_3.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _334_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_2_.Q ),
    .RESET_B(_032_),
    .Q(\mem_top_ipin_3.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _335_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_1_.Q ),
    .RESET_B(_033_),
    .Q(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _336_ (.CLK(prog_clk),
    .D(\mem_top_ipin_3.DFFR_0_.Q ),
    .RESET_B(_034_),
    .Q(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _337_ (.CLK(prog_clk),
    .D(\mem_top_ipin_2.DFFR_5_.Q ),
    .RESET_B(_035_),
    .Q(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _338_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .RESET_B(_036_),
    .Q(\mem_bottom_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _339_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .RESET_B(_037_),
    .Q(\mem_bottom_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _340_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .RESET_B(_038_),
    .Q(\mem_bottom_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _341_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .RESET_B(_039_),
    .Q(\mem_bottom_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _342_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .RESET_B(_040_),
    .Q(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _343_ (.CLK(prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .RESET_B(_041_),
    .Q(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _402__88 (.HI(net88));
 sky130_fd_sc_hd__conb_1 _416__89 (.HI(net89));
 sky130_fd_sc_hd__conb_1 _428__90 (.HI(net90));
 sky130_fd_sc_hd__conb_1 _440__91 (.HI(net91));
 sky130_fd_sc_hd__conb_1 _452__92 (.HI(net92));
 sky130_fd_sc_hd__conb_1 _462__93 (.HI(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__clkbuf_1 _351_ (.A(net30),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _352_ (.A(net29),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _353_ (.A(net28),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _354_ (.A(net27),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _355_ (.A(net26),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _356_ (.A(net25),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _357_ (.A(net24),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _358_ (.A(net23),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _359_ (.A(net22),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 _360_ (.A(net39),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _361_ (.A(net38),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(net37),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _363_ (.A(net36),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _364_ (.A(net35),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _365_ (.A(net34),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _366_ (.A(net33),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _367_ (.A(net32),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _368_ (.A(net31),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _369_ (.A(net21),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(net11),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 _371_ (.A(net10),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(net9),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 _373_ (.A(net8),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _374_ (.A(net7),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(net6),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _376_ (.A(net5),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _377_ (.A(net4),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _378_ (.A(net3),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(net20),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _380_ (.A(net19),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(net18),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _382_ (.A(net17),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _383_ (.A(net16),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _384_ (.A(net15),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(net14),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _386_ (.A(net13),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 _387_ (.A(net12),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(net2),
    .X(net65));
 sky130_fd_sc_hd__ebufn_2 _389_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_046_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _390_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_047_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _391_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_048_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _392_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_049_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _393_ (.A(net87),
    .TE_B(_050_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _394_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_051_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _395_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_052_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _396_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_053_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _397_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_054_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _398_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_055_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _399_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_056_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _400_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_057_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _401_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_058_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _402_ (.A(net88),
    .TE_B(_059_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _403_ (.A(\mux_bottom_ipin_1.INVTX1_7_.out ),
    .TE_B(_060_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _404_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_061_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _405_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_062_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _406_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_063_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _407_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_064_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _408_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_065_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _409_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_066_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _410_ (.A(\mux_bottom_ipin_1.INVTX1_6_.out ),
    .TE_B(_067_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _411_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_068_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _412_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_069_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _413_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_070_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _414_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_071_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _415_ (.A(\mux_top_ipin_0.INVTX1_7_.out ),
    .TE_B(_072_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _416_ (.A(net89),
    .TE_B(_073_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _417_ (.A(\mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_074_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _418_ (.A(\mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_075_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _419_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_076_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _420_ (.A(\mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_077_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _421_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_078_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _422_ (.A(\mux_top_ipin_0.INVTX1_6_.out ),
    .TE_B(_079_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _423_ (.A(\mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_080_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _424_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_081_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _425_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_082_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _426_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_083_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _427_ (.A(\mux_top_ipin_1.INVTX1_7_.out ),
    .TE_B(_084_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _428_ (.A(net90),
    .TE_B(_085_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _429_ (.A(\mux_top_ipin_1.INVTX1_4_.out ),
    .TE_B(_086_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _430_ (.A(\mux_top_ipin_1.INVTX1_5_.out ),
    .TE_B(_087_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _431_ (.A(\mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_088_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _432_ (.A(\mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_089_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _433_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_090_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _434_ (.A(\mux_top_ipin_1.INVTX1_6_.out ),
    .TE_B(_091_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _435_ (.A(\mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_092_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _436_ (.A(\mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_093_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _437_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_094_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _438_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_095_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _439_ (.A(\mux_top_ipin_2.INVTX1_7_.out ),
    .TE_B(_096_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _440_ (.A(net91),
    .TE_B(_097_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _441_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_098_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _442_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_099_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _443_ (.A(\mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_100_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _444_ (.A(\mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_101_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _445_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_102_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _446_ (.A(\mux_top_ipin_2.INVTX1_6_.out ),
    .TE_B(_103_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _447_ (.A(\mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_104_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _448_ (.A(\mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_105_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _449_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_106_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _450_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_107_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _451_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_108_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _452_ (.A(net92),
    .TE_B(_109_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _453_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_110_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _454_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_111_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _455_ (.A(\mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_112_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _456_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_113_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _457_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_114_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _458_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_115_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _459_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_116_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _460_ (.A(\mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_117_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _461_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_118_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _462_ (.A(net93),
    .TE_B(_119_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _463_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_120_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _464_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_121_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _465_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_122_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _466_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_123_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _467_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_124_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _468_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_125_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _469_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_126_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(ccff_head),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(chanx_left_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(chanx_left_in[10]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(chanx_left_in[11]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(chanx_left_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(chanx_left_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(chanx_left_in[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(chanx_left_in[15]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(chanx_left_in[16]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(chanx_left_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(chanx_left_in[18]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(chanx_left_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(chanx_left_in[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(chanx_left_in[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(chanx_left_in[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(chanx_left_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chanx_left_in[6]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(chanx_left_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(chanx_left_in[8]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(chanx_left_in[9]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(chanx_right_in[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(chanx_right_in[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(chanx_right_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chanx_right_in[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chanx_right_in[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chanx_right_in[14]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(chanx_right_in[15]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(chanx_right_in[16]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(chanx_right_in[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chanx_right_in[18]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(chanx_right_in[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chanx_right_in[2]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(chanx_right_in[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(chanx_right_in[4]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(chanx_right_in[5]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(chanx_right_in[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chanx_right_in[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(chanx_right_in[8]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(chanx_right_in[9]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(pReset),
    .X(net40));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_));
 sky130_fd_sc_hd__conb_1 _393__87 (.HI(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(chanx_left_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(chanx_left_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(chanx_left_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(chanx_left_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(chanx_left_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(chanx_left_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(chanx_left_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(chanx_left_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(chanx_left_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(chanx_left_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chanx_left_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chanx_left_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chanx_left_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chanx_left_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chanx_left_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chanx_left_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chanx_left_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chanx_left_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chanx_left_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chanx_right_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chanx_right_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chanx_right_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chanx_right_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chanx_right_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chanx_right_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chanx_right_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chanx_right_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chanx_right_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chanx_right_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chanx_right_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chanx_right_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chanx_right_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chanx_right_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chanx_right_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chanx_right_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chanx_right_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chanx_right_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chanx_right_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__304__D (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__D (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__D (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A (.DIODE(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__310__D (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__341__D (.DIODE(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__A (.DIODE(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__A (.DIODE(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__318__D (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A (.DIODE(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__317__D (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A (.DIODE(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__316__D (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__329__D (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__328__D (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__334__D (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__A (.DIODE(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__A (.DIODE(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__403__A (.DIODE(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__423__A (.DIODE(\mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__A (.DIODE(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A (.DIODE(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__250__A (.DIODE(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(pReset));
 sky130_fd_sc_hd__diode_2 ANTENNA__343__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__342__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__341__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__340__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__339__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__337__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__336__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__335__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__334__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__333__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__332__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__331__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__330__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__329__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__328__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__327__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__326__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__325__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__324__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__323__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__322__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__321__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__320__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__319__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__318__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__317__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__316__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__315__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__314__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__313__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__310__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__309__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__308__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__307__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__306__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__305__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__304__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__303__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__302__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__307__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__374__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__373__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__232__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__372__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__386__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__385__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__383__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__382__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__221__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__381__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__380__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__369__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__359__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__358__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__357__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__355__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__354__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__353__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__352__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__365__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__363__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__360__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__301__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__147__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_378 ();
endmodule

