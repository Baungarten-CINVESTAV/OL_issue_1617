magic
tech sky130A
magscale 1 2
timestamp 1674174375
<< viali >>
rect 2973 37417 3007 37451
rect 13645 37417 13679 37451
rect 14473 37417 14507 37451
rect 35081 37417 35115 37451
rect 36737 37417 36771 37451
rect 2329 37349 2363 37383
rect 6745 37281 6779 37315
rect 20637 37281 20671 37315
rect 22753 37281 22787 37315
rect 2145 37213 2179 37247
rect 2881 37213 2915 37247
rect 4261 37213 4295 37247
rect 5273 37213 5307 37247
rect 7297 37213 7331 37247
rect 9413 37213 9447 37247
rect 10701 37213 10735 37247
rect 12633 37213 12667 37247
rect 14381 37213 14415 37247
rect 15853 37213 15887 37247
rect 17141 37213 17175 37247
rect 17601 37213 17635 37247
rect 19441 37213 19475 37247
rect 20913 37213 20947 37247
rect 22017 37213 22051 37247
rect 24593 37213 24627 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 29745 37213 29779 37247
rect 30757 37213 30791 37247
rect 32321 37213 32355 37247
rect 33609 37213 33643 37247
rect 35725 37213 35759 37247
rect 36921 37213 36955 37247
rect 37473 37213 37507 37247
rect 35541 37145 35575 37179
rect 4077 37077 4111 37111
rect 5457 37077 5491 37111
rect 7389 37077 7423 37111
rect 9229 37077 9263 37111
rect 10517 37077 10551 37111
rect 12449 37077 12483 37111
rect 15669 37077 15703 37111
rect 16957 37077 16991 37111
rect 19625 37077 19659 37111
rect 22201 37077 22235 37111
rect 24777 37077 24811 37111
rect 25513 37077 25547 37111
rect 27353 37077 27387 37111
rect 29929 37077 29963 37111
rect 30573 37077 30607 37111
rect 32505 37077 32539 37111
rect 33793 37077 33827 37111
rect 37657 37077 37691 37111
rect 2697 36873 2731 36907
rect 13553 36873 13587 36907
rect 15117 36873 15151 36907
rect 20545 36873 20579 36907
rect 21281 36873 21315 36907
rect 22661 36805 22695 36839
rect 37565 36805 37599 36839
rect 38209 36805 38243 36839
rect 1685 36737 1719 36771
rect 3157 36737 3191 36771
rect 13737 36737 13771 36771
rect 15301 36737 15335 36771
rect 21097 36737 21131 36771
rect 22017 36737 22051 36771
rect 27169 36737 27203 36771
rect 27813 36737 27847 36771
rect 14289 36669 14323 36703
rect 25237 36669 25271 36703
rect 22201 36601 22235 36635
rect 27353 36601 27387 36635
rect 38025 36601 38059 36635
rect 1777 36533 1811 36567
rect 1685 36329 1719 36363
rect 38209 36329 38243 36363
rect 2329 36261 2363 36295
rect 1869 36125 1903 36159
rect 37565 36125 37599 36159
rect 38025 36125 38059 36159
rect 38025 35649 38059 35683
rect 37473 35445 37507 35479
rect 38209 35445 38243 35479
rect 18429 34153 18463 34187
rect 18245 33949 18279 33983
rect 17693 33813 17727 33847
rect 1685 33473 1719 33507
rect 37565 33473 37599 33507
rect 38209 33473 38243 33507
rect 1869 33337 1903 33371
rect 38025 33337 38059 33371
rect 1685 33065 1719 33099
rect 5181 33065 5215 33099
rect 4997 32861 5031 32895
rect 9873 32861 9907 32895
rect 5733 32725 5767 32759
rect 9689 32725 9723 32759
rect 10425 32725 10459 32759
rect 22201 32385 22235 32419
rect 38025 32385 38059 32419
rect 22017 32181 22051 32215
rect 22753 32181 22787 32215
rect 38209 32181 38243 32215
rect 9873 31977 9907 32011
rect 1777 31909 1811 31943
rect 1593 31773 1627 31807
rect 9965 31773 9999 31807
rect 10517 31773 10551 31807
rect 1593 31365 1627 31399
rect 30297 30821 30331 30855
rect 30113 30685 30147 30719
rect 30757 30685 30791 30719
rect 19533 30209 19567 30243
rect 38025 30209 38059 30243
rect 1593 30141 1627 30175
rect 1869 30141 1903 30175
rect 19441 30005 19475 30039
rect 38209 30005 38243 30039
rect 1593 29801 1627 29835
rect 20545 29257 20579 29291
rect 30849 29257 30883 29291
rect 20361 29121 20395 29155
rect 21005 29121 21039 29155
rect 30941 29121 30975 29155
rect 31401 29121 31435 29155
rect 38025 29121 38059 29155
rect 38209 28985 38243 29019
rect 30665 28169 30699 28203
rect 1869 28033 1903 28067
rect 30573 28033 30607 28067
rect 1685 27897 1719 27931
rect 31217 27829 31251 27863
rect 23029 27557 23063 27591
rect 22569 27421 22603 27455
rect 22477 27285 22511 27319
rect 38301 27285 38335 27319
rect 18797 27081 18831 27115
rect 1869 26945 1903 26979
rect 15393 26945 15427 26979
rect 16037 26945 16071 26979
rect 18245 26945 18279 26979
rect 38025 26877 38059 26911
rect 38301 26877 38335 26911
rect 1685 26741 1719 26775
rect 15945 26741 15979 26775
rect 18153 26741 18187 26775
rect 14381 26537 14415 26571
rect 20453 26537 20487 26571
rect 37841 26537 37875 26571
rect 14473 26333 14507 26367
rect 19901 26333 19935 26367
rect 38025 26333 38059 26367
rect 15025 26265 15059 26299
rect 19809 26265 19843 26299
rect 33609 25993 33643 26027
rect 33793 25857 33827 25891
rect 34253 25653 34287 25687
rect 38117 25653 38151 25687
rect 38025 25449 38059 25483
rect 37841 25245 37875 25279
rect 1869 24769 1903 24803
rect 20821 24769 20855 24803
rect 21373 24769 21407 24803
rect 38025 24769 38059 24803
rect 2421 24633 2455 24667
rect 20637 24633 20671 24667
rect 1685 24565 1719 24599
rect 38209 24565 38243 24599
rect 25237 24361 25271 24395
rect 34161 24361 34195 24395
rect 25053 24157 25087 24191
rect 25697 24157 25731 24191
rect 33977 24157 34011 24191
rect 33425 24021 33459 24055
rect 38025 23681 38059 23715
rect 38209 23477 38243 23511
rect 1777 23273 1811 23307
rect 1961 23069 1995 23103
rect 2421 22933 2455 22967
rect 37933 22729 37967 22763
rect 1869 22593 1903 22627
rect 37841 22593 37875 22627
rect 1685 22457 1719 22491
rect 7849 21981 7883 22015
rect 7665 21845 7699 21879
rect 8401 21845 8435 21879
rect 37657 21845 37691 21879
rect 1685 21505 1719 21539
rect 38025 21505 38059 21539
rect 1869 21369 1903 21403
rect 38209 21301 38243 21335
rect 1593 21097 1627 21131
rect 38025 21097 38059 21131
rect 37841 20893 37875 20927
rect 20361 20417 20395 20451
rect 20821 20417 20855 20451
rect 20269 20213 20303 20247
rect 27905 20009 27939 20043
rect 37657 19805 37691 19839
rect 38301 19805 38335 19839
rect 27261 19737 27295 19771
rect 27813 19737 27847 19771
rect 38117 19669 38151 19703
rect 1869 19329 1903 19363
rect 1593 19261 1627 19295
rect 1593 18921 1627 18955
rect 26157 18921 26191 18955
rect 25697 18717 25731 18751
rect 33149 18717 33183 18751
rect 25605 18581 25639 18615
rect 33057 18581 33091 18615
rect 18521 18309 18555 18343
rect 1869 18241 1903 18275
rect 19625 18241 19659 18275
rect 20085 18241 20119 18275
rect 19441 18173 19475 18207
rect 24869 18173 24903 18207
rect 25053 18173 25087 18207
rect 20821 18105 20855 18139
rect 1685 18037 1719 18071
rect 19257 18037 19291 18071
rect 20177 18037 20211 18071
rect 24685 18037 24719 18071
rect 19809 17833 19843 17867
rect 21649 17833 21683 17867
rect 25697 17833 25731 17867
rect 23029 17765 23063 17799
rect 19441 17697 19475 17731
rect 22385 17697 22419 17731
rect 19625 17629 19659 17663
rect 22569 17629 22603 17663
rect 23949 17629 23983 17663
rect 24593 17629 24627 17663
rect 24777 17629 24811 17663
rect 23857 17493 23891 17527
rect 25237 17493 25271 17527
rect 25145 17289 25179 17323
rect 18613 17221 18647 17255
rect 18705 17221 18739 17255
rect 22201 17221 22235 17255
rect 23857 17221 23891 17255
rect 23949 17221 23983 17255
rect 16221 17153 16255 17187
rect 17049 17153 17083 17187
rect 21465 17153 21499 17187
rect 24685 17153 24719 17187
rect 14841 17085 14875 17119
rect 19257 17085 19291 17119
rect 19441 17085 19475 17119
rect 22109 17085 22143 17119
rect 22385 17085 22419 17119
rect 23673 17085 23707 17119
rect 18153 17017 18187 17051
rect 15485 16949 15519 16983
rect 16129 16949 16163 16983
rect 16957 16949 16991 16983
rect 19625 16949 19659 16983
rect 21373 16949 21407 16983
rect 24593 16949 24627 16983
rect 19533 16745 19567 16779
rect 24685 16677 24719 16711
rect 14841 16609 14875 16643
rect 15485 16609 15519 16643
rect 22385 16609 22419 16643
rect 23121 16609 23155 16643
rect 17417 16541 17451 16575
rect 18705 16541 18739 16575
rect 19441 16541 19475 16575
rect 23305 16541 23339 16575
rect 23765 16541 23799 16575
rect 14933 16473 14967 16507
rect 16129 16473 16163 16507
rect 16221 16473 16255 16507
rect 16773 16473 16807 16507
rect 18153 16473 18187 16507
rect 21741 16473 21775 16507
rect 22293 16473 22327 16507
rect 25136 16473 25170 16507
rect 25237 16473 25271 16507
rect 17325 16405 17359 16439
rect 18797 16405 18831 16439
rect 13829 16201 13863 16235
rect 22569 16201 22603 16235
rect 24593 16201 24627 16235
rect 25237 16201 25271 16235
rect 32965 16201 32999 16235
rect 14473 16133 14507 16167
rect 14565 16133 14599 16167
rect 15761 16133 15795 16167
rect 23857 16133 23891 16167
rect 25789 16133 25823 16167
rect 1869 16065 1903 16099
rect 17049 16065 17083 16099
rect 17785 16065 17819 16099
rect 18429 16065 18463 16099
rect 18521 16065 18555 16099
rect 20545 16065 20579 16099
rect 22477 16065 22511 16099
rect 23121 16065 23155 16099
rect 24501 16065 24535 16099
rect 25145 16065 25179 16099
rect 33057 16065 33091 16099
rect 38025 16065 38059 16099
rect 13369 15997 13403 16031
rect 15669 15997 15703 16031
rect 16313 15997 16347 16031
rect 19441 15997 19475 16031
rect 19625 15997 19659 16031
rect 20729 15997 20763 16031
rect 23213 15997 23247 16031
rect 38301 15997 38335 16031
rect 15025 15929 15059 15963
rect 17141 15929 17175 15963
rect 1685 15861 1719 15895
rect 17877 15861 17911 15895
rect 20085 15861 20119 15895
rect 20913 15861 20947 15895
rect 23949 15861 23983 15895
rect 10701 15657 10735 15691
rect 13645 15657 13679 15691
rect 14657 15657 14691 15691
rect 17601 15657 17635 15691
rect 20729 15657 20763 15691
rect 21465 15657 21499 15691
rect 22017 15657 22051 15691
rect 23397 15657 23431 15691
rect 24593 15657 24627 15691
rect 31217 15657 31251 15691
rect 38301 15657 38335 15691
rect 15945 15521 15979 15555
rect 16221 15521 16255 15555
rect 18245 15521 18279 15555
rect 18521 15521 18555 15555
rect 19533 15521 19567 15555
rect 22661 15521 22695 15555
rect 23765 15521 23799 15555
rect 10609 15453 10643 15487
rect 11253 15453 11287 15487
rect 13553 15453 13587 15487
rect 14749 15453 14783 15487
rect 15209 15453 15243 15487
rect 17509 15453 17543 15487
rect 20821 15453 20855 15487
rect 21373 15453 21407 15487
rect 22477 15453 22511 15487
rect 23581 15453 23615 15487
rect 25053 15453 25087 15487
rect 25237 15453 25271 15487
rect 31125 15453 31159 15487
rect 16037 15385 16071 15419
rect 18337 15385 18371 15419
rect 19625 15385 19659 15419
rect 20177 15385 20211 15419
rect 12173 15317 12207 15351
rect 13093 15317 13127 15351
rect 15301 15317 15335 15351
rect 1777 15113 1811 15147
rect 4077 15113 4111 15147
rect 10793 15113 10827 15147
rect 15577 15113 15611 15147
rect 19349 15113 19383 15147
rect 19993 15113 20027 15147
rect 24869 15113 24903 15147
rect 17049 15045 17083 15079
rect 18245 15045 18279 15079
rect 20821 15045 20855 15079
rect 22109 15045 22143 15079
rect 22201 15045 22235 15079
rect 24133 15045 24167 15079
rect 1961 14977 1995 15011
rect 2421 14977 2455 15011
rect 4261 14977 4295 15011
rect 4813 14977 4847 15011
rect 10149 14977 10183 15011
rect 10701 14977 10735 15011
rect 12265 14977 12299 15011
rect 13093 14977 13127 15011
rect 13553 14977 13587 15011
rect 14197 14977 14231 15011
rect 15025 14977 15059 15011
rect 15485 14977 15519 15011
rect 19257 14977 19291 15011
rect 19901 14977 19935 15011
rect 21281 14977 21315 15011
rect 24777 14977 24811 15011
rect 16313 14909 16347 14943
rect 16957 14909 16991 14943
rect 18153 14909 18187 14943
rect 21373 14909 21407 14943
rect 23121 14909 23155 14943
rect 23581 14909 23615 14943
rect 24225 14909 24259 14943
rect 14841 14841 14875 14875
rect 17509 14841 17543 14875
rect 18705 14841 18739 14875
rect 12173 14773 12207 14807
rect 13001 14773 13035 14807
rect 13645 14773 13679 14807
rect 14289 14773 14323 14807
rect 18429 14569 18463 14603
rect 15025 14433 15059 14467
rect 15945 14433 15979 14467
rect 16221 14433 16255 14467
rect 17233 14433 17267 14467
rect 17693 14433 17727 14467
rect 20085 14433 20119 14467
rect 21373 14433 21407 14467
rect 22937 14433 22971 14467
rect 23213 14433 23247 14467
rect 24685 14433 24719 14467
rect 25237 14433 25271 14467
rect 12265 14365 12299 14399
rect 13553 14365 13587 14399
rect 18521 14365 18555 14399
rect 20821 14365 20855 14399
rect 24593 14365 24627 14399
rect 26065 14365 26099 14399
rect 26709 14365 26743 14399
rect 38025 14365 38059 14399
rect 38301 14365 38335 14399
rect 10609 14297 10643 14331
rect 11161 14297 11195 14331
rect 11253 14297 11287 14331
rect 11805 14297 11839 14331
rect 13093 14297 13127 14331
rect 14381 14297 14415 14331
rect 14473 14297 14507 14331
rect 16037 14297 16071 14331
rect 17325 14297 17359 14331
rect 19441 14297 19475 14331
rect 19993 14297 20027 14331
rect 21465 14297 21499 14331
rect 22385 14297 22419 14331
rect 23029 14297 23063 14331
rect 1685 14229 1719 14263
rect 12357 14229 12391 14263
rect 13645 14229 13679 14263
rect 20729 14229 20763 14263
rect 25973 14229 26007 14263
rect 26617 14229 26651 14263
rect 27261 14229 27295 14263
rect 10609 14025 10643 14059
rect 12173 14025 12207 14059
rect 18153 14025 18187 14059
rect 38301 14025 38335 14059
rect 13277 13957 13311 13991
rect 14565 13957 14599 13991
rect 15117 13957 15151 13991
rect 15761 13957 15795 13991
rect 16957 13957 16991 13991
rect 17049 13957 17083 13991
rect 19533 13957 19567 13991
rect 19625 13957 19659 13991
rect 22201 13957 22235 13991
rect 23121 13957 23155 13991
rect 24593 13957 24627 13991
rect 26065 13957 26099 13991
rect 1685 13889 1719 13923
rect 1869 13889 1903 13923
rect 12265 13889 12299 13923
rect 18061 13889 18095 13923
rect 20453 13889 20487 13923
rect 27169 13889 27203 13923
rect 12725 13821 12759 13855
rect 13369 13821 13403 13855
rect 14473 13821 14507 13855
rect 15669 13821 15703 13855
rect 15945 13821 15979 13855
rect 19349 13821 19383 13855
rect 20637 13821 20671 13855
rect 22109 13821 22143 13855
rect 24409 13821 24443 13855
rect 24685 13821 24719 13855
rect 26157 13821 26191 13855
rect 17509 13753 17543 13787
rect 25605 13753 25639 13787
rect 11161 13685 11195 13719
rect 21097 13685 21131 13719
rect 27813 13685 27847 13719
rect 11069 13481 11103 13515
rect 13001 13481 13035 13515
rect 19901 13481 19935 13515
rect 21833 13481 21867 13515
rect 27997 13481 28031 13515
rect 9965 13413 9999 13447
rect 13645 13413 13679 13447
rect 18245 13413 18279 13447
rect 22477 13413 22511 13447
rect 12357 13345 12391 13379
rect 15025 13345 15059 13379
rect 17049 13345 17083 13379
rect 17325 13345 17359 13379
rect 20637 13345 20671 13379
rect 21281 13345 21315 13379
rect 23029 13345 23063 13379
rect 24041 13345 24075 13379
rect 25237 13345 25271 13379
rect 27353 13345 27387 13379
rect 1961 13277 1995 13311
rect 10977 13277 11011 13311
rect 11621 13277 11655 13311
rect 12265 13277 12299 13311
rect 12909 13277 12943 13311
rect 13737 13277 13771 13311
rect 14289 13277 14323 13311
rect 19809 13277 19843 13311
rect 21741 13277 21775 13311
rect 28089 13277 28123 13311
rect 28549 13277 28583 13311
rect 9413 13209 9447 13243
rect 10517 13209 10551 13243
rect 15117 13209 15151 13243
rect 15669 13209 15703 13243
rect 17233 13209 17267 13243
rect 18705 13209 18739 13243
rect 18797 13209 18831 13243
rect 20729 13209 20763 13243
rect 23121 13209 23155 13243
rect 24593 13209 24627 13243
rect 25145 13209 25179 13243
rect 26433 13209 26467 13243
rect 26525 13209 26559 13243
rect 1777 13141 1811 13175
rect 2513 13141 2547 13175
rect 11805 13141 11839 13175
rect 14381 13141 14415 13175
rect 16221 13141 16255 13175
rect 25881 13141 25915 13175
rect 9229 12937 9263 12971
rect 9873 12937 9907 12971
rect 23029 12937 23063 12971
rect 23489 12937 23523 12971
rect 24593 12937 24627 12971
rect 27261 12937 27295 12971
rect 27905 12937 27939 12971
rect 28825 12937 28859 12971
rect 7757 12869 7791 12903
rect 12081 12869 12115 12903
rect 14013 12869 14047 12903
rect 15669 12869 15703 12903
rect 17417 12869 17451 12903
rect 17509 12869 17543 12903
rect 18245 12869 18279 12903
rect 18797 12869 18831 12903
rect 20085 12869 20119 12903
rect 20177 12869 20211 12903
rect 1869 12801 1903 12835
rect 7665 12801 7699 12835
rect 8309 12801 8343 12835
rect 10333 12801 10367 12835
rect 13185 12801 13219 12835
rect 20821 12801 20855 12835
rect 22385 12801 22419 12835
rect 24133 12801 24167 12835
rect 25053 12801 25087 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 27997 12801 28031 12835
rect 28917 12801 28951 12835
rect 11161 12733 11195 12767
rect 11989 12733 12023 12767
rect 13921 12733 13955 12767
rect 14197 12733 14231 12767
rect 15301 12733 15335 12767
rect 15761 12733 15795 12767
rect 16865 12733 16899 12767
rect 18889 12733 18923 12767
rect 21005 12733 21039 12767
rect 22569 12733 22603 12767
rect 23949 12733 23983 12767
rect 25237 12733 25271 12767
rect 26249 12733 26283 12767
rect 29377 12733 29411 12767
rect 38025 12733 38059 12767
rect 38301 12733 38335 12767
rect 12541 12665 12575 12699
rect 19625 12665 19659 12699
rect 21189 12665 21223 12699
rect 26065 12665 26099 12699
rect 1685 12597 1719 12631
rect 10425 12597 10459 12631
rect 13277 12597 13311 12631
rect 30113 12597 30147 12631
rect 7481 12393 7515 12427
rect 14841 12393 14875 12427
rect 17049 12393 17083 12427
rect 18797 12393 18831 12427
rect 20453 12393 20487 12427
rect 23765 12393 23799 12427
rect 26065 12393 26099 12427
rect 27629 12393 27663 12427
rect 9229 12325 9263 12359
rect 19809 12325 19843 12359
rect 29837 12325 29871 12359
rect 38301 12325 38335 12359
rect 12725 12257 12759 12291
rect 15485 12257 15519 12291
rect 17601 12257 17635 12291
rect 22661 12257 22695 12291
rect 23121 12257 23155 12291
rect 25237 12257 25271 12291
rect 26249 12257 26283 12291
rect 7573 12189 7607 12223
rect 10241 12189 10275 12223
rect 10885 12189 10919 12223
rect 11713 12189 11747 12223
rect 13553 12189 13587 12223
rect 14749 12189 14783 12223
rect 18705 12189 18739 12223
rect 19717 12189 19751 12223
rect 20545 12189 20579 12223
rect 23857 12189 23891 12223
rect 26433 12189 26467 12223
rect 27077 12189 27111 12223
rect 27537 12189 27571 12223
rect 28181 12189 28215 12223
rect 29009 12189 29043 12223
rect 29929 12189 29963 12223
rect 9781 12121 9815 12155
rect 10333 12121 10367 12155
rect 12265 12121 12299 12155
rect 12357 12121 12391 12155
rect 13645 12121 13679 12155
rect 15577 12121 15611 12155
rect 16497 12121 16531 12155
rect 17693 12121 17727 12155
rect 18245 12121 18279 12155
rect 21005 12121 21039 12155
rect 21557 12121 21591 12155
rect 21649 12121 21683 12155
rect 23052 12121 23086 12155
rect 24593 12121 24627 12155
rect 25145 12121 25179 12155
rect 26985 12121 27019 12155
rect 8585 12053 8619 12087
rect 10977 12053 11011 12087
rect 11621 12053 11655 12087
rect 28273 12053 28307 12087
rect 28917 12053 28951 12087
rect 30389 12053 30423 12087
rect 10425 11849 10459 11883
rect 15577 11849 15611 11883
rect 16221 11849 16255 11883
rect 19625 11849 19659 11883
rect 23949 11849 23983 11883
rect 25973 11849 26007 11883
rect 27261 11849 27295 11883
rect 28549 11849 28583 11883
rect 8309 11781 8343 11815
rect 13369 11781 13403 11815
rect 14105 11781 14139 11815
rect 14197 11781 14231 11815
rect 14749 11781 14783 11815
rect 17049 11781 17083 11815
rect 18521 11781 18555 11815
rect 18613 11781 18647 11815
rect 21281 11781 21315 11815
rect 21373 11781 21407 11815
rect 22385 11781 22419 11815
rect 22477 11781 22511 11815
rect 24777 11781 24811 11815
rect 9321 11713 9355 11747
rect 10333 11713 10367 11747
rect 10977 11713 11011 11747
rect 12173 11713 12207 11747
rect 12817 11713 12851 11747
rect 15485 11713 15519 11747
rect 16129 11713 16163 11747
rect 19165 11713 19199 11747
rect 20729 11713 20763 11747
rect 23857 11713 23891 11747
rect 24593 11713 24627 11747
rect 25513 11713 25547 11747
rect 26433 11713 26467 11747
rect 27169 11713 27203 11747
rect 27997 11713 28031 11747
rect 28641 11713 28675 11747
rect 29285 11713 29319 11747
rect 8861 11645 8895 11679
rect 13461 11645 13495 11679
rect 16957 11645 16991 11679
rect 17877 11645 17911 11679
rect 20085 11645 20119 11679
rect 20269 11645 20303 11679
rect 22661 11645 22695 11679
rect 25329 11645 25363 11679
rect 26525 11645 26559 11679
rect 27905 11645 27939 11679
rect 11069 11577 11103 11611
rect 30389 11577 30423 11611
rect 9413 11509 9447 11543
rect 12265 11509 12299 11543
rect 29193 11509 29227 11543
rect 29745 11509 29779 11543
rect 30941 11509 30975 11543
rect 38301 11509 38335 11543
rect 9965 11305 9999 11339
rect 10609 11305 10643 11339
rect 21005 11305 21039 11339
rect 23949 11305 23983 11339
rect 25789 11305 25823 11339
rect 9413 11237 9447 11271
rect 11253 11237 11287 11271
rect 27077 11237 27111 11271
rect 11897 11169 11931 11203
rect 13369 11169 13403 11203
rect 17049 11169 17083 11203
rect 17877 11169 17911 11203
rect 18889 11169 18923 11203
rect 19625 11169 19659 11203
rect 20085 11169 20119 11203
rect 21649 11169 21683 11203
rect 22753 11169 22787 11203
rect 24593 11169 24627 11203
rect 27721 11169 27755 11203
rect 8493 11101 8527 11135
rect 10057 11101 10091 11135
rect 10701 11101 10735 11135
rect 11345 11101 11379 11135
rect 12541 11101 12575 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 15209 11101 15243 11135
rect 20913 11101 20947 11135
rect 22937 11101 22971 11135
rect 23397 11101 23431 11135
rect 23849 11101 23883 11135
rect 24777 11101 24811 11135
rect 25881 11101 25915 11135
rect 26525 11101 26559 11135
rect 27169 11101 27203 11135
rect 28917 11101 28951 11135
rect 29929 11101 29963 11135
rect 30389 11101 30423 11135
rect 38025 11101 38059 11135
rect 38301 11101 38335 11135
rect 11989 11033 12023 11067
rect 13553 11033 13587 11067
rect 13645 11033 13679 11067
rect 15761 11033 15795 11067
rect 15853 11033 15887 11067
rect 16405 11033 16439 11067
rect 16957 11033 16991 11067
rect 17969 11033 18003 11067
rect 19717 11033 19751 11067
rect 21741 11033 21775 11067
rect 22293 11033 22327 11067
rect 26433 11033 26467 11067
rect 28273 11033 28307 11067
rect 28365 11033 28399 11067
rect 30481 11033 30515 11067
rect 31125 11033 31159 11067
rect 25237 10965 25271 10999
rect 29837 10965 29871 10999
rect 9873 10761 9907 10795
rect 11069 10761 11103 10795
rect 21097 10761 21131 10795
rect 23581 10761 23615 10795
rect 24777 10761 24811 10795
rect 25973 10761 26007 10795
rect 27629 10761 27663 10795
rect 8677 10693 8711 10727
rect 10425 10693 10459 10727
rect 12173 10693 12207 10727
rect 12725 10693 12759 10727
rect 13369 10693 13403 10727
rect 14565 10693 14599 10727
rect 15761 10693 15795 10727
rect 17233 10693 17267 10727
rect 18429 10693 18463 10727
rect 18981 10693 19015 10727
rect 19625 10693 19659 10727
rect 22937 10693 22971 10727
rect 1869 10625 1903 10659
rect 10333 10625 10367 10659
rect 10977 10625 11011 10659
rect 13921 10625 13955 10659
rect 16313 10625 16347 10659
rect 21005 10625 21039 10659
rect 24225 10625 24259 10659
rect 28089 10625 28123 10659
rect 28273 10625 28307 10659
rect 28733 10625 28767 10659
rect 29561 10625 29595 10659
rect 30021 10625 30055 10659
rect 30849 10625 30883 10659
rect 37841 10625 37875 10659
rect 12081 10557 12115 10591
rect 13277 10557 13311 10591
rect 14473 10557 14507 10591
rect 15669 10557 15703 10591
rect 17141 10557 17175 10591
rect 17417 10557 17451 10591
rect 18337 10557 18371 10591
rect 19533 10557 19567 10591
rect 20545 10557 20579 10591
rect 22017 10557 22051 10591
rect 23029 10557 23063 10591
rect 24041 10557 24075 10591
rect 25237 10557 25271 10591
rect 25421 10557 25455 10591
rect 26433 10557 26467 10591
rect 26617 10557 26651 10591
rect 29469 10557 29503 10591
rect 15025 10489 15059 10523
rect 30757 10489 30791 10523
rect 1685 10421 1719 10455
rect 9137 10421 9171 10455
rect 28825 10421 28859 10455
rect 30113 10421 30147 10455
rect 31401 10421 31435 10455
rect 38025 10421 38059 10455
rect 9413 10217 9447 10251
rect 13001 10217 13035 10251
rect 13645 10217 13679 10251
rect 29837 10217 29871 10251
rect 16589 10149 16623 10183
rect 18889 10149 18923 10183
rect 22569 10149 22603 10183
rect 10425 10081 10459 10115
rect 11069 10081 11103 10115
rect 14289 10081 14323 10115
rect 17141 10081 17175 10115
rect 17417 10081 17451 10115
rect 21373 10081 21407 10115
rect 23305 10081 23339 10115
rect 23949 10081 23983 10115
rect 24685 10081 24719 10115
rect 26985 10081 27019 10115
rect 27261 10081 27295 10115
rect 28549 10081 28583 10115
rect 28733 10081 28767 10115
rect 30389 10081 30423 10115
rect 9505 10013 9539 10047
rect 13093 10013 13127 10047
rect 13553 10013 13587 10047
rect 16037 10013 16071 10047
rect 16497 10013 16531 10047
rect 19441 10013 19475 10047
rect 26341 10013 26375 10047
rect 29929 10013 29963 10047
rect 10977 9945 11011 9979
rect 11621 9945 11655 9979
rect 12173 9945 12207 9979
rect 12265 9945 12299 9979
rect 15761 9945 15795 9979
rect 19533 9945 19567 9979
rect 20361 9945 20395 9979
rect 21281 9945 21315 9979
rect 22006 9945 22040 9979
rect 22109 9945 22143 9979
rect 23857 9945 23891 9979
rect 24777 9945 24811 9979
rect 25697 9945 25731 9979
rect 27077 9945 27111 9979
rect 31033 9945 31067 9979
rect 26249 9877 26283 9911
rect 28089 9877 28123 9911
rect 9873 9605 9907 9639
rect 10425 9605 10459 9639
rect 12909 9605 12943 9639
rect 13461 9605 13495 9639
rect 17049 9605 17083 9639
rect 23581 9605 23615 9639
rect 24961 9605 24995 9639
rect 25053 9605 25087 9639
rect 27721 9605 27755 9639
rect 28733 9605 28767 9639
rect 29285 9605 29319 9639
rect 10333 9537 10367 9571
rect 11161 9537 11195 9571
rect 12081 9537 12115 9571
rect 21005 9537 21039 9571
rect 30389 9537 30423 9571
rect 11069 9469 11103 9503
rect 12817 9469 12851 9503
rect 15761 9469 15795 9503
rect 16313 9469 16347 9503
rect 16957 9469 16991 9503
rect 17877 9469 17911 9503
rect 20545 9469 20579 9503
rect 21097 9469 21131 9503
rect 22109 9469 22143 9503
rect 23857 9469 23891 9503
rect 26433 9469 26467 9503
rect 26617 9469 26651 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 28641 9469 28675 9503
rect 29745 9469 29779 9503
rect 9321 9401 9355 9435
rect 24501 9401 24535 9435
rect 8677 9333 8711 9367
rect 12173 9333 12207 9367
rect 14013 9333 14047 9367
rect 15503 9333 15537 9367
rect 18797 9333 18831 9367
rect 20287 9333 20321 9367
rect 26249 9333 26283 9367
rect 30481 9333 30515 9367
rect 11069 9129 11103 9163
rect 11713 9129 11747 9163
rect 13001 9129 13035 9163
rect 23397 9129 23431 9163
rect 23949 9129 23983 9163
rect 1869 9061 1903 9095
rect 12357 9061 12391 9095
rect 13645 9061 13679 9095
rect 20177 9061 20211 9095
rect 22753 9061 22787 9095
rect 31493 9061 31527 9095
rect 9413 8993 9447 9027
rect 14289 8993 14323 9027
rect 18613 8993 18647 9027
rect 25789 8993 25823 9027
rect 27353 8993 27387 9027
rect 27538 8993 27572 9027
rect 27997 8993 28031 9027
rect 29837 8993 29871 9027
rect 30481 8993 30515 9027
rect 11161 8925 11195 8959
rect 11621 8925 11655 8959
rect 12449 8925 12483 8959
rect 13093 8925 13127 8959
rect 13553 8925 13587 8959
rect 16865 8925 16899 8959
rect 21005 8925 21039 8959
rect 23489 8925 23523 8959
rect 25605 8925 25639 8959
rect 26709 8925 26743 8959
rect 26893 8925 26927 8959
rect 28917 8925 28951 8959
rect 29101 8925 29135 8959
rect 38025 8925 38059 8959
rect 1685 8857 1719 8891
rect 8585 8857 8619 8891
rect 14565 8857 14599 8891
rect 17141 8857 17175 8891
rect 19625 8857 19659 8891
rect 19717 8857 19751 8891
rect 21281 8857 21315 8891
rect 24593 8857 24627 8891
rect 29929 8857 29963 8891
rect 9873 8789 9907 8823
rect 10425 8789 10459 8823
rect 16037 8789 16071 8823
rect 25145 8789 25179 8823
rect 26249 8789 26283 8823
rect 28457 8789 28491 8823
rect 30941 8789 30975 8823
rect 38209 8789 38243 8823
rect 1685 8585 1719 8619
rect 12265 8585 12299 8619
rect 19073 8585 19107 8619
rect 26249 8585 26283 8619
rect 27261 8585 27295 8619
rect 30389 8585 30423 8619
rect 16037 8517 16071 8551
rect 21189 8517 21223 8551
rect 23765 8517 23799 8551
rect 24777 8517 24811 8551
rect 28273 8517 28307 8551
rect 29193 8517 29227 8551
rect 14013 8449 14047 8483
rect 16306 8449 16340 8483
rect 17325 8449 17359 8483
rect 21465 8449 21499 8483
rect 24041 8449 24075 8483
rect 24501 8449 24535 8483
rect 27353 8449 27387 8483
rect 29653 8449 29687 8483
rect 30481 8449 30515 8483
rect 13737 8381 13771 8415
rect 14565 8381 14599 8415
rect 17601 8381 17635 8415
rect 22017 8381 22051 8415
rect 28181 8381 28215 8415
rect 32321 8381 32355 8415
rect 19717 8313 19751 8347
rect 9505 8245 9539 8279
rect 9965 8245 9999 8279
rect 10517 8245 10551 8279
rect 11069 8245 11103 8279
rect 29745 8245 29779 8279
rect 31033 8245 31067 8279
rect 31585 8245 31619 8279
rect 11345 8041 11379 8075
rect 13645 8041 13679 8075
rect 14473 8041 14507 8075
rect 15117 8041 15151 8075
rect 21207 8041 21241 8075
rect 24685 8041 24719 8075
rect 25329 8041 25363 8075
rect 28917 8041 28951 8075
rect 29837 8041 29871 8075
rect 30481 8041 30515 8075
rect 31769 8041 31803 8075
rect 31125 7973 31159 8007
rect 15669 7905 15703 7939
rect 17693 7905 17727 7939
rect 18245 7905 18279 7939
rect 24041 7905 24075 7939
rect 26801 7905 26835 7939
rect 27077 7905 27111 7939
rect 27629 7905 27663 7939
rect 28273 7905 28307 7939
rect 11437 7837 11471 7871
rect 11897 7837 11931 7871
rect 14565 7837 14599 7871
rect 15209 7837 15243 7871
rect 18889 7837 18923 7871
rect 21465 7837 21499 7871
rect 22017 7837 22051 7871
rect 24777 7837 24811 7871
rect 25421 7837 25455 7871
rect 28825 7837 28859 7871
rect 29929 7837 29963 7871
rect 30573 7837 30607 7871
rect 31217 7837 31251 7871
rect 12173 7769 12207 7803
rect 15945 7769 15979 7803
rect 19441 7769 19475 7803
rect 22293 7769 22327 7803
rect 26985 7769 27019 7803
rect 28181 7769 28215 7803
rect 32229 7769 32263 7803
rect 9689 7701 9723 7735
rect 10241 7701 10275 7735
rect 10793 7701 10827 7735
rect 11069 7497 11103 7531
rect 18153 7497 18187 7531
rect 21373 7497 21407 7531
rect 23765 7497 23799 7531
rect 24409 7497 24443 7531
rect 25053 7497 25087 7531
rect 28457 7497 28491 7531
rect 29101 7497 29135 7531
rect 30389 7497 30423 7531
rect 1869 7429 1903 7463
rect 9965 7429 9999 7463
rect 13369 7429 13403 7463
rect 14381 7429 14415 7463
rect 16957 7429 16991 7463
rect 18981 7429 19015 7463
rect 22293 7429 22327 7463
rect 26433 7429 26467 7463
rect 27169 7429 27203 7463
rect 27721 7429 27755 7463
rect 29745 7429 29779 7463
rect 1685 7361 1719 7395
rect 11161 7361 11195 7395
rect 17601 7361 17635 7395
rect 18245 7361 18279 7395
rect 18705 7361 18739 7395
rect 20729 7361 20763 7395
rect 21281 7361 21315 7395
rect 24501 7361 24535 7395
rect 24961 7361 24995 7395
rect 28365 7361 28399 7395
rect 29009 7361 29043 7395
rect 29653 7361 29687 7395
rect 30481 7361 30515 7395
rect 31125 7361 31159 7395
rect 38025 7361 38059 7395
rect 8861 7293 8895 7327
rect 13645 7293 13679 7327
rect 14105 7293 14139 7327
rect 22017 7293 22051 7327
rect 26157 7293 26191 7327
rect 26525 7293 26559 7327
rect 27813 7293 27847 7327
rect 38301 7293 38335 7327
rect 9413 7225 9447 7259
rect 11897 7225 11931 7259
rect 15853 7225 15887 7259
rect 17509 7225 17543 7259
rect 31033 7225 31067 7259
rect 31677 7225 31711 7259
rect 10425 7157 10459 7191
rect 32321 7157 32355 7191
rect 1593 6953 1627 6987
rect 17404 6953 17438 6987
rect 19704 6953 19738 6987
rect 21833 6953 21867 6987
rect 29837 6953 29871 6987
rect 12541 6885 12575 6919
rect 28917 6885 28951 6919
rect 38301 6885 38335 6919
rect 10885 6817 10919 6851
rect 11437 6817 11471 6851
rect 13645 6817 13679 6851
rect 14289 6817 14323 6851
rect 16037 6817 16071 6851
rect 16589 6817 16623 6851
rect 17141 6817 17175 6851
rect 19441 6817 19475 6851
rect 23581 6817 23615 6851
rect 27813 6817 27847 6851
rect 9781 6749 9815 6783
rect 13553 6749 13587 6783
rect 16497 6749 16531 6783
rect 24593 6749 24627 6783
rect 25329 6749 25363 6783
rect 25421 6749 25455 6783
rect 27169 6749 27203 6783
rect 27261 6749 27295 6783
rect 29929 6749 29963 6783
rect 30573 6749 30607 6783
rect 31217 6749 31251 6783
rect 31861 6749 31895 6783
rect 9137 6681 9171 6715
rect 14565 6681 14599 6715
rect 23305 6681 23339 6715
rect 24685 6681 24719 6715
rect 25881 6681 25915 6715
rect 26433 6681 26467 6715
rect 26525 6681 26559 6715
rect 28365 6681 28399 6715
rect 28457 6681 28491 6715
rect 10241 6613 10275 6647
rect 11897 6613 11931 6647
rect 13093 6613 13127 6647
rect 18889 6613 18923 6647
rect 21189 6613 21223 6647
rect 30481 6613 30515 6647
rect 31125 6613 31159 6647
rect 31769 6613 31803 6647
rect 32413 6613 32447 6647
rect 32873 6613 32907 6647
rect 33425 6613 33459 6647
rect 33977 6613 34011 6647
rect 37657 6613 37691 6647
rect 4537 6409 4571 6443
rect 10609 6409 10643 6443
rect 16221 6409 16255 6443
rect 27905 6409 27939 6443
rect 28641 6409 28675 6443
rect 32413 6409 32447 6443
rect 19533 6341 19567 6375
rect 26525 6341 26559 6375
rect 27261 6341 27295 6375
rect 30573 6341 30607 6375
rect 4445 6273 4479 6307
rect 5181 6273 5215 6307
rect 8125 6273 8159 6307
rect 9137 6273 9171 6307
rect 16129 6273 16163 6307
rect 18797 6273 18831 6307
rect 19257 6273 19291 6307
rect 24225 6273 24259 6307
rect 26433 6273 26467 6307
rect 27353 6273 27387 6307
rect 27997 6273 28031 6307
rect 28733 6273 28767 6307
rect 29377 6273 29411 6307
rect 30021 6273 30055 6307
rect 30665 6273 30699 6307
rect 31309 6273 31343 6307
rect 32505 6273 32539 6307
rect 15301 6205 15335 6239
rect 15577 6205 15611 6239
rect 18521 6205 18555 6239
rect 22017 6205 22051 6239
rect 22293 6205 22327 6239
rect 24501 6205 24535 6239
rect 8585 6137 8619 6171
rect 11161 6137 11195 6171
rect 12173 6137 12207 6171
rect 12725 6137 12759 6171
rect 13277 6137 13311 6171
rect 17049 6137 17083 6171
rect 21005 6137 21039 6171
rect 23765 6137 23799 6171
rect 29929 6137 29963 6171
rect 33057 6137 33091 6171
rect 9229 6069 9263 6103
rect 10057 6069 10091 6103
rect 13829 6069 13863 6103
rect 25973 6069 26007 6103
rect 29285 6069 29319 6103
rect 31217 6069 31251 6103
rect 33517 6069 33551 6103
rect 34069 6069 34103 6103
rect 37473 6069 37507 6103
rect 38301 6069 38335 6103
rect 4169 5865 4203 5899
rect 8033 5865 8067 5899
rect 10057 5865 10091 5899
rect 16313 5865 16347 5899
rect 19533 5865 19567 5899
rect 23323 5865 23357 5899
rect 26341 5865 26375 5899
rect 27537 5865 27571 5899
rect 28181 5865 28215 5899
rect 29837 5865 29871 5899
rect 30481 5865 30515 5899
rect 31125 5865 31159 5899
rect 31769 5865 31803 5899
rect 35449 5865 35483 5899
rect 3341 5797 3375 5831
rect 13737 5797 13771 5831
rect 18889 5797 18923 5831
rect 20177 5797 20211 5831
rect 26893 5797 26927 5831
rect 28825 5797 28859 5831
rect 38025 5797 38059 5831
rect 10609 5729 10643 5763
rect 11989 5729 12023 5763
rect 12265 5729 12299 5763
rect 14841 5729 14875 5763
rect 17141 5729 17175 5763
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 4721 5661 4755 5695
rect 11069 5661 11103 5695
rect 14565 5661 14599 5695
rect 19441 5661 19475 5695
rect 20085 5661 20119 5695
rect 20913 5661 20947 5695
rect 23581 5661 23615 5695
rect 24593 5661 24627 5695
rect 26801 5661 26835 5695
rect 27629 5661 27663 5695
rect 28089 5661 28123 5695
rect 28917 5661 28951 5695
rect 29929 5661 29963 5695
rect 30573 5661 30607 5695
rect 31217 5661 31251 5695
rect 31861 5661 31895 5695
rect 32505 5661 32539 5695
rect 33149 5661 33183 5695
rect 34897 5661 34931 5695
rect 9505 5593 9539 5627
rect 17417 5593 17451 5627
rect 21557 5593 21591 5627
rect 24869 5593 24903 5627
rect 32413 5593 32447 5627
rect 37565 5593 37599 5627
rect 38209 5593 38243 5627
rect 8493 5525 8527 5559
rect 11161 5525 11195 5559
rect 33057 5525 33091 5559
rect 33609 5525 33643 5559
rect 34161 5525 34195 5559
rect 36093 5525 36127 5559
rect 36645 5525 36679 5559
rect 3617 5321 3651 5355
rect 10517 5321 10551 5355
rect 13461 5321 13495 5355
rect 19717 5321 19751 5355
rect 23857 5321 23891 5355
rect 24593 5321 24627 5355
rect 25697 5321 25731 5355
rect 27261 5321 27295 5355
rect 27997 5321 28031 5355
rect 28641 5321 28675 5355
rect 29929 5321 29963 5355
rect 30573 5321 30607 5355
rect 34161 5321 34195 5355
rect 35265 5321 35299 5355
rect 7849 5253 7883 5287
rect 11989 5253 12023 5287
rect 15485 5253 15519 5287
rect 19257 5253 19291 5287
rect 33057 5253 33091 5287
rect 1869 5185 1903 5219
rect 7297 5185 7331 5219
rect 11161 5185 11195 5219
rect 11713 5185 11747 5219
rect 15761 5185 15795 5219
rect 16313 5185 16347 5219
rect 17233 5185 17267 5219
rect 24685 5185 24719 5219
rect 25881 5185 25915 5219
rect 26433 5185 26467 5219
rect 27353 5185 27387 5219
rect 28089 5185 28123 5219
rect 28733 5185 28767 5219
rect 29377 5185 29411 5219
rect 29837 5185 29871 5219
rect 30665 5185 30699 5219
rect 31309 5185 31343 5219
rect 32505 5185 32539 5219
rect 33149 5185 33183 5219
rect 1593 5117 1627 5151
rect 9505 5117 9539 5151
rect 14013 5117 14047 5151
rect 17509 5117 17543 5151
rect 21189 5117 21223 5151
rect 21465 5117 21499 5151
rect 22109 5117 22143 5151
rect 22385 5117 22419 5151
rect 34713 5117 34747 5151
rect 29285 5049 29319 5083
rect 31217 5049 31251 5083
rect 32413 5049 32447 5083
rect 8309 4981 8343 5015
rect 8953 4981 8987 5015
rect 10057 4981 10091 5015
rect 25145 4981 25179 5015
rect 26525 4981 26559 5015
rect 33609 4981 33643 5015
rect 35817 4981 35851 5015
rect 36369 4981 36403 5015
rect 38025 4981 38059 5015
rect 1593 4777 1627 4811
rect 9689 4777 9723 4811
rect 10149 4777 10183 4811
rect 10793 4777 10827 4811
rect 13553 4777 13587 4811
rect 14381 4777 14415 4811
rect 15871 4777 15905 4811
rect 28733 4777 28767 4811
rect 29837 4777 29871 4811
rect 31769 4777 31803 4811
rect 6929 4709 6963 4743
rect 11345 4709 11379 4743
rect 18797 4709 18831 4743
rect 21189 4709 21223 4743
rect 35449 4709 35483 4743
rect 16129 4641 16163 4675
rect 17049 4641 17083 4675
rect 17325 4641 17359 4675
rect 19441 4641 19475 4675
rect 28089 4641 28123 4675
rect 33701 4641 33735 4675
rect 6377 4573 6411 4607
rect 22017 4573 22051 4607
rect 24685 4573 24719 4607
rect 25789 4573 25823 4607
rect 25973 4573 26007 4607
rect 28181 4573 28215 4607
rect 28825 4573 28859 4607
rect 29929 4573 29963 4607
rect 30573 4573 30607 4607
rect 31217 4573 31251 4607
rect 31861 4573 31895 4607
rect 32505 4573 32539 4607
rect 32965 4573 32999 4607
rect 38301 4573 38335 4607
rect 7481 4505 7515 4539
rect 13645 4505 13679 4539
rect 19717 4505 19751 4539
rect 22293 4505 22327 4539
rect 26433 4505 26467 4539
rect 27353 4505 27387 4539
rect 27445 4505 27479 4539
rect 31125 4505 31159 4539
rect 32413 4505 32447 4539
rect 34989 4505 35023 4539
rect 36001 4505 36035 4539
rect 37105 4505 37139 4539
rect 8033 4437 8067 4471
rect 8493 4437 8527 4471
rect 11897 4437 11931 4471
rect 12449 4437 12483 4471
rect 13001 4437 13035 4471
rect 23765 4437 23799 4471
rect 24777 4437 24811 4471
rect 25329 4437 25363 4471
rect 30389 4437 30423 4471
rect 33149 4437 33183 4471
rect 34161 4437 34195 4471
rect 36553 4437 36587 4471
rect 38117 4437 38151 4471
rect 10057 4233 10091 4267
rect 10609 4233 10643 4267
rect 11897 4233 11931 4267
rect 12357 4233 12391 4267
rect 23765 4233 23799 4267
rect 25973 4233 26007 4267
rect 34805 4233 34839 4267
rect 36461 4233 36495 4267
rect 21465 4165 21499 4199
rect 27721 4165 27755 4199
rect 30113 4165 30147 4199
rect 38209 4165 38243 4199
rect 7297 4097 7331 4131
rect 14105 4097 14139 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 17601 4097 17635 4131
rect 19901 4097 19935 4131
rect 20729 4097 20763 4131
rect 22017 4097 22051 4131
rect 24225 4097 24259 4131
rect 26433 4097 26467 4131
rect 28917 4097 28951 4131
rect 29561 4097 29595 4131
rect 30205 4097 30239 4131
rect 30849 4097 30883 4131
rect 31493 4097 31527 4131
rect 32505 4097 32539 4131
rect 33149 4097 33183 4131
rect 33793 4097 33827 4131
rect 35357 4097 35391 4131
rect 35909 4097 35943 4131
rect 38025 4097 38059 4131
rect 6009 4029 6043 4063
rect 13829 4029 13863 4063
rect 14565 4029 14599 4063
rect 16037 4029 16071 4063
rect 17877 4029 17911 4063
rect 19349 4029 19383 4063
rect 22293 4029 22327 4063
rect 24501 4029 24535 4063
rect 27537 4029 27571 4063
rect 27813 4029 27847 4063
rect 29469 4029 29503 4063
rect 7757 3961 7791 3995
rect 8309 3961 8343 3995
rect 8861 3961 8895 3995
rect 9505 3961 9539 3995
rect 20637 3961 20671 3995
rect 28825 3961 28859 3995
rect 31401 3961 31435 3995
rect 34253 3961 34287 3995
rect 37473 3961 37507 3995
rect 1685 3893 1719 3927
rect 4445 3893 4479 3927
rect 6745 3893 6779 3927
rect 11161 3893 11195 3927
rect 17049 3893 17083 3927
rect 19993 3893 20027 3927
rect 26525 3893 26559 3927
rect 30757 3893 30791 3927
rect 32413 3893 32447 3927
rect 33057 3893 33091 3927
rect 33701 3893 33735 3927
rect 5549 3689 5583 3723
rect 9689 3689 9723 3723
rect 10333 3689 10367 3723
rect 29837 3689 29871 3723
rect 34345 3689 34379 3723
rect 34897 3689 34931 3723
rect 36001 3689 36035 3723
rect 7665 3621 7699 3655
rect 19625 3621 19659 3655
rect 1869 3553 1903 3587
rect 4261 3553 4295 3587
rect 11989 3553 12023 3587
rect 13737 3553 13771 3587
rect 16865 3553 16899 3587
rect 31769 3553 31803 3587
rect 35449 3553 35483 3587
rect 1685 3485 1719 3519
rect 4169 3485 4203 3519
rect 4905 3485 4939 3519
rect 7849 3485 7883 3519
rect 8309 3485 8343 3519
rect 10149 3485 10183 3519
rect 11253 3485 11287 3519
rect 14381 3485 14415 3519
rect 16405 3485 16439 3519
rect 19441 3485 19475 3519
rect 22569 3485 22603 3519
rect 23305 3485 23339 3519
rect 24041 3485 24075 3519
rect 24593 3485 24627 3519
rect 27537 3485 27571 3519
rect 28181 3485 28215 3519
rect 28733 3485 28767 3519
rect 28825 3485 28859 3519
rect 29745 3485 29779 3519
rect 30573 3485 30607 3519
rect 31217 3485 31251 3519
rect 31861 3485 31895 3519
rect 32505 3485 32539 3519
rect 33149 3485 33183 3519
rect 33793 3485 33827 3519
rect 37289 3485 37323 3519
rect 38025 3485 38059 3519
rect 7205 3417 7239 3451
rect 12265 3417 12299 3451
rect 14657 3417 14691 3451
rect 17141 3417 17175 3451
rect 20545 3417 20579 3451
rect 22293 3417 22327 3451
rect 24869 3417 24903 3451
rect 26893 3417 26927 3451
rect 26985 3417 27019 3451
rect 31125 3417 31159 3451
rect 33057 3417 33091 3451
rect 37013 3417 37047 3451
rect 3341 3349 3375 3383
rect 6009 3349 6043 3383
rect 6653 3349 6687 3383
rect 8493 3349 8527 3383
rect 11161 3349 11195 3383
rect 18613 3349 18647 3383
rect 23121 3349 23155 3383
rect 23857 3349 23891 3383
rect 26341 3349 26375 3383
rect 28089 3349 28123 3383
rect 30481 3349 30515 3383
rect 32413 3349 32447 3383
rect 33701 3349 33735 3383
rect 38209 3349 38243 3383
rect 2421 3145 2455 3179
rect 9781 3145 9815 3179
rect 11713 3145 11747 3179
rect 12357 3145 12391 3179
rect 23765 3145 23799 3179
rect 31585 3145 31619 3179
rect 4261 3077 4295 3111
rect 10333 3077 10367 3111
rect 10885 3077 10919 3111
rect 13829 3077 13863 3111
rect 19993 3077 20027 3111
rect 22293 3077 22327 3111
rect 33701 3077 33735 3111
rect 36277 3077 36311 3111
rect 1869 3009 1903 3043
rect 3709 3009 3743 3043
rect 4169 3009 4203 3043
rect 4813 3009 4847 3043
rect 7573 3009 7607 3043
rect 8033 3009 8067 3043
rect 8953 3009 8987 3043
rect 10241 3009 10275 3043
rect 11069 3009 11103 3043
rect 11897 3009 11931 3043
rect 14105 3009 14139 3043
rect 14565 3009 14599 3043
rect 16865 3009 16899 3043
rect 19257 3009 19291 3043
rect 19717 3009 19751 3043
rect 22017 3009 22051 3043
rect 25973 3009 26007 3043
rect 26617 3009 26651 3043
rect 28273 3009 28307 3043
rect 29101 3007 29135 3041
rect 29745 3009 29779 3043
rect 30389 3009 30423 3043
rect 30941 3009 30975 3043
rect 31033 3009 31067 3043
rect 31677 3009 31711 3043
rect 32505 3009 32539 3043
rect 33141 3009 33175 3043
rect 33793 3009 33827 3043
rect 34437 3009 34471 3043
rect 35081 3009 35115 3043
rect 36553 3009 36587 3043
rect 37473 3009 37507 3043
rect 7389 2941 7423 2975
rect 8309 2941 8343 2975
rect 14841 2941 14875 2975
rect 17141 2941 17175 2975
rect 21465 2941 21499 2975
rect 24225 2941 24259 2975
rect 25697 2941 25731 2975
rect 27629 2941 27663 2975
rect 27813 2941 27847 2975
rect 30297 2941 30331 2975
rect 35541 2941 35575 2975
rect 37657 2941 37691 2975
rect 3157 2873 3191 2907
rect 4905 2873 4939 2907
rect 27169 2873 27203 2907
rect 29653 2873 29687 2907
rect 32413 2873 32447 2907
rect 34345 2873 34379 2907
rect 1685 2805 1719 2839
rect 6009 2805 6043 2839
rect 6561 2805 6595 2839
rect 9137 2805 9171 2839
rect 16313 2805 16347 2839
rect 18613 2805 18647 2839
rect 26525 2805 26559 2839
rect 28457 2805 28491 2839
rect 29009 2805 29043 2839
rect 33057 2805 33091 2839
rect 34989 2805 35023 2839
rect 6009 2601 6043 2635
rect 7481 2601 7515 2635
rect 9229 2601 9263 2635
rect 33149 2601 33183 2635
rect 35817 2601 35851 2635
rect 2421 2533 2455 2567
rect 4169 2533 4203 2567
rect 11161 2533 11195 2567
rect 11989 2533 12023 2567
rect 17141 2533 17175 2567
rect 21281 2533 21315 2567
rect 32321 2533 32355 2567
rect 33609 2533 33643 2567
rect 10057 2465 10091 2499
rect 13737 2465 13771 2499
rect 14565 2465 14599 2499
rect 14841 2465 14875 2499
rect 16313 2465 16347 2499
rect 18889 2465 18923 2499
rect 19533 2465 19567 2499
rect 22109 2465 22143 2499
rect 22385 2465 22419 2499
rect 23857 2465 23891 2499
rect 25053 2465 25087 2499
rect 25513 2465 25547 2499
rect 36645 2465 36679 2499
rect 37473 2465 37507 2499
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 6837 2397 6871 2431
rect 8033 2397 8067 2431
rect 9781 2397 9815 2431
rect 25697 2397 25731 2431
rect 26433 2397 26467 2431
rect 27169 2397 27203 2431
rect 28733 2397 28767 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 31309 2397 31343 2431
rect 32505 2397 32539 2431
rect 33793 2397 33827 2431
rect 35173 2397 35207 2431
rect 35909 2397 35943 2431
rect 36921 2397 36955 2431
rect 37749 2397 37783 2431
rect 4905 2329 4939 2363
rect 8309 2329 8343 2363
rect 13461 2329 13495 2363
rect 18613 2329 18647 2363
rect 19809 2329 19843 2363
rect 27905 2329 27939 2363
rect 1685 2261 1719 2295
rect 3433 2261 3467 2295
rect 5457 2261 5491 2295
rect 6653 2261 6687 2295
rect 26249 2261 26283 2295
rect 27353 2261 27387 2295
rect 28549 2261 28583 2295
rect 29929 2261 29963 2295
rect 30573 2261 30607 2295
rect 31217 2261 31251 2295
rect 34989 2261 35023 2295
<< metal1 >>
rect 2958 37612 2964 37664
rect 3016 37652 3022 37664
rect 21818 37652 21824 37664
rect 3016 37624 21824 37652
rect 3016 37612 3022 37624
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 2958 37448 2964 37460
rect 2919 37420 2964 37448
rect 2958 37408 2964 37420
rect 3016 37408 3022 37460
rect 13538 37408 13544 37460
rect 13596 37448 13602 37460
rect 13633 37451 13691 37457
rect 13633 37448 13645 37451
rect 13596 37420 13645 37448
rect 13596 37408 13602 37420
rect 13633 37417 13645 37420
rect 13679 37417 13691 37451
rect 13633 37411 13691 37417
rect 14461 37451 14519 37457
rect 14461 37417 14473 37451
rect 14507 37448 14519 37451
rect 23014 37448 23020 37460
rect 14507 37420 23020 37448
rect 14507 37417 14519 37420
rect 14461 37411 14519 37417
rect 23014 37408 23020 37420
rect 23072 37408 23078 37460
rect 35069 37451 35127 37457
rect 35069 37417 35081 37451
rect 35115 37448 35127 37451
rect 35434 37448 35440 37460
rect 35115 37420 35440 37448
rect 35115 37417 35127 37420
rect 35069 37411 35127 37417
rect 35434 37408 35440 37420
rect 35492 37408 35498 37460
rect 36722 37448 36728 37460
rect 36683 37420 36728 37448
rect 36722 37408 36728 37420
rect 36780 37408 36786 37460
rect 2317 37383 2375 37389
rect 2317 37349 2329 37383
rect 2363 37380 2375 37383
rect 20530 37380 20536 37392
rect 2363 37352 20536 37380
rect 2363 37349 2375 37352
rect 2317 37343 2375 37349
rect 20530 37340 20536 37352
rect 20588 37340 20594 37392
rect 6733 37315 6791 37321
rect 6733 37281 6745 37315
rect 6779 37312 6791 37315
rect 7098 37312 7104 37324
rect 6779 37284 7104 37312
rect 6779 37281 6791 37284
rect 6733 37275 6791 37281
rect 7098 37272 7104 37284
rect 7156 37312 7162 37324
rect 7156 37284 7328 37312
rect 7156 37272 7162 37284
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2133 37247 2191 37253
rect 2133 37244 2145 37247
rect 2004 37216 2145 37244
rect 2004 37204 2010 37216
rect 2133 37213 2145 37216
rect 2179 37213 2191 37247
rect 2866 37244 2872 37256
rect 2827 37216 2872 37244
rect 2133 37207 2191 37213
rect 2866 37204 2872 37216
rect 2924 37204 2930 37256
rect 4249 37247 4307 37253
rect 4249 37213 4261 37247
rect 4295 37213 4307 37247
rect 5258 37244 5264 37256
rect 5219 37216 5264 37244
rect 4249 37207 4307 37213
rect 4264 37176 4292 37207
rect 5258 37204 5264 37216
rect 5316 37204 5322 37256
rect 7300 37253 7328 37284
rect 13538 37272 13544 37324
rect 13596 37312 13602 37324
rect 20622 37312 20628 37324
rect 13596 37284 14412 37312
rect 20583 37284 20628 37312
rect 13596 37272 13602 37284
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37213 7343 37247
rect 9398 37244 9404 37256
rect 9359 37216 9404 37244
rect 7285 37207 7343 37213
rect 9398 37204 9404 37216
rect 9456 37204 9462 37256
rect 10686 37244 10692 37256
rect 10647 37216 10692 37244
rect 10686 37204 10692 37216
rect 10744 37204 10750 37256
rect 12621 37247 12679 37253
rect 12621 37213 12633 37247
rect 12667 37244 12679 37247
rect 14274 37244 14280 37256
rect 12667 37216 14280 37244
rect 12667 37213 12679 37216
rect 12621 37207 12679 37213
rect 14274 37204 14280 37216
rect 14332 37204 14338 37256
rect 14384 37253 14412 37284
rect 20622 37272 20628 37284
rect 20680 37312 20686 37324
rect 22741 37315 22799 37321
rect 22741 37312 22753 37315
rect 20680 37284 22753 37312
rect 20680 37272 20686 37284
rect 22741 37281 22753 37284
rect 22787 37281 22799 37315
rect 22741 37275 22799 37281
rect 14369 37247 14427 37253
rect 14369 37213 14381 37247
rect 14415 37213 14427 37247
rect 15838 37244 15844 37256
rect 15799 37216 15844 37244
rect 14369 37207 14427 37213
rect 15838 37204 15844 37216
rect 15896 37204 15902 37256
rect 17126 37244 17132 37256
rect 17087 37216 17132 37244
rect 17126 37204 17132 37216
rect 17184 37244 17190 37256
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17184 37216 17601 37244
rect 17184 37204 17190 37216
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 17589 37207 17647 37213
rect 18414 37204 18420 37256
rect 18472 37244 18478 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 18472 37216 19441 37244
rect 18472 37204 18478 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 9490 37176 9496 37188
rect 4264 37148 9496 37176
rect 9490 37136 9496 37148
rect 9548 37136 9554 37188
rect 19334 37136 19340 37188
rect 19392 37176 19398 37188
rect 20916 37176 20944 37207
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21324 37216 22017 37244
rect 21324 37204 21330 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22005 37207 22063 37213
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25314 37244 25320 37256
rect 25275 37216 25320 37244
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26206 37216 27169 37244
rect 19392 37148 20944 37176
rect 19392 37136 19398 37148
rect 25222 37136 25228 37188
rect 25280 37176 25286 37188
rect 26206 37176 26234 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 27157 37207 27215 37213
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 30742 37244 30748 37256
rect 30703 37216 30748 37244
rect 30742 37204 30748 37216
rect 30800 37204 30806 37256
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37213 32367 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32309 37207 32367 37213
rect 25280 37148 26234 37176
rect 25280 37136 25286 37148
rect 30650 37136 30656 37188
rect 30708 37176 30714 37188
rect 32324 37176 32352 37207
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 35434 37204 35440 37256
rect 35492 37244 35498 37256
rect 35713 37247 35771 37253
rect 35713 37244 35725 37247
rect 35492 37216 35725 37244
rect 35492 37204 35498 37216
rect 35713 37213 35725 37216
rect 35759 37213 35771 37247
rect 36906 37244 36912 37256
rect 36867 37216 36912 37244
rect 35713 37207 35771 37213
rect 36906 37204 36912 37216
rect 36964 37204 36970 37256
rect 37458 37244 37464 37256
rect 37419 37216 37464 37244
rect 37458 37204 37464 37216
rect 37516 37204 37522 37256
rect 35526 37176 35532 37188
rect 30708 37148 32352 37176
rect 35487 37148 35532 37176
rect 30708 37136 30714 37148
rect 35526 37136 35532 37148
rect 35584 37136 35590 37188
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 4065 37111 4123 37117
rect 4065 37108 4077 37111
rect 3936 37080 4077 37108
rect 3936 37068 3942 37080
rect 4065 37077 4077 37080
rect 4111 37077 4123 37111
rect 4065 37071 4123 37077
rect 5166 37068 5172 37120
rect 5224 37108 5230 37120
rect 5445 37111 5503 37117
rect 5445 37108 5457 37111
rect 5224 37080 5457 37108
rect 5224 37068 5230 37080
rect 5445 37077 5457 37080
rect 5491 37077 5503 37111
rect 7374 37108 7380 37120
rect 7335 37080 7380 37108
rect 5445 37071 5503 37077
rect 7374 37068 7380 37080
rect 7432 37068 7438 37120
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 9217 37111 9275 37117
rect 9217 37108 9229 37111
rect 8444 37080 9229 37108
rect 8444 37068 8450 37080
rect 9217 37077 9229 37080
rect 9263 37077 9275 37111
rect 9217 37071 9275 37077
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10505 37111 10563 37117
rect 10505 37108 10517 37111
rect 10376 37080 10517 37108
rect 10376 37068 10382 37080
rect 10505 37077 10517 37080
rect 10551 37077 10563 37111
rect 12434 37108 12440 37120
rect 12395 37080 12440 37108
rect 10505 37071 10563 37077
rect 12434 37068 12440 37080
rect 12492 37068 12498 37120
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15657 37111 15715 37117
rect 15657 37108 15669 37111
rect 15528 37080 15669 37108
rect 15528 37068 15534 37080
rect 15657 37077 15669 37080
rect 15703 37077 15715 37111
rect 15657 37071 15715 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 16945 37111 17003 37117
rect 16945 37108 16957 37111
rect 16816 37080 16957 37108
rect 16816 37068 16822 37080
rect 16945 37077 16957 37080
rect 16991 37077 17003 37111
rect 16945 37071 17003 37077
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 19484 37080 19625 37108
rect 19484 37068 19490 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 19613 37071 19671 37077
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 22152 37080 22201 37108
rect 22152 37068 22158 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 23900 37080 24777 37108
rect 23900 37068 23906 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 25501 37071 25559 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30561 37111 30619 37117
rect 30561 37108 30573 37111
rect 30432 37080 30573 37108
rect 30432 37068 30438 37080
rect 30561 37077 30573 37080
rect 30607 37077 30619 37111
rect 30561 37071 30619 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 37366 37068 37372 37120
rect 37424 37108 37430 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 37424 37080 37657 37108
rect 37424 37068 37430 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 2685 36907 2743 36913
rect 2685 36873 2697 36907
rect 2731 36904 2743 36907
rect 2866 36904 2872 36916
rect 2731 36876 2872 36904
rect 2731 36873 2743 36876
rect 2685 36867 2743 36873
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 10686 36864 10692 36916
rect 10744 36904 10750 36916
rect 13541 36907 13599 36913
rect 13541 36904 13553 36907
rect 10744 36876 13553 36904
rect 10744 36864 10750 36876
rect 13541 36873 13553 36876
rect 13587 36873 13599 36907
rect 13541 36867 13599 36873
rect 14274 36864 14280 36916
rect 14332 36904 14338 36916
rect 15105 36907 15163 36913
rect 15105 36904 15117 36907
rect 14332 36876 15117 36904
rect 14332 36864 14338 36876
rect 15105 36873 15117 36876
rect 15151 36873 15163 36907
rect 20530 36904 20536 36916
rect 20491 36876 20536 36904
rect 15105 36867 15163 36873
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 21266 36904 21272 36916
rect 21227 36876 21272 36904
rect 21266 36864 21272 36876
rect 21324 36864 21330 36916
rect 1670 36768 1676 36780
rect 1631 36740 1676 36768
rect 1670 36728 1676 36740
rect 1728 36768 1734 36780
rect 3145 36771 3203 36777
rect 3145 36768 3157 36771
rect 1728 36740 3157 36768
rect 1728 36728 1734 36740
rect 3145 36737 3157 36740
rect 3191 36737 3203 36771
rect 3145 36731 3203 36737
rect 13725 36771 13783 36777
rect 13725 36737 13737 36771
rect 13771 36737 13783 36771
rect 13725 36731 13783 36737
rect 15289 36771 15347 36777
rect 15289 36737 15301 36771
rect 15335 36768 15347 36771
rect 19334 36768 19340 36780
rect 15335 36740 19340 36768
rect 15335 36737 15347 36740
rect 15289 36731 15347 36737
rect 13740 36700 13768 36731
rect 19334 36728 19340 36740
rect 19392 36728 19398 36780
rect 20548 36768 20576 36864
rect 22649 36839 22707 36845
rect 22649 36836 22661 36839
rect 22020 36808 22661 36836
rect 22020 36780 22048 36808
rect 22649 36805 22661 36808
rect 22695 36805 22707 36839
rect 22649 36799 22707 36805
rect 23014 36796 23020 36848
rect 23072 36836 23078 36848
rect 37553 36839 37611 36845
rect 23072 36808 26234 36836
rect 23072 36796 23078 36808
rect 21085 36771 21143 36777
rect 21085 36768 21097 36771
rect 20548 36740 21097 36768
rect 21085 36737 21097 36740
rect 21131 36737 21143 36771
rect 21085 36731 21143 36737
rect 21818 36728 21824 36780
rect 21876 36768 21882 36780
rect 22002 36768 22008 36780
rect 21876 36740 22008 36768
rect 21876 36728 21882 36740
rect 22002 36728 22008 36740
rect 22060 36728 22066 36780
rect 26206 36768 26234 36808
rect 37553 36805 37565 36839
rect 37599 36836 37611 36839
rect 38197 36839 38255 36845
rect 38197 36836 38209 36839
rect 37599 36808 38209 36836
rect 37599 36805 37611 36808
rect 37553 36799 37611 36805
rect 38197 36805 38209 36808
rect 38243 36836 38255 36839
rect 38654 36836 38660 36848
rect 38243 36808 38660 36836
rect 38243 36805 38255 36808
rect 38197 36799 38255 36805
rect 38654 36796 38660 36808
rect 38712 36796 38718 36848
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 22112 36740 25452 36768
rect 26206 36740 27169 36768
rect 14277 36703 14335 36709
rect 14277 36700 14289 36703
rect 13740 36672 14289 36700
rect 14277 36669 14289 36672
rect 14323 36700 14335 36703
rect 18782 36700 18788 36712
rect 14323 36672 18788 36700
rect 14323 36669 14335 36672
rect 14277 36663 14335 36669
rect 18782 36660 18788 36672
rect 18840 36700 18846 36712
rect 22112 36700 22140 36740
rect 18840 36672 22140 36700
rect 25225 36703 25283 36709
rect 18840 36660 18846 36672
rect 25225 36669 25237 36703
rect 25271 36700 25283 36703
rect 25314 36700 25320 36712
rect 25271 36672 25320 36700
rect 25271 36669 25283 36672
rect 25225 36663 25283 36669
rect 25314 36660 25320 36672
rect 25372 36660 25378 36712
rect 22189 36635 22247 36641
rect 22189 36601 22201 36635
rect 22235 36632 22247 36635
rect 25424 36632 25452 36740
rect 27157 36737 27169 36740
rect 27203 36768 27215 36771
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 27203 36740 27813 36768
rect 27203 36737 27215 36740
rect 27157 36731 27215 36737
rect 27801 36737 27813 36740
rect 27847 36737 27859 36771
rect 27801 36731 27859 36737
rect 35526 36700 35532 36712
rect 26206 36672 35532 36700
rect 26206 36632 26234 36672
rect 35526 36660 35532 36672
rect 35584 36660 35590 36712
rect 37458 36700 37464 36712
rect 35866 36672 37464 36700
rect 22235 36604 25268 36632
rect 25424 36604 26234 36632
rect 27341 36635 27399 36641
rect 22235 36601 22247 36604
rect 22189 36595 22247 36601
rect 1762 36564 1768 36576
rect 1723 36536 1768 36564
rect 1762 36524 1768 36536
rect 1820 36524 1826 36576
rect 25240 36564 25268 36604
rect 27341 36601 27353 36635
rect 27387 36632 27399 36635
rect 35866 36632 35894 36672
rect 37458 36660 37464 36672
rect 37516 36660 37522 36712
rect 27387 36604 35894 36632
rect 27387 36601 27399 36604
rect 27341 36595 27399 36601
rect 37918 36592 37924 36644
rect 37976 36632 37982 36644
rect 38013 36635 38071 36641
rect 38013 36632 38025 36635
rect 37976 36604 38025 36632
rect 37976 36592 37982 36604
rect 38013 36601 38025 36604
rect 38059 36601 38071 36635
rect 38013 36595 38071 36601
rect 29730 36564 29736 36576
rect 25240 36536 29736 36564
rect 29730 36524 29736 36536
rect 29788 36524 29794 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 14 36320 20 36372
rect 72 36360 78 36372
rect 1673 36363 1731 36369
rect 1673 36360 1685 36363
rect 72 36332 1685 36360
rect 72 36320 78 36332
rect 1673 36329 1685 36332
rect 1719 36329 1731 36363
rect 1673 36323 1731 36329
rect 1762 36320 1768 36372
rect 1820 36360 1826 36372
rect 13814 36360 13820 36372
rect 1820 36332 13820 36360
rect 1820 36320 1826 36332
rect 13814 36320 13820 36332
rect 13872 36320 13878 36372
rect 38194 36360 38200 36372
rect 38155 36332 38200 36360
rect 38194 36320 38200 36332
rect 38252 36320 38258 36372
rect 1946 36252 1952 36304
rect 2004 36292 2010 36304
rect 2317 36295 2375 36301
rect 2317 36292 2329 36295
rect 2004 36264 2329 36292
rect 2004 36252 2010 36264
rect 2317 36261 2329 36264
rect 2363 36261 2375 36295
rect 2317 36255 2375 36261
rect 1857 36159 1915 36165
rect 1857 36125 1869 36159
rect 1903 36156 1915 36159
rect 5442 36156 5448 36168
rect 1903 36128 5448 36156
rect 1903 36125 1915 36128
rect 1857 36119 1915 36125
rect 5442 36116 5448 36128
rect 5500 36116 5506 36168
rect 37553 36159 37611 36165
rect 37553 36125 37565 36159
rect 37599 36156 37611 36159
rect 37734 36156 37740 36168
rect 37599 36128 37740 36156
rect 37599 36125 37611 36128
rect 37553 36119 37611 36125
rect 37734 36116 37740 36128
rect 37792 36156 37798 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37792 36128 38025 36156
rect 37792 36116 37798 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 19426 35816 19432 35828
rect 18748 35788 19432 35816
rect 18748 35776 18754 35788
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37476 35652 38025 35680
rect 27890 35436 27896 35488
rect 27948 35476 27954 35488
rect 37476 35485 37504 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 37461 35479 37519 35485
rect 37461 35476 37473 35479
rect 27948 35448 37473 35476
rect 27948 35436 27954 35448
rect 37461 35445 37473 35448
rect 37507 35445 37519 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 37461 35439 37519 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 18414 34184 18420 34196
rect 18375 34156 18420 34184
rect 18414 34144 18420 34156
rect 18472 34144 18478 34196
rect 18233 33983 18291 33989
rect 18233 33980 18245 33983
rect 17696 33952 18245 33980
rect 17696 33856 17724 33952
rect 18233 33949 18245 33952
rect 18279 33949 18291 33983
rect 18233 33943 18291 33949
rect 17678 33844 17684 33856
rect 17639 33816 17684 33844
rect 17678 33804 17684 33816
rect 17736 33804 17742 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1670 33504 1676 33516
rect 1631 33476 1676 33504
rect 1670 33464 1676 33476
rect 1728 33464 1734 33516
rect 37553 33507 37611 33513
rect 37553 33473 37565 33507
rect 37599 33504 37611 33507
rect 38194 33504 38200 33516
rect 37599 33476 38200 33504
rect 37599 33473 37611 33476
rect 37553 33467 37611 33473
rect 38194 33464 38200 33476
rect 38252 33464 38258 33516
rect 1857 33371 1915 33377
rect 1857 33337 1869 33371
rect 1903 33368 1915 33371
rect 9306 33368 9312 33380
rect 1903 33340 9312 33368
rect 1903 33337 1915 33340
rect 1857 33331 1915 33337
rect 9306 33328 9312 33340
rect 9364 33328 9370 33380
rect 38013 33371 38071 33377
rect 38013 33368 38025 33371
rect 26206 33340 38025 33368
rect 26206 33312 26234 33340
rect 38013 33337 38025 33340
rect 38059 33337 38071 33371
rect 38013 33331 38071 33337
rect 26142 33260 26148 33312
rect 26200 33272 26234 33312
rect 26200 33260 26206 33272
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1670 33096 1676 33108
rect 1631 33068 1676 33096
rect 1670 33056 1676 33068
rect 1728 33056 1734 33108
rect 5169 33099 5227 33105
rect 5169 33065 5181 33099
rect 5215 33096 5227 33099
rect 5258 33096 5264 33108
rect 5215 33068 5264 33096
rect 5215 33065 5227 33068
rect 5169 33059 5227 33065
rect 5258 33056 5264 33068
rect 5316 33056 5322 33108
rect 4985 32895 5043 32901
rect 4985 32861 4997 32895
rect 5031 32861 5043 32895
rect 4985 32855 5043 32861
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32892 9919 32895
rect 9907 32864 10456 32892
rect 9907 32861 9919 32864
rect 9861 32855 9919 32861
rect 5000 32756 5028 32855
rect 5442 32784 5448 32836
rect 5500 32824 5506 32836
rect 5500 32796 9720 32824
rect 5500 32784 5506 32796
rect 5721 32759 5779 32765
rect 5721 32756 5733 32759
rect 5000 32728 5733 32756
rect 5721 32725 5733 32728
rect 5767 32756 5779 32759
rect 9214 32756 9220 32768
rect 5767 32728 9220 32756
rect 5767 32725 5779 32728
rect 5721 32719 5779 32725
rect 9214 32716 9220 32728
rect 9272 32716 9278 32768
rect 9692 32765 9720 32796
rect 10428 32765 10456 32864
rect 9677 32759 9735 32765
rect 9677 32725 9689 32759
rect 9723 32725 9735 32759
rect 9677 32719 9735 32725
rect 10413 32759 10471 32765
rect 10413 32725 10425 32759
rect 10459 32756 10471 32759
rect 25498 32756 25504 32768
rect 10459 32728 25504 32756
rect 10459 32725 10471 32728
rect 10413 32719 10471 32725
rect 25498 32716 25504 32728
rect 25556 32716 25562 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 38013 32419 38071 32425
rect 22235 32388 22784 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 15838 32172 15844 32224
rect 15896 32212 15902 32224
rect 22756 32221 22784 32388
rect 38013 32385 38025 32419
rect 38059 32416 38071 32419
rect 38102 32416 38108 32428
rect 38059 32388 38108 32416
rect 38059 32385 38071 32388
rect 38013 32379 38071 32385
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 15896 32184 22017 32212
rect 15896 32172 15902 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 22005 32175 22063 32181
rect 22741 32215 22799 32221
rect 22741 32181 22753 32215
rect 22787 32212 22799 32215
rect 28626 32212 28632 32224
rect 22787 32184 28632 32212
rect 22787 32181 22799 32184
rect 22741 32175 22799 32181
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 9490 31968 9496 32020
rect 9548 32008 9554 32020
rect 9861 32011 9919 32017
rect 9861 32008 9873 32011
rect 9548 31980 9873 32008
rect 9548 31968 9554 31980
rect 9861 31977 9873 31980
rect 9907 31977 9919 32011
rect 9861 31971 9919 31977
rect 1765 31943 1823 31949
rect 1765 31909 1777 31943
rect 1811 31940 1823 31943
rect 1811 31912 16574 31940
rect 1811 31909 1823 31912
rect 1765 31903 1823 31909
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 9953 31807 10011 31813
rect 9953 31773 9965 31807
rect 9999 31804 10011 31807
rect 10502 31804 10508 31816
rect 9999 31776 10508 31804
rect 9999 31773 10011 31776
rect 9953 31767 10011 31773
rect 10502 31764 10508 31776
rect 10560 31764 10566 31816
rect 16546 31804 16574 31912
rect 30098 31804 30104 31816
rect 16546 31776 30104 31804
rect 30098 31764 30104 31776
rect 30156 31764 30162 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1578 31396 1584 31408
rect 1539 31368 1584 31396
rect 1578 31356 1584 31368
rect 1636 31356 1642 31408
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 30285 30855 30343 30861
rect 30285 30821 30297 30855
rect 30331 30852 30343 30855
rect 38010 30852 38016 30864
rect 30331 30824 38016 30852
rect 30331 30821 30343 30824
rect 30285 30815 30343 30821
rect 38010 30812 38016 30824
rect 38068 30812 38074 30864
rect 30098 30716 30104 30728
rect 30059 30688 30104 30716
rect 30098 30676 30104 30688
rect 30156 30716 30162 30728
rect 30745 30719 30803 30725
rect 30745 30716 30757 30719
rect 30156 30688 30757 30716
rect 30156 30676 30162 30688
rect 30745 30685 30757 30688
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 19334 30200 19340 30252
rect 19392 30240 19398 30252
rect 19521 30243 19579 30249
rect 19521 30240 19533 30243
rect 19392 30212 19533 30240
rect 19392 30200 19398 30212
rect 19521 30209 19533 30212
rect 19567 30209 19579 30243
rect 38010 30240 38016 30252
rect 37971 30212 38016 30240
rect 19521 30203 19579 30209
rect 38010 30200 38016 30212
rect 38068 30200 38074 30252
rect 1578 30172 1584 30184
rect 1539 30144 1584 30172
rect 1578 30132 1584 30144
rect 1636 30132 1642 30184
rect 1857 30175 1915 30181
rect 1857 30141 1869 30175
rect 1903 30172 1915 30175
rect 2498 30172 2504 30184
rect 1903 30144 2504 30172
rect 1903 30141 1915 30144
rect 1857 30135 1915 30141
rect 2498 30132 2504 30144
rect 2556 30132 2562 30184
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19429 30039 19487 30045
rect 19429 30036 19441 30039
rect 19392 30008 19441 30036
rect 19392 29996 19398 30008
rect 19429 30005 19441 30008
rect 19475 30005 19487 30039
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 19429 29999 19487 30005
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 20533 29291 20591 29297
rect 20533 29257 20545 29291
rect 20579 29288 20591 29291
rect 24578 29288 24584 29300
rect 20579 29260 24584 29288
rect 20579 29257 20591 29260
rect 20533 29251 20591 29257
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 30742 29248 30748 29300
rect 30800 29288 30806 29300
rect 30837 29291 30895 29297
rect 30837 29288 30849 29291
rect 30800 29260 30849 29288
rect 30800 29248 30806 29260
rect 30837 29257 30849 29260
rect 30883 29257 30895 29291
rect 30837 29251 30895 29257
rect 12066 29112 12072 29164
rect 12124 29152 12130 29164
rect 20349 29155 20407 29161
rect 20349 29152 20361 29155
rect 12124 29124 20361 29152
rect 12124 29112 12130 29124
rect 20349 29121 20361 29124
rect 20395 29152 20407 29155
rect 20993 29155 21051 29161
rect 20993 29152 21005 29155
rect 20395 29124 21005 29152
rect 20395 29121 20407 29124
rect 20349 29115 20407 29121
rect 20993 29121 21005 29124
rect 21039 29121 21051 29155
rect 30926 29152 30932 29164
rect 30887 29124 30932 29152
rect 20993 29115 21051 29121
rect 30926 29112 30932 29124
rect 30984 29152 30990 29164
rect 31389 29155 31447 29161
rect 31389 29152 31401 29155
rect 30984 29124 31401 29152
rect 30984 29112 30990 29124
rect 31389 29121 31401 29124
rect 31435 29121 31447 29155
rect 31389 29115 31447 29121
rect 34146 29112 34152 29164
rect 34204 29152 34210 29164
rect 38013 29155 38071 29161
rect 38013 29152 38025 29155
rect 34204 29124 38025 29152
rect 34204 29112 34210 29124
rect 38013 29121 38025 29124
rect 38059 29121 38071 29155
rect 38013 29115 38071 29121
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 30650 28200 30656 28212
rect 30611 28172 30656 28200
rect 30650 28160 30656 28172
rect 30708 28160 30714 28212
rect 1854 28064 1860 28076
rect 1815 28036 1860 28064
rect 1854 28024 1860 28036
rect 1912 28024 1918 28076
rect 30561 28067 30619 28073
rect 30561 28033 30573 28067
rect 30607 28064 30619 28067
rect 31202 28064 31208 28076
rect 30607 28036 31208 28064
rect 30607 28033 30619 28036
rect 30561 28027 30619 28033
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 31202 27860 31208 27872
rect 31163 27832 31208 27860
rect 31202 27820 31208 27832
rect 31260 27820 31266 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 23014 27588 23020 27600
rect 22975 27560 23020 27588
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27452 22615 27455
rect 23032 27452 23060 27548
rect 22603 27424 23060 27452
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 22094 27276 22100 27328
rect 22152 27316 22158 27328
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 22152 27288 22477 27316
rect 22152 27276 22158 27288
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 38286 27316 38292 27328
rect 38247 27288 38292 27316
rect 22465 27279 22523 27285
rect 38286 27276 38292 27288
rect 38344 27276 38350 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 18782 27112 18788 27124
rect 18743 27084 18788 27112
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 6822 26976 6828 26988
rect 1903 26948 6828 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 15381 26979 15439 26985
rect 15381 26945 15393 26979
rect 15427 26976 15439 26979
rect 16025 26979 16083 26985
rect 16025 26976 16037 26979
rect 15427 26948 16037 26976
rect 15427 26945 15439 26948
rect 15381 26939 15439 26945
rect 16025 26945 16037 26948
rect 16071 26976 16083 26979
rect 18233 26979 18291 26985
rect 16071 26948 16574 26976
rect 16071 26945 16083 26948
rect 16025 26939 16083 26945
rect 16546 26908 16574 26948
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18800 26976 18828 27072
rect 18279 26948 18828 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 20530 26908 20536 26920
rect 16546 26880 20536 26908
rect 20530 26868 20536 26880
rect 20588 26868 20594 26920
rect 37366 26868 37372 26920
rect 37424 26908 37430 26920
rect 38013 26911 38071 26917
rect 38013 26908 38025 26911
rect 37424 26880 38025 26908
rect 37424 26868 37430 26880
rect 38013 26877 38025 26880
rect 38059 26877 38071 26911
rect 38286 26908 38292 26920
rect 38247 26880 38292 26908
rect 38013 26871 38071 26877
rect 38286 26868 38292 26880
rect 38344 26868 38350 26920
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 15654 26732 15660 26784
rect 15712 26772 15718 26784
rect 15933 26775 15991 26781
rect 15933 26772 15945 26775
rect 15712 26744 15945 26772
rect 15712 26732 15718 26744
rect 15933 26741 15945 26744
rect 15979 26741 15991 26775
rect 15933 26735 15991 26741
rect 18141 26775 18199 26781
rect 18141 26741 18153 26775
rect 18187 26772 18199 26775
rect 18322 26772 18328 26784
rect 18187 26744 18328 26772
rect 18187 26741 18199 26744
rect 18141 26735 18199 26741
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 9398 26528 9404 26580
rect 9456 26568 9462 26580
rect 14369 26571 14427 26577
rect 14369 26568 14381 26571
rect 9456 26540 14381 26568
rect 9456 26528 9462 26540
rect 14369 26537 14381 26540
rect 14415 26537 14427 26571
rect 14369 26531 14427 26537
rect 20441 26571 20499 26577
rect 20441 26537 20453 26571
rect 20487 26568 20499 26571
rect 22002 26568 22008 26580
rect 20487 26540 22008 26568
rect 20487 26537 20499 26540
rect 20441 26531 20499 26537
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26364 14519 26367
rect 19889 26367 19947 26373
rect 14507 26336 15056 26364
rect 14507 26333 14519 26336
rect 14461 26327 14519 26333
rect 15028 26305 15056 26336
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 20456 26364 20484 26531
rect 22002 26528 22008 26540
rect 22060 26528 22066 26580
rect 36906 26528 36912 26580
rect 36964 26568 36970 26580
rect 37829 26571 37887 26577
rect 37829 26568 37841 26571
rect 36964 26540 37841 26568
rect 36964 26528 36970 26540
rect 37829 26537 37841 26540
rect 37875 26537 37887 26571
rect 37829 26531 37887 26537
rect 38010 26364 38016 26376
rect 19935 26336 20484 26364
rect 37971 26336 38016 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 38010 26324 38016 26336
rect 38068 26324 38074 26376
rect 15013 26299 15071 26305
rect 15013 26265 15025 26299
rect 15059 26296 15071 26299
rect 18138 26296 18144 26308
rect 15059 26268 18144 26296
rect 15059 26265 15071 26268
rect 15013 26259 15071 26265
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 19797 26299 19855 26305
rect 19797 26265 19809 26299
rect 19843 26296 19855 26299
rect 20070 26296 20076 26308
rect 19843 26268 20076 26296
rect 19843 26265 19855 26268
rect 19797 26259 19855 26265
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 33594 26024 33600 26036
rect 33555 25996 33600 26024
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25888 33839 25891
rect 34238 25888 34244 25900
rect 33827 25860 34244 25888
rect 33827 25857 33839 25860
rect 33781 25851 33839 25857
rect 34238 25848 34244 25860
rect 34296 25848 34302 25900
rect 34238 25684 34244 25696
rect 34199 25656 34244 25684
rect 34238 25644 34244 25656
rect 34296 25644 34302 25696
rect 38010 25644 38016 25696
rect 38068 25684 38074 25696
rect 38105 25687 38163 25693
rect 38105 25684 38117 25687
rect 38068 25656 38117 25684
rect 38068 25644 38074 25656
rect 38105 25653 38117 25656
rect 38151 25653 38163 25687
rect 38105 25647 38163 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 38013 25483 38071 25489
rect 38013 25449 38025 25483
rect 38059 25480 38071 25483
rect 38194 25480 38200 25492
rect 38059 25452 38200 25480
rect 38059 25449 38071 25452
rect 38013 25443 38071 25449
rect 38194 25440 38200 25452
rect 38252 25440 38258 25492
rect 37826 25276 37832 25288
rect 37787 25248 37832 25276
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 37458 24896 37464 24948
rect 37516 24936 37522 24948
rect 38010 24936 38016 24948
rect 37516 24908 38016 24936
rect 37516 24896 37522 24908
rect 38010 24896 38016 24908
rect 38068 24896 38074 24948
rect 25498 24828 25504 24880
rect 25556 24868 25562 24880
rect 26694 24868 26700 24880
rect 25556 24840 26700 24868
rect 25556 24828 25562 24840
rect 26694 24828 26700 24840
rect 26752 24828 26758 24880
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 20809 24803 20867 24809
rect 1903 24772 2452 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2424 24673 2452 24772
rect 20809 24769 20821 24803
rect 20855 24800 20867 24803
rect 21361 24803 21419 24809
rect 21361 24800 21373 24803
rect 20855 24772 21373 24800
rect 20855 24769 20867 24772
rect 20809 24763 20867 24769
rect 21361 24769 21373 24772
rect 21407 24800 21419 24803
rect 21634 24800 21640 24812
rect 21407 24772 21640 24800
rect 21407 24769 21419 24772
rect 21361 24763 21419 24769
rect 21634 24760 21640 24772
rect 21692 24800 21698 24812
rect 37918 24800 37924 24812
rect 21692 24772 37924 24800
rect 21692 24760 21698 24772
rect 37918 24760 37924 24772
rect 37976 24760 37982 24812
rect 38013 24803 38071 24809
rect 38013 24769 38025 24803
rect 38059 24800 38071 24803
rect 38102 24800 38108 24812
rect 38059 24772 38108 24800
rect 38059 24769 38071 24772
rect 38013 24763 38071 24769
rect 38102 24760 38108 24772
rect 38160 24760 38166 24812
rect 2409 24667 2467 24673
rect 2409 24633 2421 24667
rect 2455 24664 2467 24667
rect 20625 24667 20683 24673
rect 20625 24664 20637 24667
rect 2455 24636 20637 24664
rect 2455 24633 2467 24636
rect 2409 24627 2467 24633
rect 20625 24633 20637 24636
rect 20671 24633 20683 24667
rect 20625 24627 20683 24633
rect 1670 24596 1676 24608
rect 1631 24568 1676 24596
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 25222 24392 25228 24404
rect 25183 24364 25228 24392
rect 25222 24352 25228 24364
rect 25280 24352 25286 24404
rect 34146 24392 34152 24404
rect 34107 24364 34152 24392
rect 34146 24352 34152 24364
rect 34204 24352 34210 24404
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 25004 24160 25053 24188
rect 25004 24148 25010 24160
rect 25041 24157 25053 24160
rect 25087 24188 25099 24191
rect 25685 24191 25743 24197
rect 25685 24188 25697 24191
rect 25087 24160 25697 24188
rect 25087 24157 25099 24160
rect 25041 24151 25099 24157
rect 25685 24157 25697 24160
rect 25731 24157 25743 24191
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 25685 24151 25743 24157
rect 33428 24160 33977 24188
rect 33428 24064 33456 24160
rect 33965 24157 33977 24160
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 33410 24052 33416 24064
rect 33371 24024 33416 24052
rect 33410 24012 33416 24024
rect 33468 24012 33474 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 38010 23712 38016 23724
rect 37971 23684 38016 23712
rect 38010 23672 38016 23684
rect 38068 23672 38074 23724
rect 38194 23508 38200 23520
rect 38155 23480 38200 23508
rect 38194 23468 38200 23480
rect 38252 23468 38258 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1765 23307 1823 23313
rect 1765 23273 1777 23307
rect 1811 23304 1823 23307
rect 1854 23304 1860 23316
rect 1811 23276 1860 23304
rect 1811 23273 1823 23276
rect 1765 23267 1823 23273
rect 1854 23264 1860 23276
rect 1912 23264 1918 23316
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23100 2007 23103
rect 1995 23072 2452 23100
rect 1995 23069 2007 23072
rect 1949 23063 2007 23069
rect 2424 22976 2452 23072
rect 2406 22964 2412 22976
rect 2367 22936 2412 22964
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 37921 22763 37979 22769
rect 37921 22729 37933 22763
rect 37967 22760 37979 22763
rect 38010 22760 38016 22772
rect 37967 22732 38016 22760
rect 37967 22729 37979 22732
rect 37921 22723 37979 22729
rect 38010 22720 38016 22732
rect 38068 22720 38074 22772
rect 1762 22584 1768 22636
rect 1820 22624 1826 22636
rect 1857 22627 1915 22633
rect 1857 22624 1869 22627
rect 1820 22596 1869 22624
rect 1820 22584 1826 22596
rect 1857 22593 1869 22596
rect 1903 22593 1915 22627
rect 1857 22587 1915 22593
rect 37274 22584 37280 22636
rect 37332 22624 37338 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37332 22596 37841 22624
rect 37332 22584 37338 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 1670 22488 1676 22500
rect 1631 22460 1676 22488
rect 1670 22448 1676 22460
rect 1728 22448 1734 22500
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7883 21984 8432 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 8404 21885 8432 21984
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 6880 21848 7665 21876
rect 6880 21836 6886 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 8389 21879 8447 21885
rect 8389 21845 8401 21879
rect 8435 21876 8447 21879
rect 9858 21876 9864 21888
rect 8435 21848 9864 21876
rect 8435 21845 8447 21848
rect 8389 21839 8447 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 37274 21836 37280 21888
rect 37332 21876 37338 21888
rect 37645 21879 37703 21885
rect 37645 21876 37657 21879
rect 37332 21848 37657 21876
rect 37332 21836 37338 21848
rect 37645 21845 37657 21848
rect 37691 21845 37703 21879
rect 37645 21839 37703 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1578 21496 1584 21548
rect 1636 21536 1642 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1636 21508 1685 21536
rect 1636 21496 1642 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 1673 21499 1731 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 1854 21400 1860 21412
rect 1815 21372 1860 21400
rect 1854 21360 1860 21372
rect 1912 21360 1918 21412
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 38013 21131 38071 21137
rect 38013 21097 38025 21131
rect 38059 21128 38071 21131
rect 38102 21128 38108 21140
rect 38059 21100 38108 21128
rect 38059 21097 38071 21100
rect 38013 21091 38071 21097
rect 38102 21088 38108 21100
rect 38160 21088 38166 21140
rect 37829 20927 37887 20933
rect 37829 20893 37841 20927
rect 37875 20924 37887 20927
rect 38102 20924 38108 20936
rect 37875 20896 38108 20924
rect 37875 20893 37887 20896
rect 37829 20887 37887 20893
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1854 20408 1860 20460
rect 1912 20448 1918 20460
rect 20349 20451 20407 20457
rect 20349 20448 20361 20451
rect 1912 20420 20361 20448
rect 1912 20408 1918 20420
rect 20349 20417 20361 20420
rect 20395 20448 20407 20451
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20395 20420 20821 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 20254 20244 20260 20256
rect 20215 20216 20260 20244
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 20824 20244 20852 20411
rect 33410 20244 33416 20256
rect 20824 20216 33416 20244
rect 33410 20204 33416 20216
rect 33468 20204 33474 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 27890 20040 27896 20052
rect 27851 20012 27896 20040
rect 27890 20000 27896 20012
rect 27948 20000 27954 20052
rect 37645 19839 37703 19845
rect 37645 19805 37657 19839
rect 37691 19836 37703 19839
rect 38286 19836 38292 19848
rect 37691 19808 38292 19836
rect 37691 19805 37703 19808
rect 37645 19799 37703 19805
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 27249 19771 27307 19777
rect 27249 19737 27261 19771
rect 27295 19768 27307 19771
rect 27801 19771 27859 19777
rect 27801 19768 27813 19771
rect 27295 19740 27813 19768
rect 27295 19737 27307 19740
rect 27249 19731 27307 19737
rect 27801 19737 27813 19740
rect 27847 19768 27859 19771
rect 29270 19768 29276 19780
rect 27847 19740 29276 19768
rect 27847 19737 27859 19740
rect 27801 19731 27859 19737
rect 29270 19728 29276 19740
rect 29328 19728 29334 19780
rect 38102 19700 38108 19712
rect 38063 19672 38108 19700
rect 38102 19660 38108 19672
rect 38160 19660 38166 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 1946 19360 1952 19372
rect 1903 19332 1952 19360
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 26142 18952 26148 18964
rect 26103 18924 26148 18952
rect 26142 18912 26148 18924
rect 26200 18912 26206 18964
rect 25682 18748 25688 18760
rect 25595 18720 25688 18748
rect 25682 18708 25688 18720
rect 25740 18748 25746 18760
rect 26142 18748 26148 18760
rect 25740 18720 26148 18748
rect 25740 18708 25746 18720
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18748 33195 18751
rect 38102 18748 38108 18760
rect 33183 18720 38108 18748
rect 33183 18717 33195 18720
rect 33137 18711 33195 18717
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 25590 18612 25596 18624
rect 25551 18584 25596 18612
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 33042 18612 33048 18624
rect 33003 18584 33048 18612
rect 33042 18572 33048 18584
rect 33100 18572 33106 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 18509 18343 18567 18349
rect 18509 18309 18521 18343
rect 18555 18340 18567 18343
rect 19426 18340 19432 18352
rect 18555 18312 19432 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19392 18244 19625 18272
rect 19392 18232 19398 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20073 18275 20131 18281
rect 20073 18241 20085 18275
rect 20119 18272 20131 18275
rect 20119 18244 20852 18272
rect 20119 18241 20131 18244
rect 20073 18235 20131 18241
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 19352 18176 19441 18204
rect 19352 18148 19380 18176
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 19334 18096 19340 18148
rect 19392 18096 19398 18148
rect 20824 18145 20852 18244
rect 24854 18204 24860 18216
rect 24815 18176 24860 18204
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 33042 18204 33048 18216
rect 25087 18176 33048 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 33042 18164 33048 18176
rect 33100 18164 33106 18216
rect 20809 18139 20867 18145
rect 20809 18105 20821 18139
rect 20855 18136 20867 18139
rect 30098 18136 30104 18148
rect 20855 18108 30104 18136
rect 20855 18105 20867 18108
rect 20809 18099 20867 18105
rect 30098 18096 30104 18108
rect 30156 18096 30162 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 19242 18068 19248 18080
rect 19203 18040 19248 18068
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 24673 18071 24731 18077
rect 24673 18037 24685 18071
rect 24719 18068 24731 18071
rect 25130 18068 25136 18080
rect 24719 18040 25136 18068
rect 24719 18037 24731 18040
rect 24673 18031 24731 18037
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 19242 17824 19248 17876
rect 19300 17864 19306 17876
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 19300 17836 19809 17864
rect 19300 17824 19306 17836
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 21634 17864 21640 17876
rect 21595 17836 21640 17864
rect 19797 17827 19855 17833
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 25682 17864 25688 17876
rect 25643 17836 25688 17864
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 23017 17799 23075 17805
rect 23017 17765 23029 17799
rect 23063 17796 23075 17799
rect 23934 17796 23940 17808
rect 23063 17768 23940 17796
rect 23063 17765 23075 17768
rect 23017 17759 23075 17765
rect 23934 17756 23940 17768
rect 23992 17756 23998 17808
rect 19426 17728 19432 17740
rect 19387 17700 19432 17728
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 22094 17688 22100 17740
rect 22152 17728 22158 17740
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 22152 17700 22385 17728
rect 22152 17688 22158 17700
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 25700 17728 25728 17824
rect 22373 17691 22431 17697
rect 23952 17700 25728 17728
rect 19518 17620 19524 17672
rect 19576 17660 19582 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 19576 17632 19625 17660
rect 19576 17620 19582 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17660 22615 17663
rect 23198 17660 23204 17672
rect 22603 17632 23204 17660
rect 22603 17629 22615 17632
rect 22557 17623 22615 17629
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 23952 17669 23980 17700
rect 23937 17663 23995 17669
rect 23937 17629 23949 17663
rect 23983 17629 23995 17663
rect 24578 17660 24584 17672
rect 24539 17632 24584 17660
rect 23937 17623 23995 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 23658 17592 23664 17604
rect 22066 17564 23664 17592
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 22066 17524 22094 17564
rect 23658 17552 23664 17564
rect 23716 17552 23722 17604
rect 18196 17496 22094 17524
rect 18196 17484 18202 17496
rect 23106 17484 23112 17536
rect 23164 17524 23170 17536
rect 23845 17527 23903 17533
rect 23845 17524 23857 17527
rect 23164 17496 23857 17524
rect 23164 17484 23170 17496
rect 23845 17493 23857 17496
rect 23891 17493 23903 17527
rect 23845 17487 23903 17493
rect 25130 17484 25136 17536
rect 25188 17524 25194 17536
rect 25225 17527 25283 17533
rect 25225 17524 25237 17527
rect 25188 17496 25237 17524
rect 25188 17484 25194 17496
rect 25225 17493 25237 17496
rect 25271 17493 25283 17527
rect 25225 17487 25283 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 23106 17320 23112 17332
rect 3476 17292 23112 17320
rect 3476 17280 3482 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23860 17292 24624 17320
rect 18598 17252 18604 17264
rect 18559 17224 18604 17252
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 18693 17255 18751 17261
rect 18693 17221 18705 17255
rect 18739 17252 18751 17255
rect 19242 17252 19248 17264
rect 18739 17224 19248 17252
rect 18739 17221 18751 17224
rect 18693 17215 18751 17221
rect 19242 17212 19248 17224
rect 19300 17212 19306 17264
rect 22189 17255 22247 17261
rect 22189 17221 22201 17255
rect 22235 17252 22247 17255
rect 22278 17252 22284 17264
rect 22235 17224 22284 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 23860 17261 23888 17292
rect 23845 17255 23903 17261
rect 23845 17221 23857 17255
rect 23891 17221 23903 17255
rect 23845 17215 23903 17221
rect 23934 17212 23940 17264
rect 23992 17252 23998 17264
rect 23992 17224 24037 17252
rect 23992 17212 23998 17224
rect 16206 17184 16212 17196
rect 16167 17156 16212 17184
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17310 17184 17316 17196
rect 17083 17156 17316 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17184 21511 17187
rect 21634 17184 21640 17196
rect 21499 17156 21640 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 14826 17116 14832 17128
rect 14787 17088 14832 17116
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 19245 17119 19303 17125
rect 19245 17116 19257 17119
rect 15528 17088 19257 17116
rect 15528 17076 15534 17088
rect 19245 17085 19257 17088
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17116 19487 17119
rect 20806 17116 20812 17128
rect 19475 17088 20812 17116
rect 19475 17085 19487 17088
rect 19429 17079 19487 17085
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22373 17119 22431 17125
rect 22152 17088 22197 17116
rect 22152 17076 22158 17088
rect 22373 17085 22385 17119
rect 22419 17085 22431 17119
rect 23658 17116 23664 17128
rect 23619 17088 23664 17116
rect 22373 17079 22431 17085
rect 18138 17048 18144 17060
rect 18099 17020 18144 17048
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 21726 17008 21732 17060
rect 21784 17048 21790 17060
rect 22388 17048 22416 17079
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 24596 17116 24624 17292
rect 24946 17280 24952 17332
rect 25004 17320 25010 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 25004 17292 25145 17320
rect 25004 17280 25010 17292
rect 25133 17289 25145 17292
rect 25179 17289 25191 17323
rect 25133 17283 25191 17289
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17184 24731 17187
rect 24964 17184 24992 17280
rect 24719 17156 24992 17184
rect 24719 17153 24731 17156
rect 24673 17147 24731 17153
rect 25866 17116 25872 17128
rect 24596 17088 25872 17116
rect 25866 17076 25872 17088
rect 25924 17076 25930 17128
rect 32950 17116 32956 17128
rect 28966 17088 32956 17116
rect 21784 17020 22416 17048
rect 21784 17008 21790 17020
rect 23106 17008 23112 17060
rect 23164 17048 23170 17060
rect 28966 17048 28994 17088
rect 32950 17076 32956 17088
rect 33008 17076 33014 17128
rect 23164 17020 28994 17048
rect 23164 17008 23170 17020
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 15436 16952 15485 16980
rect 15436 16940 15442 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 16080 16952 16129 16980
rect 16080 16940 16086 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16632 16952 16957 16980
rect 16632 16940 16638 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19300 16952 19625 16980
rect 19300 16940 19306 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 21361 16983 21419 16989
rect 21361 16949 21373 16983
rect 21407 16980 21419 16983
rect 21450 16980 21456 16992
rect 21407 16952 21456 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 24578 16980 24584 16992
rect 22428 16952 24584 16980
rect 22428 16940 22434 16952
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2096 16748 6914 16776
rect 2096 16736 2102 16748
rect 6886 16708 6914 16748
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 17586 16776 17592 16788
rect 14332 16748 17592 16776
rect 14332 16736 14338 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 19484 16748 19533 16776
rect 19484 16736 19490 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 24946 16776 24952 16788
rect 19521 16739 19579 16745
rect 22066 16748 24952 16776
rect 22066 16708 22094 16748
rect 24946 16736 24952 16748
rect 25004 16736 25010 16788
rect 6886 16680 22094 16708
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 24673 16711 24731 16717
rect 24673 16708 24685 16711
rect 23716 16680 24685 16708
rect 23716 16668 23722 16680
rect 24673 16677 24685 16680
rect 24719 16677 24731 16711
rect 24673 16671 24731 16677
rect 14826 16640 14832 16652
rect 14787 16612 14832 16640
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 15562 16640 15568 16652
rect 15519 16612 15568 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 22094 16640 22100 16652
rect 16264 16612 18736 16640
rect 16264 16600 16270 16612
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 18708 16581 18736 16612
rect 19444 16612 22100 16640
rect 19444 16581 19472 16612
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 22370 16640 22376 16652
rect 22331 16612 22376 16640
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23106 16640 23112 16652
rect 23067 16612 23112 16640
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 25130 16640 25136 16652
rect 23768 16612 25136 16640
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17368 16544 17417 16572
rect 17368 16532 17374 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 23290 16572 23296 16584
rect 23251 16544 23296 16572
rect 19429 16535 19487 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23768 16581 23796 16612
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 23753 16575 23811 16581
rect 23753 16541 23765 16575
rect 23799 16541 23811 16575
rect 23753 16535 23811 16541
rect 13630 16464 13636 16516
rect 13688 16504 13694 16516
rect 14921 16507 14979 16513
rect 14921 16504 14933 16507
rect 13688 16476 14933 16504
rect 13688 16464 13694 16476
rect 14921 16473 14933 16476
rect 14967 16473 14979 16507
rect 16114 16504 16120 16516
rect 16075 16476 16120 16504
rect 14921 16467 14979 16473
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 16574 16504 16580 16516
rect 16255 16476 16580 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 16758 16504 16764 16516
rect 16719 16476 16764 16504
rect 16758 16464 16764 16476
rect 16816 16464 16822 16516
rect 18141 16507 18199 16513
rect 18141 16504 18153 16507
rect 16868 16476 18153 16504
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 16868 16436 16896 16476
rect 18141 16473 18153 16476
rect 18187 16504 18199 16507
rect 18414 16504 18420 16516
rect 18187 16476 18420 16504
rect 18187 16473 18199 16476
rect 18141 16467 18199 16473
rect 18414 16464 18420 16476
rect 18472 16464 18478 16516
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21726 16504 21732 16516
rect 21324 16476 21732 16504
rect 21324 16464 21330 16476
rect 21726 16464 21732 16476
rect 21784 16464 21790 16516
rect 21910 16464 21916 16516
rect 21968 16504 21974 16516
rect 22281 16507 22339 16513
rect 22281 16504 22293 16507
rect 21968 16476 22293 16504
rect 21968 16464 21974 16476
rect 22281 16473 22293 16476
rect 22327 16473 22339 16507
rect 22281 16467 22339 16473
rect 24946 16464 24952 16516
rect 25004 16504 25010 16516
rect 25124 16507 25182 16513
rect 25124 16504 25136 16507
rect 25004 16476 25136 16504
rect 25004 16464 25010 16476
rect 25124 16473 25136 16476
rect 25170 16473 25182 16507
rect 25124 16467 25182 16473
rect 25222 16464 25228 16516
rect 25280 16504 25286 16516
rect 25280 16476 25325 16504
rect 25280 16464 25286 16476
rect 10928 16408 16896 16436
rect 10928 16396 10934 16408
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17313 16439 17371 16445
rect 17313 16436 17325 16439
rect 17276 16408 17325 16436
rect 17276 16396 17282 16408
rect 17313 16405 17325 16408
rect 17359 16405 17371 16439
rect 17313 16399 17371 16405
rect 18785 16439 18843 16445
rect 18785 16405 18797 16439
rect 18831 16436 18843 16439
rect 22186 16436 22192 16448
rect 18831 16408 22192 16436
rect 18831 16405 18843 16408
rect 18785 16399 18843 16405
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 16114 16232 16120 16244
rect 14476 16204 16120 16232
rect 14476 16173 14504 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 22557 16235 22615 16241
rect 16500 16204 22094 16232
rect 14461 16167 14519 16173
rect 14461 16164 14473 16167
rect 12406 16136 14473 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 4062 16096 4068 16108
rect 1903 16068 4068 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 12406 16028 12434 16136
rect 14461 16133 14473 16136
rect 14507 16133 14519 16167
rect 14461 16127 14519 16133
rect 14553 16167 14611 16173
rect 14553 16133 14565 16167
rect 14599 16164 14611 16167
rect 14642 16164 14648 16176
rect 14599 16136 14648 16164
rect 14599 16133 14611 16136
rect 14553 16127 14611 16133
rect 14642 16124 14648 16136
rect 14700 16124 14706 16176
rect 15746 16164 15752 16176
rect 15707 16136 15752 16164
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 10744 16000 12434 16028
rect 13357 16031 13415 16037
rect 10744 15988 10750 16000
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13814 16028 13820 16040
rect 13403 16000 13820 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 15654 16028 15660 16040
rect 15615 16000 15660 16028
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 16390 16028 16396 16040
rect 16347 16000 16396 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 15013 15963 15071 15969
rect 15013 15929 15025 15963
rect 15059 15929 15071 15963
rect 15013 15923 15071 15929
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 15028 15892 15056 15923
rect 15102 15920 15108 15972
rect 15160 15960 15166 15972
rect 16500 15960 16528 16204
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 20070 16164 20076 16176
rect 19484 16136 20076 16164
rect 19484 16124 19490 16136
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 22066 16164 22094 16204
rect 22557 16201 22569 16235
rect 22603 16232 22615 16235
rect 23290 16232 23296 16244
rect 22603 16204 23296 16232
rect 22603 16201 22615 16204
rect 22557 16195 22615 16201
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 24581 16235 24639 16241
rect 24581 16201 24593 16235
rect 24627 16232 24639 16235
rect 24762 16232 24768 16244
rect 24627 16204 24768 16232
rect 24627 16201 24639 16204
rect 24581 16195 24639 16201
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25225 16235 25283 16241
rect 25225 16232 25237 16235
rect 24912 16204 25237 16232
rect 24912 16192 24918 16204
rect 25225 16201 25237 16204
rect 25271 16201 25283 16235
rect 32950 16232 32956 16244
rect 32911 16204 32956 16232
rect 25225 16195 25283 16201
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 23845 16167 23903 16173
rect 23845 16164 23857 16167
rect 22066 16136 23857 16164
rect 23845 16133 23857 16136
rect 23891 16164 23903 16167
rect 25777 16167 25835 16173
rect 25777 16164 25789 16167
rect 23891 16136 25789 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 25777 16133 25789 16136
rect 25823 16133 25835 16167
rect 25777 16127 25835 16133
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16632 16068 17049 16096
rect 16632 16056 16638 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 18414 16096 18420 16108
rect 18375 16068 18420 16096
rect 17773 16059 17831 16065
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17788 16028 17816 16059
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 19978 16096 19984 16108
rect 18555 16068 19984 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20312 16068 20545 16096
rect 20312 16056 20318 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 22152 16068 22477 16096
rect 22152 16056 22158 16068
rect 22465 16065 22477 16068
rect 22511 16096 22523 16099
rect 23109 16099 23167 16105
rect 23109 16096 23121 16099
rect 22511 16068 23121 16096
rect 22511 16065 22523 16068
rect 22465 16059 22523 16065
rect 23109 16065 23121 16068
rect 23155 16065 23167 16099
rect 24486 16096 24492 16108
rect 24447 16068 24492 16096
rect 23109 16059 23167 16065
rect 24486 16056 24492 16068
rect 24544 16056 24550 16108
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24820 16068 25145 16096
rect 24820 16056 24826 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 33045 16099 33103 16105
rect 33045 16065 33057 16099
rect 33091 16096 33103 16099
rect 37826 16096 37832 16108
rect 33091 16068 37832 16096
rect 33091 16065 33103 16068
rect 33045 16059 33103 16065
rect 37826 16056 37832 16068
rect 37884 16096 37890 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 37884 16068 38025 16096
rect 37884 16056 37890 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 19426 16028 19432 16040
rect 16908 16000 17816 16028
rect 19387 16000 19432 16028
rect 16908 15988 16914 16000
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 19576 16000 19625 16028
rect 19576 15988 19582 16000
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 20714 16028 20720 16040
rect 20675 16000 20720 16028
rect 19613 15991 19671 15997
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 23198 16028 23204 16040
rect 23159 16000 23204 16028
rect 23198 15988 23204 16000
rect 23256 15988 23262 16040
rect 38286 16028 38292 16040
rect 38247 16000 38292 16028
rect 38286 15988 38292 16000
rect 38344 15988 38350 16040
rect 15160 15932 16528 15960
rect 17129 15963 17187 15969
rect 15160 15920 15166 15932
rect 17129 15929 17141 15963
rect 17175 15960 17187 15963
rect 17175 15932 19656 15960
rect 17175 15929 17187 15932
rect 17129 15923 17187 15929
rect 19628 15904 19656 15932
rect 16298 15892 16304 15904
rect 15028 15864 16304 15892
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18230 15892 18236 15904
rect 17911 15864 18236 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 19610 15852 19616 15904
rect 19668 15852 19674 15904
rect 20073 15895 20131 15901
rect 20073 15861 20085 15895
rect 20119 15892 20131 15895
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20119 15864 20913 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 20901 15861 20913 15864
rect 20947 15892 20959 15895
rect 22002 15892 22008 15904
rect 20947 15864 22008 15892
rect 20947 15861 20959 15864
rect 20901 15855 20959 15861
rect 22002 15852 22008 15864
rect 22060 15852 22066 15904
rect 23934 15892 23940 15904
rect 23895 15864 23940 15892
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 10686 15688 10692 15700
rect 10647 15660 10692 15688
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 13630 15688 13636 15700
rect 13591 15660 13636 15688
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 14642 15688 14648 15700
rect 14603 15660 14648 15688
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 16574 15688 16580 15700
rect 14792 15660 16580 15688
rect 14792 15648 14798 15660
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 17589 15691 17647 15697
rect 17589 15657 17601 15691
rect 17635 15688 17647 15691
rect 19518 15688 19524 15700
rect 17635 15660 19524 15688
rect 17635 15657 17647 15660
rect 17589 15651 17647 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 20806 15688 20812 15700
rect 20763 15660 20812 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 21453 15691 21511 15697
rect 21453 15657 21465 15691
rect 21499 15688 21511 15691
rect 21818 15688 21824 15700
rect 21499 15660 21824 15688
rect 21499 15657 21511 15660
rect 21453 15651 21511 15657
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 22002 15688 22008 15700
rect 21963 15660 22008 15688
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 23385 15691 23443 15697
rect 23385 15657 23397 15691
rect 23431 15688 23443 15691
rect 23842 15688 23848 15700
rect 23431 15660 23848 15688
rect 23431 15657 23443 15660
rect 23385 15651 23443 15657
rect 23842 15648 23848 15660
rect 23900 15688 23906 15700
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 23900 15660 24593 15688
rect 23900 15648 23906 15660
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 31205 15691 31263 15697
rect 31205 15657 31217 15691
rect 31251 15688 31263 15691
rect 38010 15688 38016 15700
rect 31251 15660 38016 15688
rect 31251 15657 31263 15660
rect 31205 15651 31263 15657
rect 38010 15648 38016 15660
rect 38068 15648 38074 15700
rect 38286 15688 38292 15700
rect 38247 15660 38292 15688
rect 38286 15648 38292 15660
rect 38344 15648 38350 15700
rect 15010 15580 15016 15632
rect 15068 15620 15074 15632
rect 15068 15592 16252 15620
rect 15068 15580 15074 15592
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 15102 15552 15108 15564
rect 13964 15524 15108 15552
rect 13964 15512 13970 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15160 15524 15240 15552
rect 15160 15512 15166 15524
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 10594 15484 10600 15496
rect 2464 15456 10600 15484
rect 2464 15444 2470 15456
rect 10594 15444 10600 15456
rect 10652 15484 10658 15496
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 10652 15456 11253 15484
rect 10652 15444 10658 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 13814 15484 13820 15496
rect 13587 15456 13820 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 13814 15444 13820 15456
rect 13872 15484 13878 15496
rect 14642 15484 14648 15496
rect 13872 15456 14648 15484
rect 13872 15444 13878 15456
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15212 15493 15240 15524
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16224 15561 16252 15592
rect 16758 15580 16764 15632
rect 16816 15620 16822 15632
rect 17678 15620 17684 15632
rect 16816 15592 17684 15620
rect 16816 15580 16822 15592
rect 17678 15580 17684 15592
rect 17736 15620 17742 15632
rect 17736 15592 18552 15620
rect 17736 15580 17742 15592
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15712 15524 15945 15552
rect 15712 15512 15718 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 18322 15552 18328 15564
rect 18279 15524 18328 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18524 15561 18552 15592
rect 19426 15580 19432 15632
rect 19484 15580 19490 15632
rect 23474 15620 23480 15632
rect 20824 15592 23480 15620
rect 18509 15555 18567 15561
rect 18509 15521 18521 15555
rect 18555 15521 18567 15555
rect 19444 15552 19472 15580
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 19444 15524 19533 15552
rect 18509 15515 18567 15521
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 15197 15487 15255 15493
rect 14792 15456 14837 15484
rect 14792 15444 14798 15456
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 20824 15493 20852 15592
rect 23474 15580 23480 15592
rect 23532 15580 23538 15632
rect 23934 15580 23940 15632
rect 23992 15620 23998 15632
rect 35434 15620 35440 15632
rect 23992 15592 35440 15620
rect 23992 15580 23998 15592
rect 35434 15580 35440 15592
rect 35492 15580 35498 15632
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 22388 15524 22661 15552
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 17368 15456 17509 15484
rect 17368 15444 17374 15456
rect 17497 15453 17509 15456
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 16080 15388 16125 15416
rect 16080 15376 16086 15388
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 18380 15388 18425 15416
rect 18380 15376 18386 15388
rect 19610 15376 19616 15428
rect 19668 15416 19674 15428
rect 20165 15419 20223 15425
rect 19668 15388 19713 15416
rect 19668 15376 19674 15388
rect 20165 15385 20177 15419
rect 20211 15416 20223 15419
rect 21266 15416 21272 15428
rect 20211 15388 21272 15416
rect 20211 15385 20223 15388
rect 20165 15379 20223 15385
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 12158 15348 12164 15360
rect 12119 15320 12164 15348
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15348 13139 15351
rect 14550 15348 14556 15360
rect 13127 15320 14556 15348
rect 13127 15317 13139 15320
rect 13081 15311 13139 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15930 15348 15936 15360
rect 15335 15320 15936 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 21376 15348 21404 15447
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 22388 15484 22416 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 23753 15555 23811 15561
rect 23753 15521 23765 15555
rect 23799 15552 23811 15555
rect 25314 15552 25320 15564
rect 23799 15524 25320 15552
rect 23799 15521 23811 15524
rect 23753 15515 23811 15521
rect 25314 15512 25320 15524
rect 25372 15552 25378 15564
rect 25590 15552 25596 15564
rect 25372 15524 25596 15552
rect 25372 15512 25378 15524
rect 25590 15512 25596 15524
rect 25648 15512 25654 15564
rect 21508 15456 22416 15484
rect 22465 15487 22523 15493
rect 21508 15444 21514 15456
rect 22465 15453 22477 15487
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 22480 15416 22508 15447
rect 22738 15444 22744 15496
rect 22796 15484 22802 15496
rect 23569 15487 23627 15493
rect 23569 15484 23581 15487
rect 22796 15456 23581 15484
rect 22796 15444 22802 15456
rect 23569 15453 23581 15456
rect 23615 15453 23627 15487
rect 25038 15484 25044 15496
rect 24999 15456 25044 15484
rect 23569 15447 23627 15453
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25130 15444 25136 15496
rect 25188 15484 25194 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 25188 15456 25237 15484
rect 25188 15444 25194 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 31113 15487 31171 15493
rect 31113 15484 31125 15487
rect 29880 15456 31125 15484
rect 29880 15444 29886 15456
rect 31113 15453 31125 15456
rect 31159 15453 31171 15487
rect 31113 15447 31171 15453
rect 24670 15416 24676 15428
rect 22480 15388 24676 15416
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 16908 15320 21404 15348
rect 16908 15308 16914 15320
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 15470 15144 15476 15156
rect 10827 15116 15476 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 15565 15147 15623 15153
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 15746 15144 15752 15156
rect 15611 15116 15752 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 19334 15144 19340 15156
rect 16540 15116 18368 15144
rect 19295 15116 19340 15144
rect 16540 15104 16546 15116
rect 14366 15076 14372 15088
rect 13096 15048 14372 15076
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2130 15008 2136 15020
rect 1995 14980 2136 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2130 14968 2136 14980
rect 2188 15008 2194 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2188 14980 2421 15008
rect 2188 14968 2194 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4295 14980 4813 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4801 14977 4813 14980
rect 4847 15008 4859 15011
rect 7374 15008 7380 15020
rect 4847 14980 7380 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 7374 14968 7380 14980
rect 7432 15008 7438 15020
rect 10137 15011 10195 15017
rect 10137 15008 10149 15011
rect 7432 14980 10149 15008
rect 7432 14968 7438 14980
rect 10137 14977 10149 14980
rect 10183 15008 10195 15011
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10183 14980 10701 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 13096 15017 13124 15048
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 15378 15076 15384 15088
rect 15028 15048 15384 15076
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 11756 14980 12265 15008
rect 11756 14968 11762 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 13722 15008 13728 15020
rect 13587 14980 13728 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 15008 14243 15011
rect 14550 15008 14556 15020
rect 14231 14980 14556 15008
rect 14231 14977 14243 14980
rect 14185 14971 14243 14977
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 15028 15017 15056 15048
rect 15378 15036 15384 15048
rect 15436 15076 15442 15088
rect 16942 15076 16948 15088
rect 15436 15048 16948 15076
rect 15436 15036 15442 15048
rect 16942 15036 16948 15048
rect 17000 15036 17006 15088
rect 17037 15079 17095 15085
rect 17037 15045 17049 15079
rect 17083 15076 17095 15079
rect 17218 15076 17224 15088
rect 17083 15048 17224 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 18230 15076 18236 15088
rect 18191 15048 18236 15076
rect 18230 15036 18236 15048
rect 18288 15036 18294 15088
rect 18340 15076 18368 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20714 15144 20720 15156
rect 20027 15116 20720 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 21542 15144 21548 15156
rect 20824 15116 21548 15144
rect 20824 15088 20852 15116
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 22002 15104 22008 15156
rect 22060 15104 22066 15156
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 24762 15144 24768 15156
rect 23532 15116 24768 15144
rect 23532 15104 23538 15116
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 24857 15147 24915 15153
rect 24857 15113 24869 15147
rect 24903 15144 24915 15147
rect 25038 15144 25044 15156
rect 24903 15116 25044 15144
rect 24903 15113 24915 15116
rect 24857 15107 24915 15113
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 20806 15076 20812 15088
rect 18340 15048 20812 15076
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 22020 15076 22048 15104
rect 22097 15079 22155 15085
rect 22097 15076 22109 15079
rect 22020 15048 22109 15076
rect 22097 15045 22109 15048
rect 22143 15045 22155 15079
rect 22097 15039 22155 15045
rect 22189 15079 22247 15085
rect 22189 15045 22201 15079
rect 22235 15076 22247 15079
rect 22278 15076 22284 15088
rect 22235 15048 22284 15076
rect 22235 15045 22247 15048
rect 22189 15039 22247 15045
rect 22278 15036 22284 15048
rect 22336 15036 22342 15088
rect 24118 15076 24124 15088
rect 24079 15048 24124 15076
rect 24118 15036 24124 15048
rect 24176 15036 24182 15088
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 15028 14940 15056 14971
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15344 14980 15485 15008
rect 15344 14968 15350 14980
rect 15473 14977 15485 14980
rect 15519 15008 15531 15011
rect 16022 15008 16028 15020
rect 15519 14980 16028 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 16022 14968 16028 14980
rect 16080 15008 16086 15020
rect 16206 15008 16212 15020
rect 16080 14980 16212 15008
rect 16080 14968 16086 14980
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 19150 14968 19156 15020
rect 19208 15008 19214 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 19208 14980 19257 15008
rect 19208 14968 19214 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19886 15008 19892 15020
rect 19847 14980 19892 15008
rect 19245 14971 19303 14977
rect 10836 14912 15056 14940
rect 16301 14943 16359 14949
rect 10836 14900 10842 14912
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 16347 14912 16957 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 16945 14903 17003 14909
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 18141 14943 18199 14949
rect 17092 14912 17632 14940
rect 17092 14900 17098 14912
rect 1854 14832 1860 14884
rect 1912 14872 1918 14884
rect 14829 14875 14887 14881
rect 14829 14872 14841 14875
rect 1912 14844 14841 14872
rect 1912 14832 1918 14844
rect 14829 14841 14841 14844
rect 14875 14841 14887 14875
rect 14829 14835 14887 14841
rect 15194 14832 15200 14884
rect 15252 14872 15258 14884
rect 16390 14872 16396 14884
rect 15252 14844 16396 14872
rect 15252 14832 15258 14844
rect 16390 14832 16396 14844
rect 16448 14872 16454 14884
rect 17494 14872 17500 14884
rect 16448 14844 17500 14872
rect 16448 14832 16454 14844
rect 17494 14832 17500 14844
rect 17552 14832 17558 14884
rect 17604 14872 17632 14912
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18414 14940 18420 14952
rect 18187 14912 18420 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 19260 14940 19288 14971
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 24780 15017 24808 15104
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 24765 15011 24823 15017
rect 24765 14977 24777 15011
rect 24811 14977 24823 15011
rect 24765 14971 24823 14977
rect 21284 14940 21312 14971
rect 19260 14912 21312 14940
rect 21361 14943 21419 14949
rect 18506 14872 18512 14884
rect 17604 14844 18512 14872
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 18693 14875 18751 14881
rect 18693 14841 18705 14875
rect 18739 14841 18751 14875
rect 18693 14835 18751 14841
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 11296 14776 12173 14804
rect 11296 14764 11302 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13538 14804 13544 14816
rect 13035 14776 13544 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13633 14807 13691 14813
rect 13633 14773 13645 14807
rect 13679 14804 13691 14807
rect 13998 14804 14004 14816
rect 13679 14776 14004 14804
rect 13679 14773 13691 14776
rect 13633 14767 13691 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14277 14807 14335 14813
rect 14277 14773 14289 14807
rect 14323 14804 14335 14807
rect 15102 14804 15108 14816
rect 14323 14776 15108 14804
rect 14323 14773 14335 14776
rect 14277 14767 14335 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16298 14764 16304 14816
rect 16356 14804 16362 14816
rect 18708 14804 18736 14835
rect 19058 14804 19064 14816
rect 16356 14776 19064 14804
rect 16356 14764 16362 14776
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 21192 14804 21220 14912
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 22738 14940 22744 14952
rect 21407 14912 22744 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 22738 14900 22744 14912
rect 22796 14900 22802 14952
rect 23106 14940 23112 14952
rect 23067 14912 23112 14940
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 23569 14943 23627 14949
rect 23569 14940 23581 14943
rect 23256 14912 23581 14940
rect 23256 14900 23262 14912
rect 23569 14909 23581 14912
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 24213 14943 24271 14949
rect 24213 14909 24225 14943
rect 24259 14940 24271 14943
rect 25222 14940 25228 14952
rect 24259 14912 25228 14940
rect 24259 14909 24271 14912
rect 24213 14903 24271 14909
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 21542 14832 21548 14884
rect 21600 14872 21606 14884
rect 27154 14872 27160 14884
rect 21600 14844 27160 14872
rect 21600 14832 21606 14844
rect 27154 14832 27160 14844
rect 27212 14832 27218 14884
rect 24486 14804 24492 14816
rect 21192 14776 24492 14804
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 14182 14600 14188 14612
rect 12406 14572 14188 14600
rect 11698 14492 11704 14544
rect 11756 14492 11762 14544
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12406 14532 12434 14572
rect 14182 14560 14188 14572
rect 14240 14600 14246 14612
rect 14734 14600 14740 14612
rect 14240 14572 14740 14600
rect 14240 14560 14246 14572
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 17862 14600 17868 14612
rect 15712 14572 17868 14600
rect 15712 14560 15718 14572
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18380 14572 18429 14600
rect 18380 14560 18386 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 18417 14563 18475 14569
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18564 14572 24624 14600
rect 18564 14560 18570 14572
rect 12308 14504 12434 14532
rect 12308 14492 12314 14504
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 15746 14532 15752 14544
rect 14424 14504 15752 14532
rect 14424 14492 14430 14504
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 16482 14532 16488 14544
rect 15948 14504 16488 14532
rect 11716 14464 11744 14492
rect 15948 14476 15976 14504
rect 16482 14492 16488 14504
rect 16540 14532 16546 14544
rect 16540 14504 17264 14532
rect 16540 14492 16546 14504
rect 15010 14464 15016 14476
rect 11716 14436 12434 14464
rect 14971 14436 15016 14464
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12216 14368 12265 14396
rect 12216 14356 12222 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12406 14396 12434 14436
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15930 14464 15936 14476
rect 15891 14436 15936 14464
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 16206 14464 16212 14476
rect 16167 14436 16212 14464
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 17236 14473 17264 14504
rect 17494 14492 17500 14544
rect 17552 14532 17558 14544
rect 17552 14504 21404 14532
rect 17552 14492 17558 14504
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 17678 14464 17684 14476
rect 17639 14436 17684 14464
rect 17221 14427 17279 14433
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 19886 14464 19892 14476
rect 18524 14436 19892 14464
rect 18524 14405 18552 14436
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14464 20131 14467
rect 20254 14464 20260 14476
rect 20119 14436 20260 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 21376 14473 21404 14504
rect 21542 14492 21548 14544
rect 21600 14532 21606 14544
rect 24596 14532 24624 14572
rect 31294 14532 31300 14544
rect 21600 14504 23704 14532
rect 24596 14504 31300 14532
rect 21600 14492 21606 14504
rect 21361 14467 21419 14473
rect 21361 14433 21373 14467
rect 21407 14433 21419 14467
rect 22925 14467 22983 14473
rect 22925 14464 22937 14467
rect 21361 14427 21419 14433
rect 22204 14436 22937 14464
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 12406 14368 13553 14396
rect 12253 14359 12311 14365
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14365 18567 14399
rect 20806 14396 20812 14408
rect 20767 14368 20812 14396
rect 18509 14359 18567 14365
rect 10597 14331 10655 14337
rect 10597 14297 10609 14331
rect 10643 14328 10655 14331
rect 11149 14331 11207 14337
rect 11149 14328 11161 14331
rect 10643 14300 11161 14328
rect 10643 14297 10655 14300
rect 10597 14291 10655 14297
rect 11149 14297 11161 14300
rect 11195 14297 11207 14331
rect 11149 14291 11207 14297
rect 11238 14288 11244 14340
rect 11296 14328 11302 14340
rect 11793 14331 11851 14337
rect 11296 14300 11341 14328
rect 11296 14288 11302 14300
rect 11793 14297 11805 14331
rect 11839 14328 11851 14331
rect 12526 14328 12532 14340
rect 11839 14300 12532 14328
rect 11839 14297 11851 14300
rect 11793 14291 11851 14297
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 13081 14331 13139 14337
rect 13081 14297 13093 14331
rect 13127 14328 13139 14331
rect 14369 14331 14427 14337
rect 14369 14328 14381 14331
rect 13127 14300 14381 14328
rect 13127 14297 13139 14300
rect 13081 14291 13139 14297
rect 14369 14297 14381 14300
rect 14415 14297 14427 14331
rect 14369 14291 14427 14297
rect 14458 14288 14464 14340
rect 14516 14328 14522 14340
rect 16025 14331 16083 14337
rect 16025 14328 16037 14331
rect 14516 14300 14561 14328
rect 15856 14300 16037 14328
rect 14516 14288 14522 14300
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 12345 14263 12403 14269
rect 12345 14229 12357 14263
rect 12391 14260 12403 14263
rect 13354 14260 13360 14272
rect 12391 14232 13360 14260
rect 12391 14229 12403 14232
rect 12345 14223 12403 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15856 14260 15884 14300
rect 16025 14297 16037 14300
rect 16071 14297 16083 14331
rect 16025 14291 16083 14297
rect 16574 14288 16580 14340
rect 16632 14328 16638 14340
rect 17313 14331 17371 14337
rect 17313 14328 17325 14331
rect 16632 14300 17325 14328
rect 16632 14288 16638 14300
rect 17313 14297 17325 14300
rect 17359 14297 17371 14331
rect 17313 14291 17371 14297
rect 14976 14232 15884 14260
rect 14976 14220 14982 14232
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 18524 14260 18552 14359
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 19426 14328 19432 14340
rect 19387 14300 19432 14328
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19978 14328 19984 14340
rect 19939 14300 19984 14328
rect 19978 14288 19984 14300
rect 20036 14288 20042 14340
rect 21453 14331 21511 14337
rect 21453 14297 21465 14331
rect 21499 14297 21511 14331
rect 21453 14291 21511 14297
rect 15988 14232 18552 14260
rect 15988 14220 15994 14232
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 18840 14232 20729 14260
rect 18840 14220 18846 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 21468 14260 21496 14291
rect 21542 14288 21548 14340
rect 21600 14328 21606 14340
rect 22204 14328 22232 14436
rect 22925 14433 22937 14436
rect 22971 14433 22983 14467
rect 23198 14464 23204 14476
rect 23159 14436 23204 14464
rect 22925 14427 22983 14433
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 23676 14396 23704 14504
rect 31294 14492 31300 14504
rect 31352 14492 31358 14544
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 25222 14464 25228 14476
rect 24728 14436 24773 14464
rect 25183 14436 25228 14464
rect 24728 14424 24734 14436
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 23676 14368 24593 14396
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 26053 14399 26111 14405
rect 26053 14365 26065 14399
rect 26099 14396 26111 14399
rect 26326 14396 26332 14408
rect 26099 14368 26332 14396
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 26326 14356 26332 14368
rect 26384 14356 26390 14408
rect 26697 14399 26755 14405
rect 26697 14365 26709 14399
rect 26743 14396 26755 14399
rect 38010 14396 38016 14408
rect 26743 14368 27292 14396
rect 37971 14368 38016 14396
rect 26743 14365 26755 14368
rect 26697 14359 26755 14365
rect 22370 14328 22376 14340
rect 21600 14300 22232 14328
rect 22331 14300 22376 14328
rect 21600 14288 21606 14300
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 23014 14328 23020 14340
rect 22975 14300 23020 14328
rect 23014 14288 23020 14300
rect 23072 14288 23078 14340
rect 23382 14260 23388 14272
rect 21468 14232 23388 14260
rect 20717 14223 20775 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 25958 14260 25964 14272
rect 25919 14232 25964 14260
rect 25958 14220 25964 14232
rect 26016 14220 26022 14272
rect 26602 14260 26608 14272
rect 26563 14232 26608 14260
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 27264 14269 27292 14368
rect 38010 14356 38016 14368
rect 38068 14356 38074 14408
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 27249 14263 27307 14269
rect 27249 14229 27261 14263
rect 27295 14260 27307 14263
rect 34238 14260 34244 14272
rect 27295 14232 34244 14260
rect 27295 14229 27307 14232
rect 27249 14223 27307 14229
rect 34238 14220 34244 14232
rect 34296 14220 34302 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 10870 14056 10876 14068
rect 10643 14028 10876 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 14458 14056 14464 14068
rect 12207 14028 14464 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 18141 14059 18199 14065
rect 15620 14028 17080 14056
rect 15620 14016 15626 14028
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 13265 13991 13323 13997
rect 13265 13988 13277 13991
rect 11112 13960 13277 13988
rect 11112 13948 11118 13960
rect 13265 13957 13277 13960
rect 13311 13957 13323 13991
rect 13265 13951 13323 13957
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 13596 13960 14565 13988
rect 13596 13948 13602 13960
rect 14553 13957 14565 13960
rect 14599 13957 14611 13991
rect 14553 13951 14611 13957
rect 15105 13991 15163 13997
rect 15105 13957 15117 13991
rect 15151 13988 15163 13991
rect 15194 13988 15200 14000
rect 15151 13960 15200 13988
rect 15151 13957 15163 13960
rect 15105 13951 15163 13957
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15746 13988 15752 14000
rect 15707 13960 15752 13988
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 16482 13948 16488 14000
rect 16540 13988 16546 14000
rect 17052 13997 17080 14028
rect 18141 14025 18153 14059
rect 18187 14056 18199 14059
rect 18598 14056 18604 14068
rect 18187 14028 18604 14056
rect 18187 14025 18199 14028
rect 18141 14019 18199 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 37274 14056 37280 14068
rect 18708 14028 21588 14056
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 16540 13960 16957 13988
rect 16540 13948 16546 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 16945 13951 17003 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 18708 13988 18736 14028
rect 17736 13960 18736 13988
rect 17736 13948 17742 13960
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 19521 13991 19579 13997
rect 19521 13988 19533 13991
rect 19392 13960 19533 13988
rect 19392 13948 19398 13960
rect 19521 13957 19533 13960
rect 19567 13957 19579 13991
rect 19521 13951 19579 13957
rect 19613 13991 19671 13997
rect 19613 13957 19625 13991
rect 19659 13988 19671 13991
rect 21450 13988 21456 14000
rect 19659 13960 21456 13988
rect 19659 13957 19671 13960
rect 19613 13951 19671 13957
rect 21450 13948 21456 13960
rect 21508 13948 21514 14000
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 12158 13920 12164 13932
rect 1903 13892 12164 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 13906 13920 13912 13932
rect 12308 13892 12353 13920
rect 13556 13892 13912 13920
rect 12308 13880 12314 13892
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12584 13824 12725 13852
rect 12584 13812 12590 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 13354 13852 13360 13864
rect 13267 13824 13360 13852
rect 12713 13815 12771 13821
rect 13354 13812 13360 13824
rect 13412 13852 13418 13864
rect 13556 13852 13584 13892
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 18046 13920 18052 13932
rect 18007 13892 18052 13920
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 20312 13892 20453 13920
rect 20312 13880 20318 13892
rect 20441 13889 20453 13892
rect 20487 13889 20499 13923
rect 20441 13883 20499 13889
rect 13412 13824 13584 13852
rect 13412 13812 13418 13824
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 13688 13824 14473 13852
rect 13688 13812 13694 13824
rect 14461 13821 14473 13824
rect 14507 13821 14519 13855
rect 15654 13852 15660 13864
rect 14461 13815 14519 13821
rect 15028 13824 15660 13852
rect 7742 13744 7748 13796
rect 7800 13784 7806 13796
rect 15028 13784 15056 13824
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 7800 13756 15056 13784
rect 7800 13744 7806 13756
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 15948 13784 15976 13815
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16356 13824 16988 13852
rect 16356 13812 16362 13824
rect 15528 13756 15976 13784
rect 16960 13784 16988 13824
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 19337 13855 19395 13861
rect 19337 13852 19349 13855
rect 17092 13824 19349 13852
rect 17092 13812 17098 13824
rect 19337 13821 19349 13824
rect 19383 13852 19395 13855
rect 19426 13852 19432 13864
rect 19383 13824 19432 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20622 13852 20628 13864
rect 20583 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 21560 13852 21588 14028
rect 24412 14028 37280 14056
rect 22186 13988 22192 14000
rect 22147 13960 22192 13988
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 22370 13948 22376 14000
rect 22428 13988 22434 14000
rect 23106 13988 23112 14000
rect 22428 13960 23112 13988
rect 22428 13948 22434 13960
rect 23106 13948 23112 13960
rect 23164 13988 23170 14000
rect 24412 13988 24440 14028
rect 37274 14016 37280 14028
rect 37332 14016 37338 14068
rect 38286 14056 38292 14068
rect 38247 14028 38292 14056
rect 38286 14016 38292 14028
rect 38344 14016 38350 14068
rect 23164 13960 24440 13988
rect 24581 13991 24639 13997
rect 23164 13948 23170 13960
rect 24581 13957 24593 13991
rect 24627 13988 24639 13991
rect 25038 13988 25044 14000
rect 24627 13960 25044 13988
rect 24627 13957 24639 13960
rect 24581 13951 24639 13957
rect 25038 13948 25044 13960
rect 25096 13948 25102 14000
rect 26053 13991 26111 13997
rect 26053 13957 26065 13991
rect 26099 13988 26111 13991
rect 27522 13988 27528 14000
rect 26099 13960 27528 13988
rect 26099 13957 26111 13960
rect 26053 13951 26111 13957
rect 27522 13948 27528 13960
rect 27580 13948 27586 14000
rect 27154 13920 27160 13932
rect 27115 13892 27160 13920
rect 27154 13880 27160 13892
rect 27212 13880 27218 13932
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 21560 13824 22109 13852
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 24394 13852 24400 13864
rect 24355 13824 24400 13852
rect 22097 13815 22155 13821
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24670 13852 24676 13864
rect 24631 13824 24676 13852
rect 24670 13812 24676 13824
rect 24728 13812 24734 13864
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 28810 13852 28816 13864
rect 26191 13824 28816 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 28810 13812 28816 13824
rect 28868 13812 28874 13864
rect 34238 13812 34244 13864
rect 34296 13852 34302 13864
rect 35802 13852 35808 13864
rect 34296 13824 35808 13852
rect 34296 13812 34302 13824
rect 35802 13812 35808 13824
rect 35860 13812 35866 13864
rect 17497 13787 17555 13793
rect 17497 13784 17509 13787
rect 16960 13756 17509 13784
rect 15528 13744 15534 13756
rect 17497 13753 17509 13756
rect 17543 13753 17555 13787
rect 21542 13784 21548 13796
rect 17497 13747 17555 13753
rect 19306 13756 21548 13784
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 10560 13688 11161 13716
rect 10560 13676 10566 13688
rect 11149 13685 11161 13688
rect 11195 13716 11207 13719
rect 12894 13716 12900 13728
rect 11195 13688 12900 13716
rect 11195 13685 11207 13688
rect 11149 13679 11207 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 15194 13716 15200 13728
rect 13872 13688 15200 13716
rect 13872 13676 13878 13688
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 19306 13716 19334 13756
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 24302 13744 24308 13796
rect 24360 13784 24366 13796
rect 25593 13787 25651 13793
rect 25593 13784 25605 13787
rect 24360 13756 25605 13784
rect 24360 13744 24366 13756
rect 25593 13753 25605 13756
rect 25639 13753 25651 13787
rect 25593 13747 25651 13753
rect 15344 13688 19334 13716
rect 21085 13719 21143 13725
rect 15344 13676 15350 13688
rect 21085 13685 21097 13719
rect 21131 13716 21143 13719
rect 21174 13716 21180 13728
rect 21131 13688 21180 13716
rect 21131 13685 21143 13688
rect 21085 13679 21143 13685
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 24210 13716 24216 13728
rect 22244 13688 24216 13716
rect 22244 13676 22250 13688
rect 24210 13676 24216 13688
rect 24268 13676 24274 13728
rect 27801 13719 27859 13725
rect 27801 13685 27813 13719
rect 27847 13716 27859 13719
rect 27982 13716 27988 13728
rect 27847 13688 27988 13716
rect 27847 13685 27859 13688
rect 27801 13679 27859 13685
rect 27982 13676 27988 13688
rect 28040 13676 28046 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 11054 13512 11060 13524
rect 11015 13484 11060 13512
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 12989 13515 13047 13521
rect 12989 13481 13001 13515
rect 13035 13512 13047 13515
rect 14918 13512 14924 13524
rect 13035 13484 14924 13512
rect 13035 13481 13047 13484
rect 12989 13475 13047 13481
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 19889 13515 19947 13521
rect 15528 13484 18276 13512
rect 15528 13472 15534 13484
rect 1946 13404 1952 13456
rect 2004 13404 2010 13456
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 9953 13447 10011 13453
rect 9953 13444 9965 13447
rect 9916 13416 9965 13444
rect 9916 13404 9922 13416
rect 9953 13413 9965 13416
rect 9999 13444 10011 13447
rect 13538 13444 13544 13456
rect 9999 13416 13544 13444
rect 9999 13413 10011 13416
rect 9953 13407 10011 13413
rect 13538 13404 13544 13416
rect 13596 13404 13602 13456
rect 13633 13447 13691 13453
rect 13633 13413 13645 13447
rect 13679 13444 13691 13447
rect 13722 13444 13728 13456
rect 13679 13416 13728 13444
rect 13679 13413 13691 13416
rect 13633 13407 13691 13413
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 18248 13453 18276 13484
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20622 13512 20628 13524
rect 19935 13484 20628 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21821 13515 21879 13521
rect 21821 13481 21833 13515
rect 21867 13512 21879 13515
rect 23014 13512 23020 13524
rect 21867 13484 23020 13512
rect 21867 13481 21879 13484
rect 21821 13475 21879 13481
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 27985 13515 28043 13521
rect 27985 13512 27997 13515
rect 26476 13484 27997 13512
rect 26476 13472 26482 13484
rect 27985 13481 27997 13484
rect 28031 13481 28043 13515
rect 27985 13475 28043 13481
rect 18233 13447 18291 13453
rect 14752 13416 15148 13444
rect 1964 13376 1992 13404
rect 12345 13379 12403 13385
rect 1964 13348 11652 13376
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 1995 13280 2544 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2516 13184 2544 13280
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10962 13308 10968 13320
rect 10376 13280 10968 13308
rect 10376 13268 10382 13280
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11624 13317 11652 13348
rect 12345 13345 12357 13379
rect 12391 13376 12403 13379
rect 14752 13376 14780 13416
rect 15120 13388 15148 13416
rect 18233 13413 18245 13447
rect 18279 13413 18291 13447
rect 18233 13407 18291 13413
rect 21726 13404 21732 13456
rect 21784 13444 21790 13456
rect 22465 13447 22523 13453
rect 22465 13444 22477 13447
rect 21784 13416 22477 13444
rect 21784 13404 21790 13416
rect 22465 13413 22477 13416
rect 22511 13444 22523 13447
rect 23842 13444 23848 13456
rect 22511 13416 23848 13444
rect 22511 13413 22523 13416
rect 22465 13407 22523 13413
rect 23842 13404 23848 13416
rect 23900 13444 23906 13456
rect 24394 13444 24400 13456
rect 23900 13416 23980 13444
rect 23900 13404 23906 13416
rect 15028 13385 15148 13388
rect 12391 13348 14780 13376
rect 15013 13379 15148 13385
rect 12391 13345 12403 13348
rect 12345 13339 12403 13345
rect 15013 13345 15025 13379
rect 15059 13376 15148 13379
rect 15286 13376 15292 13388
rect 15059 13360 15292 13376
rect 15059 13345 15071 13360
rect 15120 13348 15292 13360
rect 15013 13339 15071 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 17034 13376 17040 13388
rect 16724 13348 17040 13376
rect 16724 13336 16730 13348
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 17313 13379 17371 13385
rect 17313 13345 17325 13379
rect 17359 13376 17371 13379
rect 19242 13376 19248 13388
rect 17359 13348 19248 13376
rect 17359 13345 17371 13348
rect 17313 13339 17371 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 20162 13336 20168 13388
rect 20220 13376 20226 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20220 13348 20637 13376
rect 20220 13336 20226 13348
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 21269 13379 21327 13385
rect 21269 13345 21281 13379
rect 21315 13376 21327 13379
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 21315 13348 23029 13376
rect 21315 13345 21327 13348
rect 21269 13339 21327 13345
rect 23017 13345 23029 13348
rect 23063 13376 23075 13379
rect 23198 13376 23204 13388
rect 23063 13348 23204 13376
rect 23063 13345 23075 13348
rect 23017 13339 23075 13345
rect 23198 13336 23204 13348
rect 23256 13336 23262 13388
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13308 11667 13311
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 11655 13280 12265 13308
rect 11655 13277 11667 13280
rect 11609 13271 11667 13277
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12894 13308 12900 13320
rect 12855 13280 12900 13308
rect 12253 13271 12311 13277
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 13814 13308 13820 13320
rect 13771 13280 13820 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 14274 13308 14280 13320
rect 13924 13280 14280 13308
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9364 13212 9413 13240
rect 9364 13200 9370 13212
rect 9401 13209 9413 13212
rect 9447 13240 9459 13243
rect 10226 13240 10232 13252
rect 9447 13212 10232 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13240 10563 13243
rect 10686 13240 10692 13252
rect 10551 13212 10692 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 10686 13200 10692 13212
rect 10744 13240 10750 13252
rect 13924 13240 13952 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 16298 13308 16304 13320
rect 16080 13280 16304 13308
rect 16080 13268 16086 13280
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 19794 13308 19800 13320
rect 19755 13280 19800 13308
rect 19794 13268 19800 13280
rect 19852 13268 19858 13320
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 23952 13308 23980 13416
rect 24044 13416 24400 13444
rect 24044 13385 24072 13416
rect 24394 13404 24400 13416
rect 24452 13444 24458 13456
rect 31202 13444 31208 13456
rect 24452 13416 31208 13444
rect 24452 13404 24458 13416
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13345 24087 13379
rect 24029 13339 24087 13345
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25188 13348 25237 13376
rect 25188 13336 25194 13348
rect 25225 13345 25237 13348
rect 25271 13376 25283 13379
rect 26142 13376 26148 13388
rect 25271 13348 26148 13376
rect 25271 13345 25283 13348
rect 25225 13339 25283 13345
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 27356 13385 27384 13416
rect 31202 13404 31208 13416
rect 31260 13404 31266 13456
rect 27341 13379 27399 13385
rect 27341 13345 27353 13379
rect 27387 13345 27399 13379
rect 27341 13339 27399 13345
rect 24486 13308 24492 13320
rect 23952 13280 24492 13308
rect 24486 13268 24492 13280
rect 24544 13268 24550 13320
rect 28077 13311 28135 13317
rect 28077 13277 28089 13311
rect 28123 13308 28135 13311
rect 28537 13311 28595 13317
rect 28537 13308 28549 13311
rect 28123 13280 28549 13308
rect 28123 13277 28135 13280
rect 28077 13271 28135 13277
rect 28537 13277 28549 13280
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 10744 13212 13952 13240
rect 10744 13200 10750 13212
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 15654 13240 15660 13252
rect 15160 13212 15205 13240
rect 15615 13212 15660 13240
rect 15160 13200 15166 13212
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 17218 13200 17224 13252
rect 17276 13240 17282 13252
rect 18414 13240 18420 13252
rect 17276 13212 17321 13240
rect 17420 13212 18420 13240
rect 17276 13200 17282 13212
rect 1762 13172 1768 13184
rect 1723 13144 1768 13172
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2498 13172 2504 13184
rect 2459 13144 2504 13172
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 11790 13172 11796 13184
rect 11751 13144 11796 13172
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 14366 13172 14372 13184
rect 14327 13144 14372 13172
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 16209 13175 16267 13181
rect 16209 13172 16221 13175
rect 15252 13144 16221 13172
rect 15252 13132 15258 13144
rect 16209 13141 16221 13144
rect 16255 13172 16267 13175
rect 17420 13172 17448 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13209 18751 13243
rect 18693 13203 18751 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13209 18843 13243
rect 18785 13203 18843 13209
rect 16255 13144 17448 13172
rect 16255 13141 16267 13144
rect 16209 13135 16267 13141
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 18708 13172 18736 13203
rect 17828 13144 18736 13172
rect 18800 13172 18828 13203
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 20772 13212 20817 13240
rect 20772 13200 20778 13212
rect 21358 13200 21364 13252
rect 21416 13240 21422 13252
rect 22278 13240 22284 13252
rect 21416 13212 22284 13240
rect 21416 13200 21422 13212
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 23109 13243 23167 13249
rect 23109 13209 23121 13243
rect 23155 13209 23167 13243
rect 24578 13240 24584 13252
rect 24539 13212 24584 13240
rect 23109 13203 23167 13209
rect 21726 13172 21732 13184
rect 18800 13144 21732 13172
rect 17828 13132 17834 13144
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 23124 13172 23152 13203
rect 24578 13200 24584 13212
rect 24636 13200 24642 13252
rect 25130 13240 25136 13252
rect 25091 13212 25136 13240
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 26050 13200 26056 13252
rect 26108 13240 26114 13252
rect 26421 13243 26479 13249
rect 26421 13240 26433 13243
rect 26108 13212 26433 13240
rect 26108 13200 26114 13212
rect 26421 13209 26433 13212
rect 26467 13209 26479 13243
rect 26421 13203 26479 13209
rect 26513 13243 26571 13249
rect 26513 13209 26525 13243
rect 26559 13240 26571 13243
rect 27338 13240 27344 13252
rect 26559 13212 27344 13240
rect 26559 13209 26571 13212
rect 26513 13203 26571 13209
rect 27338 13200 27344 13212
rect 27396 13200 27402 13252
rect 24394 13172 24400 13184
rect 23124 13144 24400 13172
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 24544 13144 25881 13172
rect 24544 13132 24550 13144
rect 25869 13141 25881 13144
rect 25915 13172 25927 13175
rect 28092 13172 28120 13271
rect 25915 13144 28120 13172
rect 25915 13141 25927 13144
rect 25869 13135 25927 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 2188 12940 9229 12968
rect 2188 12928 2194 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9217 12931 9275 12937
rect 9861 12971 9919 12977
rect 9861 12937 9873 12971
rect 9907 12968 9919 12971
rect 9907 12940 14136 12968
rect 9907 12937 9919 12940
rect 9861 12931 9919 12937
rect 2498 12860 2504 12912
rect 2556 12900 2562 12912
rect 7742 12900 7748 12912
rect 2556 12872 6914 12900
rect 7703 12872 7748 12900
rect 2556 12860 2562 12872
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 5534 12832 5540 12844
rect 1903 12804 5540 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 6886 12832 6914 12872
rect 7742 12860 7748 12872
rect 7800 12860 7806 12912
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 6886 12804 7665 12832
rect 7653 12801 7665 12804
rect 7699 12832 7711 12835
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7699 12804 8309 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 9232 12832 9260 12931
rect 10410 12860 10416 12912
rect 10468 12900 10474 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 10468 12872 12081 12900
rect 10468 12860 10474 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 13998 12900 14004 12912
rect 13959 12872 14004 12900
rect 12069 12863 12127 12869
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 14108 12900 14136 12940
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 23017 12971 23075 12977
rect 14424 12940 22416 12968
rect 14424 12928 14430 12940
rect 14108 12872 14596 12900
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 9232 12804 10333 12832
rect 8297 12795 8355 12801
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13538 12832 13544 12844
rect 13219 12804 13544 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12250 12764 12256 12776
rect 12023 12736 12256 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 11164 12696 11192 12727
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 13906 12764 13912 12776
rect 12406 12736 12664 12764
rect 13867 12736 13912 12764
rect 12406 12696 12434 12736
rect 12526 12696 12532 12708
rect 11164 12668 12434 12696
rect 12487 12668 12532 12696
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12636 12696 12664 12736
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14182 12764 14188 12776
rect 14143 12736 14188 12764
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14568 12764 14596 12872
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 15436 12872 15669 12900
rect 15436 12860 15442 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 15657 12863 15715 12869
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 17512 12909 17540 12940
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 16080 12872 17417 12900
rect 16080 12860 16086 12872
rect 17405 12869 17417 12872
rect 17451 12869 17463 12903
rect 17405 12863 17463 12869
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 17678 12900 17684 12912
rect 17543 12872 17684 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 18233 12903 18291 12909
rect 18233 12869 18245 12903
rect 18279 12900 18291 12903
rect 18598 12900 18604 12912
rect 18279 12872 18604 12900
rect 18279 12869 18291 12872
rect 18233 12863 18291 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 18782 12900 18788 12912
rect 18743 12872 18788 12900
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 20070 12900 20076 12912
rect 20031 12872 20076 12900
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 22278 12900 22284 12912
rect 20220 12872 20265 12900
rect 20364 12872 22284 12900
rect 20220 12860 20226 12872
rect 15286 12764 15292 12776
rect 14332 12736 14596 12764
rect 15247 12736 15292 12764
rect 14332 12724 14338 12736
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15712 12736 15761 12764
rect 15712 12724 15718 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 15749 12727 15807 12733
rect 14090 12696 14096 12708
rect 12636 12668 14096 12696
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 15764 12696 15792 12727
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16816 12736 16865 12764
rect 16816 12724 16822 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 17092 12736 18889 12764
rect 17092 12724 17098 12736
rect 18877 12733 18889 12736
rect 18923 12764 18935 12767
rect 20162 12764 20168 12776
rect 18923 12736 20168 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 20162 12724 20168 12736
rect 20220 12764 20226 12776
rect 20364 12764 20392 12872
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21450 12832 21456 12844
rect 20855 12804 21456 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 22388 12841 22416 12940
rect 23017 12937 23029 12971
rect 23063 12968 23075 12971
rect 23477 12971 23535 12977
rect 23477 12968 23489 12971
rect 23063 12940 23489 12968
rect 23063 12937 23075 12940
rect 23017 12931 23075 12937
rect 23477 12937 23489 12940
rect 23523 12968 23535 12971
rect 24581 12971 24639 12977
rect 24581 12968 24593 12971
rect 23523 12940 24593 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 24581 12937 24593 12940
rect 24627 12968 24639 12971
rect 24670 12968 24676 12980
rect 24627 12940 24676 12968
rect 24627 12937 24639 12940
rect 24581 12931 24639 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 25130 12928 25136 12980
rect 25188 12968 25194 12980
rect 27249 12971 27307 12977
rect 27249 12968 27261 12971
rect 25188 12940 27261 12968
rect 25188 12928 25194 12940
rect 27249 12937 27261 12940
rect 27295 12937 27307 12971
rect 27249 12931 27307 12937
rect 27522 12928 27528 12980
rect 27580 12968 27586 12980
rect 27893 12971 27951 12977
rect 27893 12968 27905 12971
rect 27580 12940 27905 12968
rect 27580 12928 27586 12940
rect 27893 12937 27905 12940
rect 27939 12937 27951 12971
rect 27893 12931 27951 12937
rect 28442 12928 28448 12980
rect 28500 12968 28506 12980
rect 28810 12968 28816 12980
rect 28500 12940 28816 12968
rect 28500 12928 28506 12940
rect 28810 12928 28816 12940
rect 28868 12928 28874 12980
rect 26602 12900 26608 12912
rect 24136 12872 26608 12900
rect 24136 12841 24164 12872
rect 26602 12860 26608 12872
rect 26660 12860 26666 12912
rect 38010 12900 38016 12912
rect 35866 12872 38016 12900
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 24121 12835 24179 12841
rect 24121 12832 24133 12835
rect 22373 12795 22431 12801
rect 22480 12804 24133 12832
rect 20990 12764 20996 12776
rect 20220 12736 20392 12764
rect 20951 12736 20996 12764
rect 20220 12724 20226 12736
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 22480 12764 22508 12804
rect 24121 12801 24133 12804
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25958 12832 25964 12844
rect 25087 12804 25964 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25958 12792 25964 12804
rect 26016 12792 26022 12844
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26160 12804 26433 12832
rect 21876 12736 22508 12764
rect 22557 12767 22615 12773
rect 21876 12724 21882 12736
rect 22557 12733 22569 12767
rect 22603 12764 22615 12767
rect 23750 12764 23756 12776
rect 22603 12736 23756 12764
rect 22603 12733 22615 12736
rect 22557 12727 22615 12733
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 23934 12764 23940 12776
rect 23895 12736 23940 12764
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 24688 12736 25237 12764
rect 19613 12699 19671 12705
rect 19613 12696 19625 12699
rect 14792 12668 19625 12696
rect 14792 12656 14798 12668
rect 19613 12665 19625 12668
rect 19659 12665 19671 12699
rect 21174 12696 21180 12708
rect 21135 12668 21180 12696
rect 19613 12659 19671 12665
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 24688 12640 24716 12736
rect 25225 12733 25237 12736
rect 25271 12733 25283 12767
rect 25225 12727 25283 12733
rect 25682 12724 25688 12776
rect 25740 12764 25746 12776
rect 26160 12764 26188 12804
rect 26421 12801 26433 12804
rect 26467 12832 26479 12835
rect 26786 12832 26792 12844
rect 26467 12804 26792 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 26786 12792 26792 12804
rect 26844 12792 26850 12844
rect 27154 12832 27160 12844
rect 27115 12804 27160 12832
rect 27154 12792 27160 12804
rect 27212 12792 27218 12844
rect 27982 12832 27988 12844
rect 27943 12804 27988 12832
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 28905 12835 28963 12841
rect 28905 12801 28917 12835
rect 28951 12832 28963 12835
rect 35866 12832 35894 12872
rect 38010 12860 38016 12872
rect 38068 12860 38074 12912
rect 28951 12804 35894 12832
rect 28951 12801 28963 12804
rect 28905 12795 28963 12801
rect 25740 12736 26188 12764
rect 26237 12767 26295 12773
rect 25740 12724 25746 12736
rect 26237 12733 26249 12767
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 26050 12696 26056 12708
rect 26011 12668 26056 12696
rect 26050 12656 26056 12668
rect 26108 12656 26114 12708
rect 26252 12696 26280 12727
rect 27062 12724 27068 12776
rect 27120 12764 27126 12776
rect 29365 12767 29423 12773
rect 29365 12764 29377 12767
rect 27120 12736 29377 12764
rect 27120 12724 27126 12736
rect 29365 12733 29377 12736
rect 29411 12733 29423 12767
rect 29365 12727 29423 12733
rect 34146 12724 34152 12776
rect 34204 12764 34210 12776
rect 38013 12767 38071 12773
rect 38013 12764 38025 12767
rect 34204 12736 38025 12764
rect 34204 12724 34210 12736
rect 38013 12733 38025 12736
rect 38059 12733 38071 12767
rect 38286 12764 38292 12776
rect 38247 12736 38292 12764
rect 38013 12727 38071 12733
rect 38286 12724 38292 12736
rect 38344 12724 38350 12776
rect 27522 12696 27528 12708
rect 26252 12668 27528 12696
rect 27522 12656 27528 12668
rect 27580 12656 27586 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 13170 12628 13176 12640
rect 10459 12600 13176 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12628 13323 12631
rect 24670 12628 24676 12640
rect 13311 12600 24676 12628
rect 13311 12597 13323 12600
rect 13265 12591 13323 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 30098 12628 30104 12640
rect 30059 12600 30104 12628
rect 30098 12588 30104 12600
rect 30156 12588 30162 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 5592 12396 7481 12424
rect 5592 12384 5598 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 14829 12427 14887 12433
rect 14829 12393 14841 12427
rect 14875 12424 14887 12427
rect 15746 12424 15752 12436
rect 14875 12396 15752 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 15896 12396 17049 12424
rect 15896 12384 15902 12396
rect 17037 12393 17049 12396
rect 17083 12424 17095 12427
rect 18785 12427 18843 12433
rect 17083 12396 18368 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 9217 12359 9275 12365
rect 9217 12325 9229 12359
rect 9263 12356 9275 12359
rect 13446 12356 13452 12368
rect 9263 12328 13452 12356
rect 9263 12325 9275 12328
rect 9217 12319 9275 12325
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 18340 12356 18368 12396
rect 18785 12393 18797 12427
rect 18831 12424 18843 12427
rect 19334 12424 19340 12436
rect 18831 12396 19340 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 20441 12427 20499 12433
rect 20441 12393 20453 12427
rect 20487 12424 20499 12427
rect 20714 12424 20720 12436
rect 20487 12396 20720 12424
rect 20487 12393 20499 12396
rect 20441 12387 20499 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 23750 12424 23756 12436
rect 23711 12396 23756 12424
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 25682 12424 25688 12436
rect 24504 12396 25688 12424
rect 19797 12359 19855 12365
rect 18340 12328 19334 12356
rect 12618 12288 12624 12300
rect 10152 12260 12624 12288
rect 10152 12232 10180 12260
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 14182 12288 14188 12300
rect 12768 12260 14188 12288
rect 12768 12248 12774 12260
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17678 12288 17684 12300
rect 17635 12260 17684 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 19306 12288 19334 12328
rect 19797 12325 19809 12359
rect 19843 12356 19855 12359
rect 20990 12356 20996 12368
rect 19843 12328 20996 12356
rect 19843 12325 19855 12328
rect 19797 12319 19855 12325
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 24302 12356 24308 12368
rect 22480 12328 24308 12356
rect 20898 12288 20904 12300
rect 19306 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 10134 12220 10140 12232
rect 7607 12192 10140 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10284 12192 10329 12220
rect 10612 12192 10885 12220
rect 10284 12180 10290 12192
rect 9766 12152 9772 12164
rect 9727 12124 9772 12152
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 9916 12124 10333 12152
rect 9916 12112 9922 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 8570 12084 8576 12096
rect 8531 12056 8576 12084
rect 8570 12044 8576 12056
rect 8628 12084 8634 12096
rect 10612 12084 10640 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 10873 12183 10931 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13504 12192 13553 12220
rect 13504 12180 13510 12192
rect 13541 12189 13553 12192
rect 13587 12220 13599 12223
rect 13998 12220 14004 12232
rect 13587 12192 14004 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14550 12220 14556 12232
rect 14332 12192 14556 12220
rect 14332 12180 14338 12192
rect 14550 12180 14556 12192
rect 14608 12220 14614 12232
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14608 12192 14749 12220
rect 14608 12180 14614 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18472 12192 18705 12220
rect 18472 12180 18478 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 20346 12220 20352 12232
rect 19751 12192 20352 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20533 12223 20591 12229
rect 20533 12189 20545 12223
rect 20579 12220 20591 12223
rect 20806 12220 20812 12232
rect 20579 12192 20812 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 12066 12112 12072 12164
rect 12124 12152 12130 12164
rect 12388 12161 12394 12164
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 12124 12124 12265 12152
rect 12124 12112 12130 12124
rect 12253 12121 12265 12124
rect 12299 12121 12311 12155
rect 12253 12115 12311 12121
rect 12345 12155 12394 12161
rect 12345 12121 12357 12155
rect 12391 12121 12394 12155
rect 12345 12115 12394 12121
rect 12388 12112 12394 12115
rect 12446 12112 12452 12164
rect 13633 12155 13691 12161
rect 13633 12121 13645 12155
rect 13679 12152 13691 12155
rect 15565 12155 15623 12161
rect 13679 12124 15516 12152
rect 13679 12121 13691 12124
rect 13633 12115 13691 12121
rect 10962 12084 10968 12096
rect 8628 12056 10640 12084
rect 10923 12056 10968 12084
rect 8628 12044 8634 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11609 12087 11667 12093
rect 11609 12053 11621 12087
rect 11655 12084 11667 12087
rect 14642 12084 14648 12096
rect 11655 12056 14648 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15488 12084 15516 12124
rect 15565 12121 15577 12155
rect 15611 12152 15623 12155
rect 15654 12152 15660 12164
rect 15611 12124 15660 12152
rect 15611 12121 15623 12124
rect 15565 12115 15623 12121
rect 15654 12112 15660 12124
rect 15712 12112 15718 12164
rect 16482 12152 16488 12164
rect 16443 12124 16488 12152
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 17681 12155 17739 12161
rect 17681 12152 17693 12155
rect 16592 12124 17693 12152
rect 16592 12084 16620 12124
rect 17681 12121 17693 12124
rect 17727 12121 17739 12155
rect 18230 12152 18236 12164
rect 18143 12124 18236 12152
rect 17681 12115 17739 12121
rect 18230 12112 18236 12124
rect 18288 12152 18294 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 18288 12124 21005 12152
rect 18288 12112 18294 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 21542 12152 21548 12164
rect 21503 12124 21548 12152
rect 20993 12115 21051 12121
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 21634 12112 21640 12164
rect 21692 12152 21698 12164
rect 21818 12152 21824 12164
rect 21692 12124 21824 12152
rect 21692 12112 21698 12124
rect 21818 12112 21824 12124
rect 21876 12112 21882 12164
rect 15488 12056 16620 12084
rect 18598 12044 18604 12096
rect 18656 12084 18662 12096
rect 22480 12084 22508 12328
rect 24302 12316 24308 12328
rect 24360 12316 24366 12368
rect 22646 12288 22652 12300
rect 22607 12260 22652 12288
rect 22646 12248 22652 12260
rect 22704 12248 22710 12300
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12288 23167 12291
rect 24504 12288 24532 12396
rect 25682 12384 25688 12396
rect 25740 12384 25746 12436
rect 26050 12424 26056 12436
rect 26011 12396 26056 12424
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 27522 12384 27528 12436
rect 27580 12424 27586 12436
rect 27617 12427 27675 12433
rect 27617 12424 27629 12427
rect 27580 12396 27629 12424
rect 27580 12384 27586 12396
rect 27617 12393 27629 12396
rect 27663 12393 27675 12427
rect 27617 12387 27675 12393
rect 25314 12316 25320 12368
rect 25372 12316 25378 12368
rect 26418 12316 26424 12368
rect 26476 12316 26482 12368
rect 26786 12316 26792 12368
rect 26844 12356 26850 12368
rect 28166 12356 28172 12368
rect 26844 12328 28172 12356
rect 26844 12316 26850 12328
rect 28166 12316 28172 12328
rect 28224 12356 28230 12368
rect 29825 12359 29883 12365
rect 29825 12356 29837 12359
rect 28224 12328 29837 12356
rect 28224 12316 28230 12328
rect 29825 12325 29837 12328
rect 29871 12325 29883 12359
rect 29825 12319 29883 12325
rect 30098 12316 30104 12368
rect 30156 12356 30162 12368
rect 37458 12356 37464 12368
rect 30156 12328 37464 12356
rect 30156 12316 30162 12328
rect 37458 12316 37464 12328
rect 37516 12316 37522 12368
rect 38286 12356 38292 12368
rect 38247 12328 38292 12356
rect 38286 12316 38292 12328
rect 38344 12316 38350 12368
rect 23155 12260 24532 12288
rect 25225 12291 25283 12297
rect 23155 12257 23167 12260
rect 23109 12251 23167 12257
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25332 12288 25360 12316
rect 25271 12260 25360 12288
rect 26237 12291 26295 12297
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 26237 12257 26249 12291
rect 26283 12288 26295 12291
rect 26436 12288 26464 12316
rect 27430 12288 27436 12300
rect 26283 12260 26464 12288
rect 26712 12260 27436 12288
rect 26283 12257 26295 12260
rect 26237 12251 26295 12257
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 24026 12220 24032 12232
rect 23891 12192 24032 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 26421 12223 26479 12229
rect 26421 12189 26433 12223
rect 26467 12220 26479 12223
rect 26602 12220 26608 12232
rect 26467 12192 26608 12220
rect 26467 12189 26479 12192
rect 26421 12183 26479 12189
rect 26602 12180 26608 12192
rect 26660 12220 26666 12232
rect 26712 12220 26740 12260
rect 27430 12248 27436 12260
rect 27488 12248 27494 12300
rect 26660 12192 26740 12220
rect 26660 12180 26666 12192
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 27062 12220 27068 12232
rect 26936 12192 27068 12220
rect 26936 12180 26942 12192
rect 27062 12180 27068 12192
rect 27120 12180 27126 12232
rect 27522 12220 27528 12232
rect 27483 12192 27528 12220
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 28074 12180 28080 12232
rect 28132 12220 28138 12232
rect 28169 12223 28227 12229
rect 28169 12220 28181 12223
rect 28132 12192 28181 12220
rect 28132 12180 28138 12192
rect 28169 12189 28181 12192
rect 28215 12189 28227 12223
rect 28994 12220 29000 12232
rect 28955 12192 29000 12220
rect 28169 12183 28227 12189
rect 28994 12180 29000 12192
rect 29052 12180 29058 12232
rect 29917 12223 29975 12229
rect 29917 12189 29929 12223
rect 29963 12220 29975 12223
rect 30116 12220 30144 12316
rect 29963 12192 30144 12220
rect 29963 12189 29975 12192
rect 29917 12183 29975 12189
rect 23040 12155 23098 12161
rect 23040 12121 23052 12155
rect 23086 12152 23098 12155
rect 23086 12124 24256 12152
rect 23086 12121 23098 12124
rect 23040 12115 23098 12121
rect 18656 12056 22508 12084
rect 24228 12084 24256 12124
rect 24302 12112 24308 12164
rect 24360 12152 24366 12164
rect 24581 12155 24639 12161
rect 24581 12152 24593 12155
rect 24360 12124 24593 12152
rect 24360 12112 24366 12124
rect 24581 12121 24593 12124
rect 24627 12121 24639 12155
rect 24581 12115 24639 12121
rect 25133 12155 25191 12161
rect 25133 12121 25145 12155
rect 25179 12152 25191 12155
rect 26973 12155 27031 12161
rect 26973 12152 26985 12155
rect 25179 12124 26985 12152
rect 25179 12121 25191 12124
rect 25133 12115 25191 12121
rect 26973 12121 26985 12124
rect 27019 12121 27031 12155
rect 26973 12115 27031 12121
rect 25406 12084 25412 12096
rect 24228 12056 25412 12084
rect 18656 12044 18662 12056
rect 25406 12044 25412 12056
rect 25464 12044 25470 12096
rect 25498 12044 25504 12096
rect 25556 12084 25562 12096
rect 28261 12087 28319 12093
rect 28261 12084 28273 12087
rect 25556 12056 28273 12084
rect 25556 12044 25562 12056
rect 28261 12053 28273 12056
rect 28307 12053 28319 12087
rect 28261 12047 28319 12053
rect 28350 12044 28356 12096
rect 28408 12084 28414 12096
rect 28905 12087 28963 12093
rect 28905 12084 28917 12087
rect 28408 12056 28917 12084
rect 28408 12044 28414 12056
rect 28905 12053 28917 12056
rect 28951 12053 28963 12087
rect 28905 12047 28963 12053
rect 29270 12044 29276 12096
rect 29328 12084 29334 12096
rect 30377 12087 30435 12093
rect 30377 12084 30389 12087
rect 29328 12056 30389 12084
rect 29328 12044 29334 12056
rect 30377 12053 30389 12056
rect 30423 12053 30435 12087
rect 30377 12047 30435 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 10410 11880 10416 11892
rect 10371 11852 10416 11880
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 15562 11880 15568 11892
rect 11020 11852 14228 11880
rect 15523 11852 15568 11880
rect 11020 11840 11026 11852
rect 8297 11815 8355 11821
rect 8297 11781 8309 11815
rect 8343 11812 8355 11815
rect 8343 11784 9674 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9214 11744 9220 11756
rect 8444 11716 9220 11744
rect 8444 11704 8450 11716
rect 9214 11704 9220 11716
rect 9272 11744 9278 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9272 11716 9321 11744
rect 9272 11704 9278 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9646 11744 9674 11784
rect 9950 11772 9956 11824
rect 10008 11812 10014 11824
rect 13357 11815 13415 11821
rect 13357 11812 13369 11815
rect 10008 11784 13369 11812
rect 10008 11772 10014 11784
rect 13357 11781 13369 11784
rect 13403 11781 13415 11815
rect 14090 11812 14096 11824
rect 14051 11784 14096 11812
rect 13357 11775 13415 11781
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14200 11821 14228 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 17678 11880 17684 11892
rect 16255 11852 17684 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 19613 11883 19671 11889
rect 17788 11852 18644 11880
rect 14185 11815 14243 11821
rect 14185 11781 14197 11815
rect 14231 11781 14243 11815
rect 14734 11812 14740 11824
rect 14695 11784 14740 11812
rect 14185 11775 14243 11781
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 15838 11772 15844 11824
rect 15896 11812 15902 11824
rect 17034 11812 17040 11824
rect 15896 11784 16160 11812
rect 16995 11784 17040 11812
rect 15896 11772 15902 11784
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9646 11716 10333 11744
rect 9309 11707 9367 11713
rect 10321 11713 10333 11716
rect 10367 11744 10379 11747
rect 10502 11744 10508 11756
rect 10367 11716 10508 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 10778 11676 10784 11688
rect 8895 11648 10784 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 10778 11636 10784 11648
rect 10836 11676 10842 11688
rect 10980 11676 11008 11707
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11204 11716 12173 11744
rect 11204 11704 11210 11716
rect 12161 11713 12173 11716
rect 12207 11744 12219 11747
rect 12250 11744 12256 11756
rect 12207 11716 12256 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12676 11716 12817 11744
rect 12676 11704 12682 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 15470 11744 15476 11756
rect 15383 11716 15476 11744
rect 12805 11707 12863 11713
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 15930 11744 15936 11756
rect 15528 11716 15936 11744
rect 15528 11704 15534 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16132 11753 16160 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 17126 11772 17132 11824
rect 17184 11812 17190 11824
rect 17788 11812 17816 11852
rect 17184 11784 17816 11812
rect 17184 11772 17190 11784
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 18616 11821 18644 11852
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 21174 11880 21180 11892
rect 19659 11852 21180 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 21174 11840 21180 11852
rect 21232 11880 21238 11892
rect 23934 11880 23940 11892
rect 21232 11852 22094 11880
rect 23895 11852 23940 11880
rect 21232 11840 21238 11852
rect 18509 11815 18567 11821
rect 18509 11812 18521 11815
rect 17920 11784 18521 11812
rect 17920 11772 17926 11784
rect 18509 11781 18521 11784
rect 18555 11781 18567 11815
rect 18509 11775 18567 11781
rect 18601 11815 18659 11821
rect 18601 11781 18613 11815
rect 18647 11781 18659 11815
rect 18601 11775 18659 11781
rect 21082 11772 21088 11824
rect 21140 11812 21146 11824
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 21140 11784 21281 11812
rect 21140 11772 21146 11784
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 21269 11775 21327 11781
rect 21361 11815 21419 11821
rect 21361 11781 21373 11815
rect 21407 11812 21419 11815
rect 21726 11812 21732 11824
rect 21407 11784 21732 11812
rect 21407 11781 21419 11784
rect 21361 11775 21419 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 22066 11812 22094 11852
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 25961 11883 26019 11889
rect 25961 11849 25973 11883
rect 26007 11880 26019 11883
rect 26050 11880 26056 11892
rect 26007 11852 26056 11880
rect 26007 11849 26019 11852
rect 25961 11843 26019 11849
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 27246 11880 27252 11892
rect 27207 11852 27252 11880
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 27488 11852 28549 11880
rect 27488 11840 27494 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 28537 11843 28595 11849
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 33226 11880 33232 11892
rect 30432 11852 33232 11880
rect 30432 11840 30438 11852
rect 33226 11840 33232 11852
rect 33284 11880 33290 11892
rect 34146 11880 34152 11892
rect 33284 11852 34152 11880
rect 33284 11840 33290 11852
rect 34146 11840 34152 11852
rect 34204 11840 34210 11892
rect 22373 11815 22431 11821
rect 22373 11812 22385 11815
rect 22066 11784 22385 11812
rect 22373 11781 22385 11784
rect 22419 11781 22431 11815
rect 22373 11775 22431 11781
rect 22465 11815 22523 11821
rect 22465 11781 22477 11815
rect 22511 11812 22523 11815
rect 22554 11812 22560 11824
rect 22511 11784 22560 11812
rect 22511 11781 22523 11784
rect 22465 11775 22523 11781
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 24762 11812 24768 11824
rect 24723 11784 24768 11812
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 30926 11812 30932 11824
rect 25332 11784 28028 11812
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16390 11744 16396 11756
rect 16163 11716 16396 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11744 19211 11747
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 19199 11716 20729 11744
rect 19199 11713 19211 11716
rect 19153 11707 19211 11713
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 23842 11744 23848 11756
rect 23803 11716 23848 11744
rect 20717 11707 20775 11713
rect 10836 11648 11008 11676
rect 13449 11679 13507 11685
rect 10836 11636 10842 11648
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 16666 11676 16672 11688
rect 13495 11648 16672 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11645 17003 11679
rect 17862 11676 17868 11688
rect 17823 11648 17868 11676
rect 16945 11639 17003 11645
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 13722 11608 13728 11620
rect 11103 11580 13728 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 16960 11608 16988 11639
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 20070 11676 20076 11688
rect 20031 11648 20076 11676
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11645 20315 11679
rect 20257 11639 20315 11645
rect 14240 11580 16988 11608
rect 14240 11568 14246 11580
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 12158 11540 12164 11552
rect 9447 11512 12164 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 16022 11540 16028 11552
rect 12299 11512 16028 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 20272 11540 20300 11639
rect 20732 11608 20760 11707
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 25332 11744 25360 11784
rect 25498 11744 25504 11756
rect 24627 11716 25360 11744
rect 25459 11716 25504 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 26326 11704 26332 11756
rect 26384 11744 26390 11756
rect 28000 11753 28028 11784
rect 28644 11784 30932 11812
rect 28644 11756 28672 11784
rect 30926 11772 30932 11784
rect 30984 11772 30990 11824
rect 26421 11747 26479 11753
rect 26421 11744 26433 11747
rect 26384 11716 26433 11744
rect 26384 11704 26390 11716
rect 26421 11713 26433 11716
rect 26467 11713 26479 11747
rect 26421 11707 26479 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27985 11747 28043 11753
rect 27985 11713 27997 11747
rect 28031 11713 28043 11747
rect 28626 11744 28632 11756
rect 28587 11716 28632 11744
rect 27985 11707 28043 11713
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 22649 11679 22707 11685
rect 22649 11676 22661 11679
rect 22520 11648 22661 11676
rect 22520 11636 22526 11648
rect 22649 11645 22661 11648
rect 22695 11645 22707 11679
rect 22649 11639 22707 11645
rect 25314 11636 25320 11688
rect 25372 11676 25378 11688
rect 25372 11648 25417 11676
rect 25372 11636 25378 11648
rect 25866 11636 25872 11688
rect 25924 11676 25930 11688
rect 26513 11679 26571 11685
rect 26513 11676 26525 11679
rect 25924 11648 26525 11676
rect 25924 11636 25930 11648
rect 26513 11645 26525 11648
rect 26559 11645 26571 11679
rect 26513 11639 26571 11645
rect 22738 11608 22744 11620
rect 20732 11580 22744 11608
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 23842 11568 23848 11620
rect 23900 11608 23906 11620
rect 27172 11608 27200 11707
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27893 11679 27951 11685
rect 27893 11676 27905 11679
rect 27488 11648 27905 11676
rect 27488 11636 27494 11648
rect 27893 11645 27905 11648
rect 27939 11645 27951 11679
rect 28000 11676 28028 11707
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 29270 11744 29276 11756
rect 29231 11716 29276 11744
rect 29270 11704 29276 11716
rect 29328 11704 29334 11756
rect 35894 11676 35900 11688
rect 28000 11648 35900 11676
rect 27893 11639 27951 11645
rect 35894 11636 35900 11648
rect 35952 11636 35958 11688
rect 23900 11580 27200 11608
rect 23900 11568 23906 11580
rect 27246 11568 27252 11620
rect 27304 11608 27310 11620
rect 27304 11580 27568 11608
rect 27304 11568 27310 11580
rect 21634 11540 21640 11552
rect 20272 11512 21640 11540
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 26234 11500 26240 11552
rect 26292 11540 26298 11552
rect 27430 11540 27436 11552
rect 26292 11512 27436 11540
rect 26292 11500 26298 11512
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27540 11540 27568 11580
rect 27982 11568 27988 11620
rect 28040 11608 28046 11620
rect 30374 11608 30380 11620
rect 28040 11580 30380 11608
rect 28040 11568 28046 11580
rect 30374 11568 30380 11580
rect 30432 11568 30438 11620
rect 29181 11543 29239 11549
rect 29181 11540 29193 11543
rect 27540 11512 29193 11540
rect 29181 11509 29193 11512
rect 29227 11509 29239 11543
rect 29730 11540 29736 11552
rect 29691 11512 29736 11540
rect 29181 11503 29239 11509
rect 29730 11500 29736 11512
rect 29788 11500 29794 11552
rect 30926 11540 30932 11552
rect 30839 11512 30932 11540
rect 30926 11500 30932 11512
rect 30984 11540 30990 11552
rect 33502 11540 33508 11552
rect 30984 11512 33508 11540
rect 30984 11500 30990 11512
rect 33502 11500 33508 11512
rect 33560 11500 33566 11552
rect 38286 11540 38292 11552
rect 38247 11512 38292 11540
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 12342 11336 12348 11348
rect 10643 11308 12348 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 15378 11336 15384 11348
rect 13924 11308 15384 11336
rect 9401 11271 9459 11277
rect 9401 11237 9413 11271
rect 9447 11268 9459 11271
rect 11054 11268 11060 11280
rect 9447 11240 11060 11268
rect 9447 11237 9459 11240
rect 9401 11231 9459 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11241 11271 11299 11277
rect 11241 11237 11253 11271
rect 11287 11268 11299 11271
rect 13924 11268 13952 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 15746 11336 15752 11348
rect 15620 11308 15752 11336
rect 15620 11296 15626 11308
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 16206 11336 16212 11348
rect 16080 11308 16212 11336
rect 16080 11296 16086 11308
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16540 11308 18920 11336
rect 16540 11296 16546 11308
rect 11287 11240 13952 11268
rect 11287 11237 11299 11240
rect 11241 11231 11299 11237
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 14700 11240 17264 11268
rect 14700 11228 14706 11240
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 11885 11203 11943 11209
rect 11885 11200 11897 11203
rect 9916 11172 11897 11200
rect 9916 11160 9922 11172
rect 11885 11169 11897 11172
rect 11931 11200 11943 11203
rect 12158 11200 12164 11212
rect 11931 11172 12164 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 12860 11172 13369 11200
rect 12860 11160 12866 11172
rect 13357 11169 13369 11172
rect 13403 11200 13415 11203
rect 16390 11200 16396 11212
rect 13403 11172 14044 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 8444 11104 8493 11132
rect 8444 11092 8450 11104
rect 8481 11101 8493 11104
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 11146 11132 11152 11144
rect 10735 11104 11152 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 10060 11064 10088 11095
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11606 11132 11612 11144
rect 11379 11104 11612 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11132 12682 11144
rect 12986 11132 12992 11144
rect 12676 11104 12992 11132
rect 12676 11092 12682 11104
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 11514 11064 11520 11076
rect 8404 11036 8616 11064
rect 10060 11036 11520 11064
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 8404 10996 8432 11036
rect 1912 10968 8432 10996
rect 8588 10996 8616 11036
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11033 12035 11067
rect 13541 11067 13599 11073
rect 13541 11064 13553 11067
rect 11977 11027 12035 11033
rect 13096 11036 13553 11064
rect 9582 10996 9588 11008
rect 8588 10968 9588 10996
rect 1912 10956 1918 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11992 10996 12020 11027
rect 11204 10968 12020 10996
rect 11204 10956 11210 10968
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 13096 10996 13124 11036
rect 13541 11033 13553 11036
rect 13587 11033 13599 11067
rect 13541 11027 13599 11033
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13814 11064 13820 11076
rect 13679 11036 13820 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14016 11064 14044 11172
rect 14660 11172 16396 11200
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14660 11141 14688 11172
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 17037 11203 17095 11209
rect 17037 11200 17049 11203
rect 17000 11172 17049 11200
rect 17000 11160 17006 11172
rect 17037 11169 17049 11172
rect 17083 11169 17095 11203
rect 17037 11163 17095 11169
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 14332 11104 14565 11132
rect 14332 11092 14338 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 15194 11132 15200 11144
rect 15155 11104 15200 11132
rect 14645 11095 14703 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16080 11104 16436 11132
rect 16080 11092 16086 11104
rect 15212 11064 15240 11092
rect 15746 11064 15752 11076
rect 14016 11036 15240 11064
rect 15707 11036 15752 11064
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16408 11073 16436 11104
rect 16393 11067 16451 11073
rect 15896 11036 15941 11064
rect 15896 11024 15902 11036
rect 16393 11033 16405 11067
rect 16439 11033 16451 11067
rect 16393 11027 16451 11033
rect 16945 11067 17003 11073
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 17236 11064 17264 11240
rect 18598 11228 18604 11280
rect 18656 11228 18662 11280
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11200 17923 11203
rect 18616 11200 18644 11228
rect 18892 11209 18920 11308
rect 20070 11296 20076 11348
rect 20128 11336 20134 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20128 11308 21005 11336
rect 20128 11296 20134 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 23842 11336 23848 11348
rect 21232 11308 23848 11336
rect 21232 11296 21238 11308
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 23937 11339 23995 11345
rect 23937 11305 23949 11339
rect 23983 11336 23995 11339
rect 24118 11336 24124 11348
rect 23983 11308 24124 11336
rect 23983 11305 23995 11308
rect 23937 11299 23995 11305
rect 24118 11296 24124 11308
rect 24176 11296 24182 11348
rect 24486 11296 24492 11348
rect 24544 11336 24550 11348
rect 24670 11336 24676 11348
rect 24544 11308 24676 11336
rect 24544 11296 24550 11308
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 25406 11296 25412 11348
rect 25464 11336 25470 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 25464 11308 25789 11336
rect 25464 11296 25470 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 29730 11336 29736 11348
rect 25777 11299 25835 11305
rect 27172 11308 29736 11336
rect 22186 11268 22192 11280
rect 20088 11240 22192 11268
rect 20088 11212 20116 11240
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 27065 11271 27123 11277
rect 27065 11268 27077 11271
rect 22388 11240 27077 11268
rect 17911 11172 18644 11200
rect 18877 11203 18935 11209
rect 17911 11169 17923 11172
rect 17865 11163 17923 11169
rect 18877 11169 18889 11203
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 18892 11132 18920 11163
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19116 11172 19625 11200
rect 19116 11160 19122 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 20070 11200 20076 11212
rect 20031 11172 20076 11200
rect 19613 11163 19671 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 21637 11203 21695 11209
rect 21637 11200 21649 11203
rect 21324 11172 21649 11200
rect 21324 11160 21330 11172
rect 21637 11169 21649 11172
rect 21683 11169 21695 11203
rect 21637 11163 21695 11169
rect 21726 11160 21732 11212
rect 21784 11200 21790 11212
rect 22388 11200 22416 11240
rect 27065 11237 27077 11240
rect 27111 11237 27123 11271
rect 27065 11231 27123 11237
rect 21784 11172 22416 11200
rect 21784 11160 21790 11172
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 22741 11203 22799 11209
rect 22741 11200 22753 11203
rect 22520 11172 22753 11200
rect 22520 11160 22526 11172
rect 22741 11169 22753 11172
rect 22787 11169 22799 11203
rect 22741 11163 22799 11169
rect 23106 11160 23112 11212
rect 23164 11200 23170 11212
rect 23750 11200 23756 11212
rect 23164 11172 23756 11200
rect 23164 11160 23170 11172
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24486 11160 24492 11212
rect 24544 11200 24550 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24544 11172 24593 11200
rect 24544 11160 24550 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 27172 11200 27200 11308
rect 29730 11296 29736 11308
rect 29788 11296 29794 11348
rect 28074 11228 28080 11280
rect 28132 11268 28138 11280
rect 29638 11268 29644 11280
rect 28132 11240 29644 11268
rect 28132 11228 28138 11240
rect 29638 11228 29644 11240
rect 29696 11228 29702 11280
rect 29822 11228 29828 11280
rect 29880 11268 29886 11280
rect 30466 11268 30472 11280
rect 29880 11240 30472 11268
rect 29880 11228 29886 11240
rect 30466 11228 30472 11240
rect 30524 11228 30530 11280
rect 24581 11163 24639 11169
rect 25884 11172 27200 11200
rect 27709 11203 27767 11209
rect 19426 11132 19432 11144
rect 18892 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20898 11132 20904 11144
rect 20859 11104 20904 11132
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11132 23443 11135
rect 23566 11132 23572 11144
rect 23431 11104 23572 11132
rect 23431 11101 23443 11104
rect 23385 11095 23443 11101
rect 16991 11036 17264 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 17586 11024 17592 11076
rect 17644 11064 17650 11076
rect 17957 11067 18015 11073
rect 17957 11064 17969 11067
rect 17644 11036 17969 11064
rect 17644 11024 17650 11036
rect 17957 11033 17969 11036
rect 18003 11033 18015 11067
rect 17957 11027 18015 11033
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20622 11064 20628 11076
rect 19751 11036 20628 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 21729 11067 21787 11073
rect 21729 11033 21741 11067
rect 21775 11033 21787 11067
rect 21729 11027 21787 11033
rect 22281 11067 22339 11073
rect 22281 11033 22293 11067
rect 22327 11064 22339 11067
rect 22462 11064 22468 11076
rect 22327 11036 22468 11064
rect 22327 11033 22339 11036
rect 22281 11027 22339 11033
rect 12400 10968 13124 10996
rect 12400 10956 12406 10968
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 16022 10996 16028 11008
rect 13228 10968 16028 10996
rect 13228 10956 13234 10968
rect 16022 10956 16028 10968
rect 16080 10956 16086 11008
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 21744 10996 21772 11027
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 22940 11064 22968 11095
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23768 11132 23796 11160
rect 25884 11144 25912 11172
rect 27709 11169 27721 11203
rect 27755 11200 27767 11203
rect 31018 11200 31024 11212
rect 27755 11172 31024 11200
rect 27755 11169 27767 11172
rect 27709 11163 27767 11169
rect 31018 11160 31024 11172
rect 31076 11160 31082 11212
rect 23837 11135 23895 11141
rect 23837 11132 23849 11135
rect 23768 11104 23849 11132
rect 23837 11101 23849 11104
rect 23883 11101 23895 11135
rect 23837 11095 23895 11101
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11134 24823 11135
rect 24811 11132 24900 11134
rect 25774 11132 25780 11144
rect 24811 11106 25780 11132
rect 24811 11101 24823 11106
rect 24872 11104 25780 11106
rect 24765 11095 24823 11101
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 26510 11132 26516 11144
rect 25924 11104 26017 11132
rect 26471 11104 26516 11132
rect 25924 11092 25930 11104
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 27157 11135 27215 11141
rect 27157 11101 27169 11135
rect 27203 11132 27215 11135
rect 27982 11132 27988 11144
rect 27203 11104 27988 11132
rect 27203 11101 27215 11104
rect 27157 11095 27215 11101
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 28905 11135 28963 11141
rect 28905 11101 28917 11135
rect 28951 11132 28963 11135
rect 29822 11132 29828 11144
rect 28951 11104 29828 11132
rect 28951 11101 28963 11104
rect 28905 11095 28963 11101
rect 29822 11092 29828 11104
rect 29880 11092 29886 11144
rect 29917 11135 29975 11141
rect 29917 11101 29929 11135
rect 29963 11132 29975 11135
rect 30006 11132 30012 11144
rect 29963 11104 30012 11132
rect 29963 11101 29975 11104
rect 29917 11095 29975 11101
rect 30006 11092 30012 11104
rect 30064 11132 30070 11144
rect 30377 11135 30435 11141
rect 30377 11132 30389 11135
rect 30064 11104 30389 11132
rect 30064 11092 30070 11104
rect 30377 11101 30389 11104
rect 30423 11101 30435 11135
rect 30377 11095 30435 11101
rect 30650 11092 30656 11144
rect 30708 11132 30714 11144
rect 38013 11135 38071 11141
rect 38013 11132 38025 11135
rect 30708 11104 38025 11132
rect 30708 11092 30714 11104
rect 38013 11101 38025 11104
rect 38059 11101 38071 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 38013 11095 38071 11101
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 26421 11067 26479 11073
rect 26421 11064 26433 11067
rect 22940 11036 26433 11064
rect 26421 11033 26433 11036
rect 26467 11033 26479 11067
rect 26421 11027 26479 11033
rect 26970 11024 26976 11076
rect 27028 11064 27034 11076
rect 28258 11064 28264 11076
rect 27028 11036 28120 11064
rect 28219 11036 28264 11064
rect 27028 11024 27034 11036
rect 16724 10968 21772 10996
rect 16724 10956 16730 10968
rect 21818 10956 21824 11008
rect 21876 10996 21882 11008
rect 25130 10996 25136 11008
rect 21876 10968 25136 10996
rect 21876 10956 21882 10968
rect 25130 10956 25136 10968
rect 25188 10956 25194 11008
rect 25222 10956 25228 11008
rect 25280 10996 25286 11008
rect 25280 10968 25325 10996
rect 25280 10956 25286 10968
rect 25498 10956 25504 11008
rect 25556 10996 25562 11008
rect 27982 10996 27988 11008
rect 25556 10968 27988 10996
rect 25556 10956 25562 10968
rect 27982 10956 27988 10968
rect 28040 10956 28046 11008
rect 28092 10996 28120 11036
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 28353 11067 28411 11073
rect 28353 11033 28365 11067
rect 28399 11033 28411 11067
rect 30469 11067 30527 11073
rect 30469 11064 30481 11067
rect 28353 11027 28411 11033
rect 29012 11036 30481 11064
rect 28368 10996 28396 11027
rect 28092 10968 28396 10996
rect 28534 10956 28540 11008
rect 28592 10996 28598 11008
rect 29012 10996 29040 11036
rect 30469 11033 30481 11036
rect 30515 11033 30527 11067
rect 30469 11027 30527 11033
rect 31113 11067 31171 11073
rect 31113 11033 31125 11067
rect 31159 11064 31171 11067
rect 31386 11064 31392 11076
rect 31159 11036 31392 11064
rect 31159 11033 31171 11036
rect 31113 11027 31171 11033
rect 31386 11024 31392 11036
rect 31444 11024 31450 11076
rect 28592 10968 29040 10996
rect 28592 10956 28598 10968
rect 29638 10956 29644 11008
rect 29696 10996 29702 11008
rect 29825 10999 29883 11005
rect 29825 10996 29837 10999
rect 29696 10968 29837 10996
rect 29696 10956 29702 10968
rect 29825 10965 29837 10968
rect 29871 10965 29883 10999
rect 29825 10959 29883 10965
rect 31294 10956 31300 11008
rect 31352 10996 31358 11008
rect 37918 10996 37924 11008
rect 31352 10968 37924 10996
rect 31352 10956 31358 10968
rect 37918 10956 37924 10968
rect 37976 10956 37982 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 10870 10792 10876 10804
rect 9907 10764 10876 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 20070 10792 20076 10804
rect 11103 10764 15608 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 8665 10727 8723 10733
rect 8665 10693 8677 10727
rect 8711 10724 8723 10727
rect 10413 10727 10471 10733
rect 8711 10696 10364 10724
rect 8711 10693 8723 10696
rect 8665 10687 8723 10693
rect 10336 10668 10364 10696
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 11146 10724 11152 10736
rect 10459 10696 11152 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 11296 10696 12173 10724
rect 11296 10684 11302 10696
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12710 10724 12716 10736
rect 12671 10696 12716 10724
rect 12161 10687 12219 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 13357 10727 13415 10733
rect 13357 10724 13369 10727
rect 12952 10696 13369 10724
rect 12952 10684 12958 10696
rect 13357 10693 13369 10696
rect 13403 10693 13415 10727
rect 13357 10687 13415 10693
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 14553 10727 14611 10733
rect 14553 10724 14565 10727
rect 13504 10696 14565 10724
rect 13504 10684 13510 10696
rect 14553 10693 14565 10696
rect 14599 10693 14611 10727
rect 15580 10724 15608 10764
rect 18984 10764 20076 10792
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 15580 10696 15761 10724
rect 14553 10687 14611 10693
rect 15749 10693 15761 10696
rect 15795 10693 15807 10727
rect 15749 10687 15807 10693
rect 16574 10684 16580 10736
rect 16632 10724 16638 10736
rect 17221 10727 17279 10733
rect 17221 10724 17233 10727
rect 16632 10696 17233 10724
rect 16632 10684 16638 10696
rect 17221 10693 17233 10696
rect 17267 10693 17279 10727
rect 17221 10687 17279 10693
rect 17402 10684 17408 10736
rect 17460 10724 17466 10736
rect 18984 10733 19012 10764
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21542 10792 21548 10804
rect 21131 10764 21548 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 23566 10792 23572 10804
rect 23527 10764 23572 10792
rect 23566 10752 23572 10764
rect 23624 10792 23630 10804
rect 24762 10792 24768 10804
rect 23624 10764 24768 10792
rect 23624 10752 23630 10764
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25280 10764 25973 10792
rect 25280 10752 25286 10764
rect 25961 10761 25973 10764
rect 26007 10792 26019 10795
rect 27617 10795 27675 10801
rect 27617 10792 27629 10795
rect 26007 10764 27629 10792
rect 26007 10761 26019 10764
rect 25961 10755 26019 10761
rect 27617 10761 27629 10764
rect 27663 10792 27675 10795
rect 28258 10792 28264 10804
rect 27663 10764 28264 10792
rect 27663 10761 27675 10764
rect 27617 10755 27675 10761
rect 28258 10752 28264 10764
rect 28316 10752 28322 10804
rect 28626 10752 28632 10804
rect 28684 10792 28690 10804
rect 28684 10764 30052 10792
rect 28684 10752 28690 10764
rect 18417 10727 18475 10733
rect 18417 10724 18429 10727
rect 17460 10696 18429 10724
rect 17460 10684 17466 10696
rect 18417 10693 18429 10696
rect 18463 10693 18475 10727
rect 18417 10687 18475 10693
rect 18969 10727 19027 10733
rect 18969 10693 18981 10727
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 19613 10727 19671 10733
rect 19613 10724 19625 10727
rect 19116 10696 19625 10724
rect 19116 10684 19122 10696
rect 19613 10693 19625 10696
rect 19659 10693 19671 10727
rect 22646 10724 22652 10736
rect 19613 10687 19671 10693
rect 20364 10696 22652 10724
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 9398 10656 9404 10668
rect 1903 10628 9404 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 10318 10656 10324 10668
rect 10279 10628 10324 10656
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 10962 10656 10968 10668
rect 10923 10628 10968 10656
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 16301 10659 16359 10665
rect 13964 10628 14009 10656
rect 13964 10616 13970 10628
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16758 10656 16764 10668
rect 16347 10628 16764 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 10928 10560 12081 10588
rect 10928 10548 10934 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 12216 10560 13277 10588
rect 12216 10548 12222 10560
rect 13265 10557 13277 10560
rect 13311 10588 13323 10591
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 13311 10560 14473 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 14461 10557 14473 10560
rect 14507 10557 14519 10591
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 14461 10551 14519 10557
rect 14936 10560 15669 10588
rect 10962 10520 10968 10532
rect 9140 10492 10968 10520
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9140 10461 9168 10492
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 14936 10520 14964 10560
rect 15657 10557 15669 10560
rect 15703 10588 15715 10591
rect 16942 10588 16948 10600
rect 15703 10560 16948 10588
rect 15703 10557 15715 10560
rect 15657 10551 15715 10557
rect 16942 10548 16948 10560
rect 17000 10588 17006 10600
rect 17129 10591 17187 10597
rect 17129 10588 17141 10591
rect 17000 10560 17141 10588
rect 17000 10548 17006 10560
rect 17129 10557 17141 10560
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 17405 10591 17463 10597
rect 17405 10557 17417 10591
rect 17451 10588 17463 10591
rect 18322 10588 18328 10600
rect 17451 10560 18000 10588
rect 18283 10560 18328 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 13964 10492 14964 10520
rect 13964 10480 13970 10492
rect 15010 10480 15016 10532
rect 15068 10520 15074 10532
rect 15068 10492 15113 10520
rect 15068 10480 15074 10492
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 17420 10520 17448 10551
rect 15896 10492 17448 10520
rect 17972 10520 18000 10560
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20070 10588 20076 10600
rect 19567 10560 20076 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20364 10520 20392 10696
rect 22646 10684 22652 10696
rect 22704 10684 22710 10736
rect 22925 10727 22983 10733
rect 22925 10693 22937 10727
rect 22971 10724 22983 10727
rect 24854 10724 24860 10736
rect 22971 10696 24860 10724
rect 22971 10693 22983 10696
rect 22925 10687 22983 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 25130 10684 25136 10736
rect 25188 10724 25194 10736
rect 25188 10696 28764 10724
rect 25188 10684 25194 10696
rect 20990 10656 20996 10668
rect 20903 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10656 21054 10668
rect 21910 10656 21916 10668
rect 21048 10628 21916 10656
rect 21048 10616 21054 10628
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 23198 10616 23204 10668
rect 23256 10656 23262 10668
rect 24213 10659 24271 10665
rect 23256 10628 24164 10656
rect 23256 10616 23262 10628
rect 20530 10548 20536 10600
rect 20588 10588 20594 10600
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 20588 10560 22017 10588
rect 20588 10548 20594 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22738 10548 22744 10600
rect 22796 10588 22802 10600
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22796 10560 23029 10588
rect 22796 10548 22802 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 24026 10588 24032 10600
rect 23987 10560 24032 10588
rect 23017 10551 23075 10557
rect 24026 10548 24032 10560
rect 24084 10548 24090 10600
rect 24136 10588 24164 10628
rect 24213 10625 24225 10659
rect 24259 10656 24271 10659
rect 24486 10656 24492 10668
rect 24259 10628 24492 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 24486 10616 24492 10628
rect 24544 10616 24550 10668
rect 25498 10656 25504 10668
rect 24780 10628 25504 10656
rect 24780 10588 24808 10628
rect 25498 10616 25504 10628
rect 25556 10616 25562 10668
rect 25774 10616 25780 10668
rect 25832 10656 25838 10668
rect 28074 10656 28080 10668
rect 25832 10628 26924 10656
rect 28035 10628 28080 10656
rect 25832 10616 25838 10628
rect 24136 10560 24808 10588
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25314 10588 25320 10600
rect 25271 10560 25320 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25314 10548 25320 10560
rect 25372 10548 25378 10600
rect 25409 10591 25467 10597
rect 25409 10557 25421 10591
rect 25455 10557 25467 10591
rect 26418 10588 26424 10600
rect 26379 10560 26424 10588
rect 25409 10551 25467 10557
rect 17972 10492 20392 10520
rect 15896 10480 15902 10492
rect 20438 10480 20444 10532
rect 20496 10520 20502 10532
rect 21818 10520 21824 10532
rect 20496 10492 21824 10520
rect 20496 10480 20502 10492
rect 21818 10480 21824 10492
rect 21876 10480 21882 10532
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 23934 10520 23940 10532
rect 21968 10492 23940 10520
rect 21968 10480 21974 10492
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 25424 10520 25452 10551
rect 26418 10548 26424 10560
rect 26476 10548 26482 10600
rect 26602 10588 26608 10600
rect 26563 10560 26608 10588
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 26896 10588 26924 10628
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 28166 10616 28172 10668
rect 28224 10656 28230 10668
rect 28736 10665 28764 10696
rect 30024 10665 30052 10764
rect 28261 10659 28319 10665
rect 28261 10656 28273 10659
rect 28224 10628 28273 10656
rect 28224 10616 28230 10628
rect 28261 10625 28273 10628
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28721 10659 28779 10665
rect 28721 10625 28733 10659
rect 28767 10625 28779 10659
rect 28721 10619 28779 10625
rect 29549 10659 29607 10665
rect 29549 10625 29561 10659
rect 29595 10625 29607 10659
rect 29549 10619 29607 10625
rect 30009 10659 30067 10665
rect 30009 10625 30021 10659
rect 30055 10625 30067 10659
rect 30009 10619 30067 10625
rect 30837 10659 30895 10665
rect 30837 10625 30849 10659
rect 30883 10656 30895 10659
rect 31386 10656 31392 10668
rect 30883 10628 31392 10656
rect 30883 10625 30895 10628
rect 30837 10619 30895 10625
rect 29457 10591 29515 10597
rect 29457 10588 29469 10591
rect 26896 10560 29469 10588
rect 29457 10557 29469 10560
rect 29503 10557 29515 10591
rect 29564 10588 29592 10619
rect 30852 10588 30880 10619
rect 31386 10616 31392 10628
rect 31444 10616 31450 10668
rect 37829 10659 37887 10665
rect 37829 10625 37841 10659
rect 37875 10656 37887 10659
rect 38010 10656 38016 10668
rect 37875 10628 38016 10656
rect 37875 10625 37887 10628
rect 37829 10619 37887 10625
rect 38010 10616 38016 10628
rect 38068 10616 38074 10668
rect 29564 10560 30880 10588
rect 29457 10551 29515 10557
rect 26620 10520 26648 10548
rect 25424 10492 26648 10520
rect 27062 10480 27068 10532
rect 27120 10520 27126 10532
rect 30745 10523 30803 10529
rect 30745 10520 30757 10523
rect 27120 10492 30757 10520
rect 27120 10480 27126 10492
rect 30745 10489 30757 10492
rect 30791 10489 30803 10523
rect 30745 10483 30803 10489
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 8720 10424 9137 10452
rect 8720 10412 8726 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 17402 10452 17408 10464
rect 13044 10424 17408 10452
rect 13044 10412 13050 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 20254 10452 20260 10464
rect 18932 10424 20260 10452
rect 18932 10412 18938 10424
rect 20254 10412 20260 10424
rect 20312 10452 20318 10464
rect 26326 10452 26332 10464
rect 20312 10424 26332 10452
rect 20312 10412 20318 10424
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 26786 10412 26792 10464
rect 26844 10452 26850 10464
rect 27246 10452 27252 10464
rect 26844 10424 27252 10452
rect 26844 10412 26850 10424
rect 27246 10412 27252 10424
rect 27304 10412 27310 10464
rect 27338 10412 27344 10464
rect 27396 10452 27402 10464
rect 28813 10455 28871 10461
rect 28813 10452 28825 10455
rect 27396 10424 28825 10452
rect 27396 10412 27402 10424
rect 28813 10421 28825 10424
rect 28859 10421 28871 10455
rect 30098 10452 30104 10464
rect 30059 10424 30104 10452
rect 28813 10415 28871 10421
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 31386 10452 31392 10464
rect 31347 10424 31392 10452
rect 31386 10412 31392 10424
rect 31444 10412 31450 10464
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 12802 10248 12808 10260
rect 9508 10220 12808 10248
rect 9508 10053 9536 10220
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 12986 10248 12992 10260
rect 12947 10220 12992 10248
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 19426 10248 19432 10260
rect 13679 10220 19432 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 22094 10248 22100 10260
rect 19628 10220 22100 10248
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 16114 10180 16120 10192
rect 9640 10152 14780 10180
rect 9640 10140 9646 10152
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10413 10115 10471 10121
rect 10413 10112 10425 10115
rect 10192 10084 10425 10112
rect 10192 10072 10198 10084
rect 10413 10081 10425 10084
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 12526 10112 12532 10124
rect 11103 10084 12532 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 10428 9908 10456 10075
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10081 14335 10115
rect 14752 10112 14780 10152
rect 15948 10152 16120 10180
rect 15948 10112 15976 10152
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 16577 10183 16635 10189
rect 16577 10149 16589 10183
rect 16623 10180 16635 10183
rect 16666 10180 16672 10192
rect 16623 10152 16672 10180
rect 16623 10149 16635 10152
rect 16577 10143 16635 10149
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 18874 10180 18880 10192
rect 18835 10152 18880 10180
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 19628 10180 19656 10220
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 24578 10248 24584 10260
rect 22204 10220 24584 10248
rect 22204 10180 22232 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 29825 10251 29883 10257
rect 29825 10248 29837 10251
rect 26476 10220 29837 10248
rect 26476 10208 26482 10220
rect 29825 10217 29837 10220
rect 29871 10217 29883 10251
rect 29825 10211 29883 10217
rect 19444 10152 19656 10180
rect 22066 10152 22232 10180
rect 22557 10183 22615 10189
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 14752 10084 15976 10112
rect 16316 10084 17141 10112
rect 14277 10075 14335 10081
rect 13078 10044 13084 10056
rect 13039 10016 13084 10044
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13412 10016 13553 10044
rect 13412 10004 13418 10016
rect 13541 10013 13553 10016
rect 13587 10044 13599 10047
rect 14292 10044 14320 10075
rect 16316 10056 16344 10084
rect 17129 10081 17141 10084
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 19444 10112 19472 10152
rect 17451 10084 19472 10112
rect 21361 10115 21419 10121
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 22066 10112 22094 10152
rect 22557 10149 22569 10183
rect 22603 10180 22615 10183
rect 22738 10180 22744 10192
rect 22603 10152 22744 10180
rect 22603 10149 22615 10152
rect 22557 10143 22615 10149
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 23952 10152 24900 10180
rect 21407 10084 22094 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 22646 10072 22652 10124
rect 22704 10112 22710 10124
rect 23952 10121 23980 10152
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 22704 10084 23305 10112
rect 22704 10072 22710 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 24673 10115 24731 10121
rect 24673 10081 24685 10115
rect 24719 10112 24731 10115
rect 24762 10112 24768 10124
rect 24719 10084 24768 10112
rect 24719 10081 24731 10084
rect 24673 10075 24731 10081
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 24872 10112 24900 10152
rect 26234 10140 26240 10192
rect 26292 10180 26298 10192
rect 30098 10180 30104 10192
rect 26292 10152 30104 10180
rect 26292 10140 26298 10152
rect 30098 10140 30104 10152
rect 30156 10140 30162 10192
rect 26786 10112 26792 10124
rect 24872 10084 26792 10112
rect 26786 10072 26792 10084
rect 26844 10112 26850 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26844 10084 26985 10112
rect 26844 10072 26850 10084
rect 26973 10081 26985 10084
rect 27019 10081 27031 10115
rect 26973 10075 27031 10081
rect 27154 10072 27160 10124
rect 27212 10112 27218 10124
rect 27249 10115 27307 10121
rect 27249 10112 27261 10115
rect 27212 10084 27261 10112
rect 27212 10072 27218 10084
rect 27249 10081 27261 10084
rect 27295 10112 27307 10115
rect 28534 10112 28540 10124
rect 27295 10084 28396 10112
rect 28495 10084 28540 10112
rect 27295 10081 27307 10084
rect 27249 10075 27307 10081
rect 13587 10016 14320 10044
rect 16025 10047 16083 10053
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 16025 10013 16037 10047
rect 16071 10044 16083 10047
rect 16298 10044 16304 10056
rect 16071 10016 16304 10044
rect 16071 10013 16083 10016
rect 16025 10007 16083 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9976 11023 9979
rect 11054 9976 11060 9988
rect 11011 9948 11060 9976
rect 11011 9945 11023 9948
rect 10965 9939 11023 9945
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 11609 9979 11667 9985
rect 11609 9945 11621 9979
rect 11655 9945 11667 9979
rect 12158 9976 12164 9988
rect 12119 9948 12164 9976
rect 11609 9939 11667 9945
rect 11624 9908 11652 9939
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 12253 9979 12311 9985
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 12618 9976 12624 9988
rect 12299 9948 12624 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14366 9976 14372 9988
rect 13964 9948 14372 9976
rect 13964 9936 13970 9948
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 15102 9936 15108 9988
rect 15160 9936 15166 9988
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9976 15807 9979
rect 15838 9976 15844 9988
rect 15795 9948 15844 9976
rect 15795 9945 15807 9948
rect 15749 9939 15807 9945
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 10428 9880 11652 9908
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 16500 9908 16528 10007
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 19426 10054 19432 10056
rect 19352 10044 19432 10054
rect 19024 10026 19432 10044
rect 19024 10016 19380 10026
rect 19024 10004 19030 10016
rect 19426 10004 19432 10026
rect 19484 10044 19490 10056
rect 19484 10016 19529 10044
rect 19484 10004 19490 10016
rect 19978 10004 19984 10056
rect 20036 10044 20042 10056
rect 20438 10044 20444 10056
rect 20036 10016 20444 10044
rect 20036 10004 20042 10016
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 26234 10044 26240 10056
rect 25608 10016 26240 10044
rect 19242 9976 19248 9988
rect 18630 9948 19248 9976
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19521 9979 19579 9985
rect 19521 9976 19533 9979
rect 19392 9948 19533 9976
rect 19392 9936 19398 9948
rect 19521 9945 19533 9948
rect 19567 9945 19579 9979
rect 19521 9939 19579 9945
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 20349 9979 20407 9985
rect 20349 9976 20361 9979
rect 19944 9948 20361 9976
rect 19944 9936 19950 9948
rect 20349 9945 20361 9948
rect 20395 9945 20407 9979
rect 21266 9976 21272 9988
rect 21227 9948 21272 9976
rect 20349 9939 20407 9945
rect 21266 9936 21272 9948
rect 21324 9936 21330 9988
rect 21994 9979 22052 9985
rect 21994 9976 22006 9979
rect 21376 9948 22006 9976
rect 13872 9880 16528 9908
rect 13872 9868 13878 9880
rect 18874 9868 18880 9920
rect 18932 9908 18938 9920
rect 19426 9908 19432 9920
rect 18932 9880 19432 9908
rect 18932 9868 18938 9880
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 21376 9908 21404 9948
rect 21994 9945 22006 9948
rect 22040 9945 22052 9979
rect 21994 9939 22052 9945
rect 22097 9979 22155 9985
rect 22097 9945 22109 9979
rect 22143 9976 22155 9979
rect 22186 9976 22192 9988
rect 22143 9948 22192 9976
rect 22143 9945 22155 9948
rect 22097 9939 22155 9945
rect 22186 9936 22192 9948
rect 22244 9936 22250 9988
rect 23845 9979 23903 9985
rect 23845 9945 23857 9979
rect 23891 9945 23903 9979
rect 23845 9939 23903 9945
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9976 24823 9979
rect 25608 9976 25636 10016
rect 26234 10004 26240 10016
rect 26292 10004 26298 10056
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10013 26387 10047
rect 28368 10044 28396 10084
rect 28534 10072 28540 10084
rect 28592 10072 28598 10124
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10112 28779 10115
rect 30377 10115 30435 10121
rect 30377 10112 30389 10115
rect 28767 10084 30389 10112
rect 28767 10081 28779 10084
rect 28721 10075 28779 10081
rect 30377 10081 30389 10084
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 29822 10044 29828 10056
rect 28368 10016 29828 10044
rect 26329 10007 26387 10013
rect 24811 9948 25636 9976
rect 24811 9945 24823 9948
rect 24765 9939 24823 9945
rect 19760 9880 21404 9908
rect 23860 9908 23888 9939
rect 25682 9936 25688 9988
rect 25740 9976 25746 9988
rect 25740 9948 25785 9976
rect 25740 9936 25746 9948
rect 26142 9936 26148 9988
rect 26200 9976 26206 9988
rect 26344 9976 26372 10007
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10044 29975 10047
rect 30282 10044 30288 10056
rect 29963 10016 30288 10044
rect 29963 10013 29975 10016
rect 29917 10007 29975 10013
rect 30282 10004 30288 10016
rect 30340 10004 30346 10056
rect 26200 9948 26372 9976
rect 26200 9936 26206 9948
rect 26237 9911 26295 9917
rect 26237 9908 26249 9911
rect 23860 9880 26249 9908
rect 19760 9868 19766 9880
rect 26237 9877 26249 9880
rect 26283 9877 26295 9911
rect 26344 9908 26372 9948
rect 27062 9936 27068 9988
rect 27120 9976 27126 9988
rect 31021 9979 31079 9985
rect 31021 9976 31033 9979
rect 27120 9948 27165 9976
rect 27264 9948 31033 9976
rect 27120 9936 27126 9948
rect 27264 9908 27292 9948
rect 31021 9945 31033 9948
rect 31067 9945 31079 9979
rect 31021 9939 31079 9945
rect 26344 9880 27292 9908
rect 26237 9871 26295 9877
rect 27706 9868 27712 9920
rect 27764 9908 27770 9920
rect 28077 9911 28135 9917
rect 28077 9908 28089 9911
rect 27764 9880 28089 9908
rect 27764 9868 27770 9880
rect 28077 9877 28089 9880
rect 28123 9877 28135 9911
rect 28077 9871 28135 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 16850 9704 16856 9716
rect 13136 9676 16856 9704
rect 13136 9664 13142 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20128 9676 21220 9704
rect 20128 9664 20134 9676
rect 9858 9636 9864 9648
rect 9819 9608 9864 9636
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 10413 9639 10471 9645
rect 10413 9605 10425 9639
rect 10459 9636 10471 9639
rect 11238 9636 11244 9648
rect 10459 9608 11244 9636
rect 10459 9605 10471 9608
rect 10413 9599 10471 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 11388 9608 12909 9636
rect 11388 9596 11394 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 14182 9636 14188 9648
rect 13495 9608 14188 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 14734 9596 14740 9648
rect 14792 9596 14798 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 15252 9608 17049 9636
rect 15252 9596 15258 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 21192 9636 21220 9676
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 22186 9704 22192 9716
rect 21600 9676 22192 9704
rect 21600 9664 21606 9676
rect 22186 9664 22192 9676
rect 22244 9664 22250 9716
rect 23400 9676 23704 9704
rect 23400 9636 23428 9676
rect 19826 9608 21128 9636
rect 21192 9608 22324 9636
rect 23138 9608 23428 9636
rect 17037 9599 17095 9605
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 8720 9540 10333 9568
rect 8720 9528 8726 9540
rect 10321 9537 10333 9540
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11882 9568 11888 9580
rect 11195 9540 11888 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12066 9568 12072 9580
rect 12027 9540 12072 9568
rect 12066 9528 12072 9540
rect 12124 9568 12130 9580
rect 12124 9540 12664 9568
rect 12124 9528 12130 9540
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9500 11115 9503
rect 12342 9500 12348 9512
rect 11103 9472 12348 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 9306 9432 9312 9444
rect 9267 9404 9312 9432
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 12636 9432 12664 9540
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 16666 9568 16672 9580
rect 16264 9540 16672 9568
rect 16264 9528 16270 9540
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 20993 9571 21051 9577
rect 20993 9568 21005 9571
rect 20916 9540 21005 9568
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 13630 9500 13636 9512
rect 12860 9472 13636 9500
rect 12860 9460 12866 9472
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 15749 9503 15807 9509
rect 13780 9472 15700 9500
rect 13780 9460 13786 9472
rect 13078 9432 13084 9444
rect 12636 9404 13084 9432
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 15672 9432 15700 9472
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 16298 9500 16304 9512
rect 15795 9472 16304 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16816 9472 16957 9500
rect 16816 9460 16822 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 17862 9500 17868 9512
rect 17823 9472 17868 9500
rect 16945 9463 17003 9469
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 19610 9460 19616 9512
rect 19668 9500 19674 9512
rect 20162 9500 20168 9512
rect 19668 9472 20168 9500
rect 19668 9460 19674 9472
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 17126 9432 17132 9444
rect 13832 9404 14136 9432
rect 15672 9404 17132 9432
rect 8662 9364 8668 9376
rect 8623 9336 8668 9364
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 12161 9367 12219 9373
rect 12161 9333 12173 9367
rect 12207 9364 12219 9367
rect 13832 9364 13860 9404
rect 12207 9336 13860 9364
rect 12207 9333 12219 9336
rect 12161 9327 12219 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13964 9336 14013 9364
rect 13964 9324 13970 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14108 9364 14136 9404
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 20916 9432 20944 9540
rect 20993 9537 21005 9540
rect 21039 9537 21051 9571
rect 21100 9568 21128 9608
rect 22186 9568 22192 9580
rect 21100 9540 22192 9568
rect 20993 9531 21051 9537
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 21082 9500 21088 9512
rect 21043 9472 21088 9500
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22296 9500 22324 9608
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23569 9639 23627 9645
rect 23569 9636 23581 9639
rect 23532 9608 23581 9636
rect 23532 9596 23538 9608
rect 23569 9605 23581 9608
rect 23615 9605 23627 9639
rect 23676 9636 23704 9676
rect 24578 9664 24584 9716
rect 24636 9704 24642 9716
rect 27246 9704 27252 9716
rect 24636 9676 27252 9704
rect 24636 9664 24642 9676
rect 27246 9664 27252 9676
rect 27304 9664 27310 9716
rect 24670 9636 24676 9648
rect 23676 9608 24676 9636
rect 23569 9599 23627 9605
rect 24670 9596 24676 9608
rect 24728 9596 24734 9648
rect 24946 9636 24952 9648
rect 24907 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25041 9639 25099 9645
rect 25041 9605 25053 9639
rect 25087 9636 25099 9639
rect 27614 9636 27620 9648
rect 25087 9608 27620 9636
rect 25087 9605 25099 9608
rect 25041 9599 25099 9605
rect 27614 9596 27620 9608
rect 27672 9596 27678 9648
rect 27709 9639 27767 9645
rect 27709 9605 27721 9639
rect 27755 9636 27767 9639
rect 28350 9636 28356 9648
rect 27755 9608 28356 9636
rect 27755 9605 27767 9608
rect 27709 9599 27767 9605
rect 28350 9596 28356 9608
rect 28408 9596 28414 9648
rect 28721 9639 28779 9645
rect 28721 9636 28733 9639
rect 28460 9608 28733 9636
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26878 9568 26884 9580
rect 25924 9540 26884 9568
rect 25924 9528 25930 9540
rect 26878 9528 26884 9540
rect 26936 9528 26942 9580
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 28460 9568 28488 9608
rect 28721 9605 28733 9608
rect 28767 9605 28779 9639
rect 28721 9599 28779 9605
rect 29273 9639 29331 9645
rect 29273 9605 29285 9639
rect 29319 9636 29331 9639
rect 30466 9636 30472 9648
rect 29319 9608 30472 9636
rect 29319 9605 29331 9608
rect 29273 9599 29331 9605
rect 30466 9596 30472 9608
rect 30524 9596 30530 9648
rect 30374 9568 30380 9580
rect 28040 9540 28488 9568
rect 30335 9540 30380 9568
rect 28040 9528 28046 9540
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 22152 9472 22197 9500
rect 22296 9472 23796 9500
rect 22152 9460 22158 9472
rect 23768 9432 23796 9472
rect 23842 9460 23848 9512
rect 23900 9500 23906 9512
rect 23900 9472 23945 9500
rect 23900 9460 23906 9472
rect 24946 9460 24952 9512
rect 25004 9500 25010 9512
rect 26234 9500 26240 9512
rect 25004 9472 26240 9500
rect 25004 9460 25010 9472
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 26418 9500 26424 9512
rect 26379 9472 26424 9500
rect 26418 9460 26424 9472
rect 26476 9460 26482 9512
rect 26602 9500 26608 9512
rect 26563 9472 26608 9500
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9500 27583 9503
rect 27614 9500 27620 9512
rect 27571 9472 27620 9500
rect 27571 9469 27583 9472
rect 27525 9463 27583 9469
rect 27614 9460 27620 9472
rect 27672 9460 27678 9512
rect 27798 9460 27804 9512
rect 27856 9500 27862 9512
rect 28442 9500 28448 9512
rect 27856 9472 28448 9500
rect 27856 9460 27862 9472
rect 28442 9460 28448 9472
rect 28500 9460 28506 9512
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9469 28687 9503
rect 29730 9500 29736 9512
rect 29691 9472 29736 9500
rect 28629 9463 28687 9469
rect 24489 9435 24547 9441
rect 24489 9432 24501 9435
rect 20916 9404 21312 9432
rect 23768 9404 24501 9432
rect 15378 9364 15384 9376
rect 14108 9336 15384 9364
rect 14001 9327 14059 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15491 9367 15549 9373
rect 15491 9333 15503 9367
rect 15537 9364 15549 9367
rect 15930 9364 15936 9376
rect 15537 9336 15936 9364
rect 15537 9333 15549 9336
rect 15491 9327 15549 9333
rect 15930 9324 15936 9336
rect 15988 9364 15994 9376
rect 16942 9364 16948 9376
rect 15988 9336 16948 9364
rect 15988 9324 15994 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 18046 9324 18052 9376
rect 18104 9364 18110 9376
rect 18598 9364 18604 9376
rect 18104 9336 18604 9364
rect 18104 9324 18110 9336
rect 18598 9324 18604 9336
rect 18656 9364 18662 9376
rect 18785 9367 18843 9373
rect 18785 9364 18797 9367
rect 18656 9336 18797 9364
rect 18656 9324 18662 9336
rect 18785 9333 18797 9336
rect 18831 9333 18843 9367
rect 18785 9327 18843 9333
rect 20275 9367 20333 9373
rect 20275 9333 20287 9367
rect 20321 9364 20333 9367
rect 21174 9364 21180 9376
rect 20321 9336 21180 9364
rect 20321 9333 20333 9336
rect 20275 9327 20333 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21284 9364 21312 9404
rect 24489 9401 24501 9404
rect 24535 9432 24547 9435
rect 27338 9432 27344 9444
rect 24535 9404 27344 9432
rect 24535 9401 24547 9404
rect 24489 9395 24547 9401
rect 27338 9392 27344 9404
rect 27396 9392 27402 9444
rect 27706 9432 27712 9444
rect 27448 9404 27712 9432
rect 24578 9364 24584 9376
rect 21284 9336 24584 9364
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 26237 9367 26295 9373
rect 26237 9333 26249 9367
rect 26283 9364 26295 9367
rect 27448 9364 27476 9404
rect 27706 9392 27712 9404
rect 27764 9432 27770 9444
rect 28644 9432 28672 9463
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 27764 9404 28672 9432
rect 27764 9392 27770 9404
rect 26283 9336 27476 9364
rect 26283 9333 26295 9336
rect 26237 9327 26295 9333
rect 27522 9324 27528 9376
rect 27580 9364 27586 9376
rect 30469 9367 30527 9373
rect 30469 9364 30481 9367
rect 27580 9336 30481 9364
rect 27580 9324 27586 9336
rect 30469 9333 30481 9336
rect 30515 9333 30527 9367
rect 30469 9327 30527 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 11057 9163 11115 9169
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11330 9160 11336 9172
rect 11103 9132 11336 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 12894 9160 12900 9172
rect 11747 9132 12900 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 15194 9160 15200 9172
rect 13035 9132 15200 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15344 9132 15884 9160
rect 15344 9120 15350 9132
rect 1854 9092 1860 9104
rect 1815 9064 1860 9092
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 12345 9095 12403 9101
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 13446 9092 13452 9104
rect 12391 9064 13452 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13633 9095 13691 9101
rect 13633 9061 13645 9095
rect 13679 9092 13691 9095
rect 13722 9092 13728 9104
rect 13679 9064 13728 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 15856 9092 15884 9132
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 19702 9160 19708 9172
rect 16448 9132 19708 9160
rect 16448 9120 16454 9132
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 23382 9160 23388 9172
rect 19812 9132 23244 9160
rect 23343 9132 23388 9160
rect 15856 9064 16436 9092
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9024 9459 9027
rect 10410 9024 10416 9036
rect 9447 8996 10416 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 10410 8984 10416 8996
rect 10468 9024 10474 9036
rect 10468 8996 13584 9024
rect 10468 8984 10474 8996
rect 11146 8956 11152 8968
rect 11107 8928 11152 8956
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 12342 8956 12348 8968
rect 11655 8928 12348 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 8570 8888 8576 8900
rect 8483 8860 8576 8888
rect 8570 8848 8576 8860
rect 8628 8888 8634 8900
rect 11624 8888 11652 8919
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 13556 8965 13584 8996
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 14056 8996 14289 9024
rect 14056 8984 14062 8996
rect 14277 8993 14289 8996
rect 14323 9024 14335 9027
rect 16408 9024 16436 9064
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 19812 9092 19840 9132
rect 18196 9064 19840 9092
rect 18196 9052 18202 9064
rect 20070 9052 20076 9104
rect 20128 9092 20134 9104
rect 20165 9095 20223 9101
rect 20165 9092 20177 9095
rect 20128 9064 20177 9092
rect 20128 9052 20134 9064
rect 20165 9061 20177 9064
rect 20211 9061 20223 9095
rect 20165 9055 20223 9061
rect 22278 9052 22284 9104
rect 22336 9092 22342 9104
rect 22741 9095 22799 9101
rect 22741 9092 22753 9095
rect 22336 9064 22753 9092
rect 22336 9052 22342 9064
rect 22741 9061 22753 9064
rect 22787 9092 22799 9095
rect 23106 9092 23112 9104
rect 22787 9064 23112 9092
rect 22787 9061 22799 9064
rect 22741 9055 22799 9061
rect 23106 9052 23112 9064
rect 23164 9052 23170 9104
rect 23216 9092 23244 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 23934 9160 23940 9172
rect 23895 9132 23940 9160
rect 23934 9120 23940 9132
rect 23992 9120 23998 9172
rect 26142 9160 26148 9172
rect 24688 9132 26148 9160
rect 24688 9092 24716 9132
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 26234 9120 26240 9172
rect 26292 9160 26298 9172
rect 27430 9160 27436 9172
rect 26292 9132 27436 9160
rect 26292 9120 26298 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 27522 9120 27528 9172
rect 27580 9160 27586 9172
rect 27580 9132 27660 9160
rect 27580 9120 27586 9132
rect 23216 9064 24716 9092
rect 25792 9064 27476 9092
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 14323 8996 16344 9024
rect 16408 8996 18613 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 16316 8968 16344 8996
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 25792 9033 25820 9064
rect 27264 9033 27384 9036
rect 25777 9027 25835 9033
rect 19484 8996 25728 9024
rect 19484 8984 19490 8996
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8956 13139 8959
rect 13541 8959 13599 8965
rect 13127 8928 13492 8956
rect 13127 8925 13139 8928
rect 13081 8919 13139 8925
rect 8628 8860 11652 8888
rect 12452 8888 12480 8919
rect 13262 8888 13268 8900
rect 12452 8860 13268 8888
rect 8628 8848 8634 8860
rect 13262 8848 13268 8860
rect 13320 8848 13326 8900
rect 13464 8888 13492 8928
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16758 8956 16764 8968
rect 16356 8928 16764 8956
rect 16356 8916 16362 8928
rect 16758 8916 16764 8928
rect 16816 8956 16822 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16816 8928 16865 8956
rect 16816 8916 16822 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 20990 8956 20996 8968
rect 20588 8928 20996 8956
rect 20588 8916 20594 8928
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8956 23535 8959
rect 23658 8956 23664 8968
rect 23523 8928 23664 8956
rect 23523 8925 23535 8928
rect 23477 8919 23535 8925
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 25590 8956 25596 8968
rect 25551 8928 25596 8956
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 25700 8956 25728 8996
rect 25777 8993 25789 9027
rect 25823 8993 25835 9027
rect 27264 9027 27399 9033
rect 27264 9024 27353 9027
rect 25777 8987 25835 8993
rect 26896 9008 27353 9024
rect 26896 8996 27292 9008
rect 26896 8968 26924 8996
rect 27341 8993 27353 9008
rect 27387 8993 27399 9027
rect 27341 8987 27399 8993
rect 26142 8956 26148 8968
rect 25700 8928 26148 8956
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 26694 8956 26700 8968
rect 26655 8928 26700 8956
rect 26694 8916 26700 8928
rect 26752 8916 26758 8968
rect 26878 8956 26884 8968
rect 26839 8928 26884 8956
rect 26878 8916 26884 8928
rect 26936 8916 26942 8968
rect 27448 8956 27476 9064
rect 27526 9027 27584 9033
rect 27526 8993 27538 9027
rect 27572 9024 27584 9027
rect 27632 9024 27660 9132
rect 27890 9120 27896 9172
rect 27948 9160 27954 9172
rect 27948 9132 29868 9160
rect 27948 9120 27954 9132
rect 29730 9092 29736 9104
rect 28092 9064 29736 9092
rect 27572 8996 27660 9024
rect 27572 8993 27584 8996
rect 27526 8987 27584 8993
rect 27706 8984 27712 9036
rect 27764 9024 27770 9036
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 27764 8996 27997 9024
rect 27764 8984 27770 8996
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 27985 8987 28043 8993
rect 28092 8956 28120 9064
rect 29730 9052 29736 9064
rect 29788 9052 29794 9104
rect 29840 9092 29868 9132
rect 30926 9120 30932 9172
rect 30984 9160 30990 9172
rect 37366 9160 37372 9172
rect 30984 9132 37372 9160
rect 30984 9120 30990 9132
rect 37366 9120 37372 9132
rect 37424 9120 37430 9172
rect 31481 9095 31539 9101
rect 31481 9092 31493 9095
rect 29840 9064 31493 9092
rect 31481 9061 31493 9064
rect 31527 9061 31539 9095
rect 31481 9055 31539 9061
rect 28166 8984 28172 9036
rect 28224 9024 28230 9036
rect 29822 9024 29828 9036
rect 28224 8996 29132 9024
rect 29783 8996 29828 9024
rect 28224 8984 28230 8996
rect 28902 8956 28908 8968
rect 27448 8928 28120 8956
rect 28863 8928 28908 8956
rect 28902 8916 28908 8928
rect 28960 8916 28966 8968
rect 29104 8965 29132 8996
rect 29822 8984 29828 8996
rect 29880 8984 29886 9036
rect 30466 9024 30472 9036
rect 30427 8996 30472 9024
rect 30466 8984 30472 8996
rect 30524 8984 30530 9036
rect 29089 8959 29147 8965
rect 29089 8925 29101 8959
rect 29135 8956 29147 8959
rect 29270 8956 29276 8968
rect 29135 8928 29276 8956
rect 29135 8925 29147 8928
rect 29089 8919 29147 8925
rect 29270 8916 29276 8928
rect 29328 8916 29334 8968
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 13464 8860 14504 8888
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9732 8792 9873 8820
rect 9732 8780 9738 8792
rect 9861 8789 9873 8792
rect 9907 8820 9919 8823
rect 10413 8823 10471 8829
rect 10413 8820 10425 8823
rect 9907 8792 10425 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 10413 8789 10425 8792
rect 10459 8789 10471 8823
rect 10413 8783 10471 8789
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 12802 8820 12808 8832
rect 10560 8792 12808 8820
rect 10560 8780 10566 8792
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 14366 8820 14372 8832
rect 13044 8792 14372 8820
rect 13044 8780 13050 8792
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14476 8820 14504 8860
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 16482 8888 16488 8900
rect 14608 8860 14653 8888
rect 15778 8860 16488 8888
rect 14608 8848 14614 8860
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17129 8891 17187 8897
rect 17129 8888 17141 8891
rect 16724 8860 17141 8888
rect 16724 8848 16730 8860
rect 17129 8857 17141 8860
rect 17175 8888 17187 8891
rect 19610 8888 19616 8900
rect 17175 8860 17540 8888
rect 18354 8860 19472 8888
rect 19571 8860 19616 8888
rect 17175 8857 17187 8860
rect 17129 8851 17187 8857
rect 15930 8820 15936 8832
rect 14476 8792 15936 8820
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16025 8823 16083 8829
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 17310 8820 17316 8832
rect 16071 8792 17316 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 17512 8820 17540 8860
rect 17954 8820 17960 8832
rect 17512 8792 17960 8820
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 19444 8820 19472 8860
rect 19610 8848 19616 8860
rect 19668 8848 19674 8900
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 19760 8860 19805 8888
rect 19760 8848 19766 8860
rect 20806 8848 20812 8900
rect 20864 8888 20870 8900
rect 21269 8891 21327 8897
rect 21269 8888 21281 8891
rect 20864 8860 21281 8888
rect 20864 8848 20870 8860
rect 21269 8857 21281 8860
rect 21315 8857 21327 8891
rect 24486 8888 24492 8900
rect 22494 8860 24492 8888
rect 21269 8851 21327 8857
rect 24486 8848 24492 8860
rect 24544 8848 24550 8900
rect 24578 8848 24584 8900
rect 24636 8888 24642 8900
rect 25498 8888 25504 8900
rect 24636 8860 24681 8888
rect 25056 8860 25504 8888
rect 24636 8848 24642 8860
rect 20714 8820 20720 8832
rect 19444 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 25056 8820 25084 8860
rect 25498 8848 25504 8860
rect 25556 8848 25562 8900
rect 26418 8848 26424 8900
rect 26476 8888 26482 8900
rect 29638 8888 29644 8900
rect 26476 8860 29644 8888
rect 26476 8848 26482 8860
rect 29638 8848 29644 8860
rect 29696 8848 29702 8900
rect 29914 8848 29920 8900
rect 29972 8888 29978 8900
rect 29972 8860 30017 8888
rect 29972 8848 29978 8860
rect 22244 8792 25084 8820
rect 25133 8823 25191 8829
rect 22244 8780 22250 8792
rect 25133 8789 25145 8823
rect 25179 8820 25191 8823
rect 26237 8823 26295 8829
rect 26237 8820 26249 8823
rect 25179 8792 26249 8820
rect 25179 8789 25191 8792
rect 25133 8783 25191 8789
rect 26237 8789 26249 8792
rect 26283 8820 26295 8823
rect 27062 8820 27068 8832
rect 26283 8792 27068 8820
rect 26283 8789 26295 8792
rect 26237 8783 26295 8789
rect 27062 8780 27068 8792
rect 27120 8820 27126 8832
rect 28445 8823 28503 8829
rect 28445 8820 28457 8823
rect 27120 8792 28457 8820
rect 27120 8780 27126 8792
rect 28445 8789 28457 8792
rect 28491 8789 28503 8823
rect 30926 8820 30932 8832
rect 30887 8792 30932 8820
rect 28445 8783 28503 8789
rect 30926 8780 30932 8792
rect 30984 8780 30990 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 11204 8588 12265 8616
rect 11204 8576 11210 8588
rect 12253 8585 12265 8588
rect 12299 8616 12311 8619
rect 12986 8616 12992 8628
rect 12299 8588 12992 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 15654 8616 15660 8628
rect 13136 8588 15660 8616
rect 13136 8576 13142 8588
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 18598 8616 18604 8628
rect 16040 8588 18604 8616
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 8352 8520 12558 8548
rect 8352 8508 8358 8520
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 16040 8557 16068 8588
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19150 8616 19156 8628
rect 19107 8588 19156 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 25774 8616 25780 8628
rect 21048 8588 21496 8616
rect 21048 8576 21054 8588
rect 16025 8551 16083 8557
rect 13688 8520 14858 8548
rect 13688 8508 13694 8520
rect 16025 8517 16037 8551
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17862 8548 17868 8560
rect 16816 8520 17868 8548
rect 16816 8508 16822 8520
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 16298 8489 16304 8492
rect 14056 8452 14101 8480
rect 14056 8440 14062 8452
rect 16294 8443 16304 8489
rect 16356 8480 16362 8492
rect 17328 8489 17356 8520
rect 17862 8508 17868 8520
rect 17920 8508 17926 8560
rect 19426 8548 19432 8560
rect 18814 8520 19432 8548
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 20622 8508 20628 8560
rect 20680 8508 20686 8560
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8548 21235 8551
rect 21266 8548 21272 8560
rect 21223 8520 21272 8548
rect 21223 8517 21235 8520
rect 21177 8511 21235 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 21468 8492 21496 8588
rect 23584 8588 25780 8616
rect 23584 8548 23612 8588
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26292 8588 26337 8616
rect 26292 8576 26298 8588
rect 26418 8576 26424 8628
rect 26476 8616 26482 8628
rect 27249 8619 27307 8625
rect 27249 8616 27261 8619
rect 26476 8588 27261 8616
rect 26476 8576 26482 8588
rect 27249 8585 27261 8588
rect 27295 8585 27307 8619
rect 29454 8616 29460 8628
rect 27249 8579 27307 8585
rect 27448 8588 29460 8616
rect 23750 8548 23756 8560
rect 23322 8520 23612 8548
rect 23711 8520 23756 8548
rect 23750 8508 23756 8520
rect 23808 8508 23814 8560
rect 23842 8508 23848 8560
rect 23900 8548 23906 8560
rect 23900 8520 24072 8548
rect 23900 8508 23906 8520
rect 17313 8483 17371 8489
rect 16356 8452 16394 8480
rect 16298 8440 16304 8443
rect 16356 8440 16362 8452
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 24044 8489 24072 8520
rect 24118 8508 24124 8560
rect 24176 8548 24182 8560
rect 24762 8548 24768 8560
rect 24176 8520 24768 8548
rect 24176 8508 24182 8520
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 27448 8548 27476 8588
rect 29454 8576 29460 8588
rect 29512 8576 29518 8628
rect 30374 8616 30380 8628
rect 30335 8588 30380 8616
rect 30374 8576 30380 8588
rect 30432 8576 30438 8628
rect 28258 8548 28264 8560
rect 25990 8520 27476 8548
rect 28219 8520 28264 8548
rect 28258 8508 28264 8520
rect 28316 8508 28322 8560
rect 29178 8548 29184 8560
rect 29091 8520 29184 8548
rect 29178 8508 29184 8520
rect 29236 8548 29242 8560
rect 30834 8548 30840 8560
rect 29236 8520 30840 8548
rect 29236 8508 29242 8520
rect 30834 8508 30840 8520
rect 30892 8508 30898 8560
rect 24029 8483 24087 8489
rect 21508 8452 21553 8480
rect 21508 8440 21514 8452
rect 24029 8449 24041 8483
rect 24075 8480 24087 8483
rect 24489 8483 24547 8489
rect 24489 8480 24501 8483
rect 24075 8452 24501 8480
rect 24075 8449 24087 8452
rect 24029 8443 24087 8449
rect 24489 8449 24501 8452
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 26786 8480 26792 8492
rect 26292 8452 26792 8480
rect 26292 8440 26298 8452
rect 26786 8440 26792 8452
rect 26844 8440 26850 8492
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 27522 8480 27528 8492
rect 27387 8452 27528 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 29086 8440 29092 8492
rect 29144 8480 29150 8492
rect 29641 8483 29699 8489
rect 29641 8480 29653 8483
rect 29144 8452 29653 8480
rect 29144 8440 29150 8452
rect 29641 8449 29653 8452
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8480 30527 8483
rect 30742 8480 30748 8492
rect 30515 8452 30748 8480
rect 30515 8449 30527 8452
rect 30469 8443 30527 8449
rect 30742 8440 30748 8452
rect 30800 8440 30806 8492
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 14553 8415 14611 8421
rect 14553 8412 14565 8415
rect 13771 8384 14565 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 14553 8381 14565 8384
rect 14599 8412 14611 8415
rect 15470 8412 15476 8424
rect 14599 8384 15476 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15654 8372 15660 8424
rect 15712 8412 15718 8424
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 15712 8384 17601 8412
rect 15712 8372 15718 8384
rect 17589 8381 17601 8384
rect 17635 8381 17647 8415
rect 17589 8375 17647 8381
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 18012 8384 22017 8412
rect 18012 8372 18018 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 24504 8384 25820 8412
rect 24504 8356 24532 8384
rect 19705 8347 19763 8353
rect 19705 8313 19717 8347
rect 19751 8344 19763 8347
rect 20162 8344 20168 8356
rect 19751 8316 20168 8344
rect 19751 8313 19763 8316
rect 19705 8307 19763 8313
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 21968 8316 22416 8344
rect 21968 8304 21974 8316
rect 9493 8279 9551 8285
rect 9493 8245 9505 8279
rect 9539 8276 9551 8279
rect 9674 8276 9680 8288
rect 9539 8248 9680 8276
rect 9539 8245 9551 8248
rect 9493 8239 9551 8245
rect 9674 8236 9680 8248
rect 9732 8276 9738 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9732 8248 9965 8276
rect 9732 8236 9738 8248
rect 9953 8245 9965 8248
rect 9999 8276 10011 8279
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 9999 8248 10517 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10505 8245 10517 8248
rect 10551 8276 10563 8279
rect 11057 8279 11115 8285
rect 11057 8276 11069 8279
rect 10551 8248 11069 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 11057 8245 11069 8248
rect 11103 8245 11115 8279
rect 11057 8239 11115 8245
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 17586 8276 17592 8288
rect 14516 8248 17592 8276
rect 14516 8236 14522 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 18966 8276 18972 8288
rect 17736 8248 18972 8276
rect 17736 8236 17742 8248
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 22278 8276 22284 8288
rect 19208 8248 22284 8276
rect 19208 8236 19214 8248
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 22388 8276 22416 8316
rect 24486 8304 24492 8356
rect 24544 8304 24550 8356
rect 25792 8344 25820 8384
rect 26142 8372 26148 8424
rect 26200 8412 26206 8424
rect 27614 8412 27620 8424
rect 26200 8384 27620 8412
rect 26200 8372 26206 8384
rect 27614 8372 27620 8384
rect 27672 8412 27678 8424
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 27672 8384 28181 8412
rect 27672 8372 27678 8384
rect 28169 8381 28181 8384
rect 28215 8381 28227 8415
rect 28169 8375 28227 8381
rect 29362 8372 29368 8424
rect 29420 8412 29426 8424
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 29420 8384 32321 8412
rect 29420 8372 29426 8384
rect 32309 8381 32321 8384
rect 32355 8381 32367 8415
rect 32309 8375 32367 8381
rect 30282 8344 30288 8356
rect 25792 8316 30288 8344
rect 30282 8304 30288 8316
rect 30340 8304 30346 8356
rect 29546 8276 29552 8288
rect 22388 8248 29552 8276
rect 29546 8236 29552 8248
rect 29604 8236 29610 8288
rect 29730 8276 29736 8288
rect 29691 8248 29736 8276
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 31018 8276 31024 8288
rect 30931 8248 31024 8276
rect 31018 8236 31024 8248
rect 31076 8276 31082 8288
rect 31570 8276 31576 8288
rect 31076 8248 31576 8276
rect 31076 8236 31082 8248
rect 31570 8236 31576 8248
rect 31628 8236 31634 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 12158 8072 12164 8084
rect 11379 8044 12164 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13320 8044 13645 8072
rect 13320 8032 13326 8044
rect 13633 8041 13645 8044
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14458 8072 14464 8084
rect 14419 8044 14464 8072
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 17034 8072 17040 8084
rect 15151 8044 17040 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 20530 8072 20536 8084
rect 17368 8044 20536 8072
rect 17368 8032 17374 8044
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21195 8075 21253 8081
rect 21195 8041 21207 8075
rect 21241 8072 21253 8075
rect 23658 8072 23664 8084
rect 21241 8044 23664 8072
rect 21241 8041 21253 8044
rect 21195 8035 21253 8041
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 24026 8032 24032 8084
rect 24084 8072 24090 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24084 8044 24685 8072
rect 24084 8032 24090 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 25317 8075 25375 8081
rect 25317 8072 25329 8075
rect 24912 8044 25329 8072
rect 24912 8032 24918 8044
rect 25317 8041 25329 8044
rect 25363 8041 25375 8075
rect 25317 8035 25375 8041
rect 25590 8032 25596 8084
rect 25648 8072 25654 8084
rect 28905 8075 28963 8081
rect 28905 8072 28917 8075
rect 25648 8044 28917 8072
rect 25648 8032 25654 8044
rect 28905 8041 28917 8044
rect 28951 8041 28963 8075
rect 28905 8035 28963 8041
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 29825 8075 29883 8081
rect 29825 8072 29837 8075
rect 29696 8044 29837 8072
rect 29696 8032 29702 8044
rect 29825 8041 29837 8044
rect 29871 8041 29883 8075
rect 30466 8072 30472 8084
rect 30427 8044 30472 8072
rect 29825 8035 29883 8041
rect 30466 8032 30472 8044
rect 30524 8032 30530 8084
rect 31754 8032 31760 8084
rect 31812 8072 31818 8084
rect 37734 8072 37740 8084
rect 31812 8044 37740 8072
rect 31812 8032 31818 8044
rect 37734 8032 37740 8044
rect 37792 8032 37798 8084
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 15010 8004 15016 8016
rect 14148 7976 15016 8004
rect 14148 7964 14154 7976
rect 15010 7964 15016 7976
rect 15068 7964 15074 8016
rect 18966 8004 18972 8016
rect 17696 7976 18972 8004
rect 13170 7936 13176 7948
rect 11440 7908 13176 7936
rect 11440 7877 11468 7908
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 16298 7936 16304 7948
rect 15703 7908 16304 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 17696 7945 17724 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 31113 8007 31171 8013
rect 31113 8004 31125 8007
rect 23308 7976 31125 8004
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 16448 7908 17693 7936
rect 16448 7896 16454 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 18233 7939 18291 7945
rect 18233 7936 18245 7939
rect 17920 7908 18245 7936
rect 17920 7896 17926 7908
rect 18233 7905 18245 7908
rect 18279 7936 18291 7939
rect 19426 7936 19432 7948
rect 18279 7908 19432 7936
rect 18279 7905 18291 7908
rect 18233 7899 18291 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 20714 7936 20720 7948
rect 19852 7908 20720 7936
rect 19852 7896 19858 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 22830 7896 22836 7948
rect 22888 7936 22894 7948
rect 23308 7936 23336 7976
rect 31113 7973 31125 7976
rect 31159 7973 31171 8007
rect 31113 7967 31171 7973
rect 23934 7936 23940 7948
rect 22888 7908 23336 7936
rect 23400 7908 23940 7936
rect 22888 7896 22894 7908
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7837 11943 7871
rect 11885 7831 11943 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7837 14611 7871
rect 15194 7868 15200 7880
rect 15155 7840 15200 7868
rect 14553 7831 14611 7837
rect 11900 7800 11928 7831
rect 12158 7800 12164 7812
rect 11900 7772 12020 7800
rect 12119 7772 12164 7800
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 9732 7704 10241 7732
rect 9732 7692 9738 7704
rect 10229 7701 10241 7704
rect 10275 7732 10287 7735
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10275 7704 10793 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 10781 7701 10793 7704
rect 10827 7732 10839 7735
rect 11992 7732 12020 7772
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 13446 7800 13452 7812
rect 13359 7772 13452 7800
rect 13446 7760 13452 7772
rect 13504 7800 13510 7812
rect 14568 7800 14596 7831
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 18874 7868 18880 7880
rect 18835 7840 18880 7868
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 22002 7868 22008 7880
rect 21508 7840 22008 7868
rect 21508 7828 21514 7840
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 23400 7854 23428 7908
rect 23934 7896 23940 7908
rect 23992 7896 23998 7948
rect 24029 7939 24087 7945
rect 24029 7905 24041 7939
rect 24075 7936 24087 7939
rect 24075 7908 25452 7936
rect 24075 7905 24087 7908
rect 24029 7899 24087 7905
rect 25424 7880 25452 7908
rect 25682 7896 25688 7948
rect 25740 7936 25746 7948
rect 26786 7936 26792 7948
rect 25740 7908 26792 7936
rect 25740 7896 25746 7908
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 27062 7936 27068 7948
rect 27023 7908 27068 7936
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 27614 7936 27620 7948
rect 27575 7908 27620 7936
rect 27614 7896 27620 7908
rect 27672 7896 27678 7948
rect 28261 7939 28319 7945
rect 28261 7905 28273 7939
rect 28307 7936 28319 7939
rect 28994 7936 29000 7948
rect 28307 7908 29000 7936
rect 28307 7905 28319 7908
rect 28261 7899 28319 7905
rect 28994 7896 29000 7908
rect 29052 7896 29058 7948
rect 23584 7840 24716 7868
rect 15838 7800 15844 7812
rect 13504 7772 14504 7800
rect 14568 7772 15844 7800
rect 13504 7760 13510 7772
rect 12526 7732 12532 7744
rect 10827 7704 12532 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 14476 7732 14504 7772
rect 15838 7760 15844 7772
rect 15896 7760 15902 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 16022 7800 16028 7812
rect 15979 7772 16028 7800
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 16022 7760 16028 7772
rect 16080 7800 16086 7812
rect 16206 7800 16212 7812
rect 16080 7772 16212 7800
rect 16080 7760 16086 7772
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 17586 7800 17592 7812
rect 17158 7772 17592 7800
rect 17586 7760 17592 7772
rect 17644 7760 17650 7812
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 18656 7772 19441 7800
rect 18656 7760 18662 7772
rect 19429 7769 19441 7772
rect 19475 7800 19487 7803
rect 22281 7803 22339 7809
rect 19475 7772 19932 7800
rect 20746 7772 20852 7800
rect 19475 7769 19487 7772
rect 19429 7763 19487 7769
rect 19794 7732 19800 7744
rect 14476 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 19904 7732 19932 7772
rect 20346 7732 20352 7744
rect 19904 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 20824 7732 20852 7772
rect 22281 7769 22293 7803
rect 22327 7769 22339 7803
rect 22281 7763 22339 7769
rect 22186 7732 22192 7744
rect 20824 7704 22192 7732
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22296 7732 22324 7763
rect 23584 7732 23612 7840
rect 24688 7800 24716 7840
rect 24762 7828 24768 7880
rect 24820 7868 24826 7880
rect 25406 7868 25412 7880
rect 24820 7840 24865 7868
rect 25367 7840 25412 7868
rect 24820 7828 24826 7840
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 28718 7828 28724 7880
rect 28776 7868 28782 7880
rect 28813 7871 28871 7877
rect 28813 7868 28825 7871
rect 28776 7840 28825 7868
rect 28776 7828 28782 7840
rect 28813 7837 28825 7840
rect 28859 7837 28871 7871
rect 28813 7831 28871 7837
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 30561 7871 30619 7877
rect 30561 7837 30573 7871
rect 30607 7868 30619 7871
rect 30742 7868 30748 7880
rect 30607 7840 30748 7868
rect 30607 7837 30619 7840
rect 30561 7831 30619 7837
rect 25958 7800 25964 7812
rect 24688 7772 25964 7800
rect 25958 7760 25964 7772
rect 26016 7760 26022 7812
rect 26973 7803 27031 7809
rect 26973 7769 26985 7803
rect 27019 7800 27031 7803
rect 27062 7800 27068 7812
rect 27019 7772 27068 7800
rect 27019 7769 27031 7772
rect 26973 7763 27031 7769
rect 27062 7760 27068 7772
rect 27120 7760 27126 7812
rect 28169 7803 28227 7809
rect 28169 7769 28181 7803
rect 28215 7769 28227 7803
rect 28169 7763 28227 7769
rect 22296 7704 23612 7732
rect 23658 7692 23664 7744
rect 23716 7732 23722 7744
rect 26326 7732 26332 7744
rect 23716 7704 26332 7732
rect 23716 7692 23722 7704
rect 26326 7692 26332 7704
rect 26384 7692 26390 7744
rect 28191 7732 28219 7763
rect 28534 7760 28540 7812
rect 28592 7800 28598 7812
rect 29730 7800 29736 7812
rect 28592 7772 29736 7800
rect 28592 7760 28598 7772
rect 29730 7760 29736 7772
rect 29788 7760 29794 7812
rect 29932 7800 29960 7831
rect 30742 7828 30748 7840
rect 30800 7828 30806 7880
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7868 31263 7871
rect 31294 7868 31300 7880
rect 31251 7840 31300 7868
rect 31251 7837 31263 7840
rect 31205 7831 31263 7837
rect 31294 7828 31300 7840
rect 31352 7828 31358 7880
rect 31386 7800 31392 7812
rect 29932 7772 31392 7800
rect 28350 7732 28356 7744
rect 28191 7704 28356 7732
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 28442 7692 28448 7744
rect 28500 7732 28506 7744
rect 29932 7732 29960 7772
rect 31386 7760 31392 7772
rect 31444 7800 31450 7812
rect 32217 7803 32275 7809
rect 32217 7800 32229 7803
rect 31444 7772 32229 7800
rect 31444 7760 31450 7772
rect 32217 7769 32229 7772
rect 32263 7769 32275 7803
rect 32217 7763 32275 7769
rect 28500 7704 29960 7732
rect 28500 7692 28506 7704
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 13446 7528 13452 7540
rect 11164 7500 13452 7528
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2038 7460 2044 7472
rect 1903 7432 2044 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2038 7420 2044 7432
rect 2096 7420 2102 7472
rect 9953 7463 10011 7469
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 11164 7460 11192 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 18141 7531 18199 7537
rect 15252 7500 18092 7528
rect 15252 7488 15258 7500
rect 13354 7460 13360 7472
rect 9999 7432 11192 7460
rect 13315 7432 13360 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 14369 7463 14427 7469
rect 14369 7460 14381 7463
rect 13780 7432 14381 7460
rect 13780 7420 13786 7432
rect 14369 7429 14381 7432
rect 14415 7429 14427 7463
rect 16482 7460 16488 7472
rect 15594 7432 16488 7460
rect 14369 7423 14427 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 16945 7463 17003 7469
rect 16945 7429 16957 7463
rect 16991 7460 17003 7463
rect 17678 7460 17684 7472
rect 16991 7432 17684 7460
rect 16991 7429 17003 7432
rect 16945 7423 17003 7429
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11790 7392 11796 7404
rect 11195 7364 11796 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12250 7352 12256 7404
rect 12308 7352 12314 7404
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 16960 7392 16988 7423
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 18064 7460 18092 7500
rect 18141 7497 18153 7531
rect 18187 7528 18199 7531
rect 19058 7528 19064 7540
rect 18187 7500 19064 7528
rect 18187 7497 18199 7500
rect 18141 7491 18199 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 20898 7528 20904 7540
rect 19168 7500 20904 7528
rect 18874 7460 18880 7472
rect 18064 7432 18880 7460
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19168 7460 19196 7500
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 21358 7528 21364 7540
rect 21319 7500 21364 7528
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 22370 7488 22376 7540
rect 22428 7528 22434 7540
rect 22428 7500 23612 7528
rect 22428 7488 22434 7500
rect 21910 7460 21916 7472
rect 19024 7432 19196 7460
rect 20194 7432 21916 7460
rect 19024 7420 19030 7432
rect 21910 7420 21916 7432
rect 21968 7420 21974 7472
rect 22278 7460 22284 7472
rect 22239 7432 22284 7460
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 23584 7460 23612 7500
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 23753 7531 23811 7537
rect 23753 7528 23765 7531
rect 23716 7500 23765 7528
rect 23716 7488 23722 7500
rect 23753 7497 23765 7500
rect 23799 7497 23811 7531
rect 23753 7491 23811 7497
rect 24210 7488 24216 7540
rect 24268 7528 24274 7540
rect 24397 7531 24455 7537
rect 24397 7528 24409 7531
rect 24268 7500 24409 7528
rect 24268 7488 24274 7500
rect 24397 7497 24409 7500
rect 24443 7497 24455 7531
rect 25038 7528 25044 7540
rect 24999 7500 25044 7528
rect 24397 7491 24455 7497
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 26436 7500 27844 7528
rect 25406 7460 25412 7472
rect 23584 7432 25412 7460
rect 25406 7420 25412 7432
rect 25464 7460 25470 7472
rect 25866 7460 25872 7472
rect 25464 7432 25872 7460
rect 25464 7420 25470 7432
rect 25866 7420 25872 7432
rect 25924 7420 25930 7472
rect 26436 7469 26464 7500
rect 26421 7463 26479 7469
rect 26421 7429 26433 7463
rect 26467 7429 26479 7463
rect 27154 7460 27160 7472
rect 27115 7432 27160 7460
rect 26421 7423 26479 7429
rect 27154 7420 27160 7432
rect 27212 7420 27218 7472
rect 27706 7460 27712 7472
rect 27667 7432 27712 7460
rect 27706 7420 27712 7432
rect 27764 7420 27770 7472
rect 27816 7460 27844 7500
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 28445 7531 28503 7537
rect 28445 7528 28457 7531
rect 28408 7500 28457 7528
rect 28408 7488 28414 7500
rect 28445 7497 28457 7500
rect 28491 7497 28503 7531
rect 28445 7491 28503 7497
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 28960 7500 29101 7528
rect 28960 7488 28966 7500
rect 29089 7497 29101 7500
rect 29135 7497 29147 7531
rect 29089 7491 29147 7497
rect 30377 7531 30435 7537
rect 30377 7497 30389 7531
rect 30423 7528 30435 7531
rect 30558 7528 30564 7540
rect 30423 7500 30564 7528
rect 30423 7497 30435 7500
rect 30377 7491 30435 7497
rect 30558 7488 30564 7500
rect 30616 7488 30622 7540
rect 29733 7463 29791 7469
rect 29733 7460 29745 7463
rect 27816 7432 29745 7460
rect 29733 7429 29745 7432
rect 29779 7429 29791 7463
rect 29733 7423 29791 7429
rect 16356 7364 16988 7392
rect 17589 7395 17647 7401
rect 16356 7352 16362 7364
rect 17589 7361 17601 7395
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18506 7392 18512 7404
rect 18279 7364 18512 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7324 8907 7327
rect 12268 7324 12296 7352
rect 8895 7296 12296 7324
rect 13633 7327 13691 7333
rect 8895 7293 8907 7296
rect 8849 7287 8907 7293
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 14090 7324 14096 7336
rect 13679 7296 14096 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 14918 7284 14924 7336
rect 14976 7324 14982 7336
rect 17310 7324 17316 7336
rect 14976 7296 17316 7324
rect 14976 7284 14982 7296
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17604 7324 17632 7355
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 20530 7352 20536 7404
rect 20588 7392 20594 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20588 7364 20729 7392
rect 20588 7352 20594 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21358 7392 21364 7404
rect 21315 7364 21364 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 23382 7352 23388 7404
rect 23440 7352 23446 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24854 7392 24860 7404
rect 24535 7364 24860 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 24946 7352 24952 7404
rect 25004 7392 25010 7404
rect 25004 7364 25049 7392
rect 25004 7352 25010 7364
rect 28166 7352 28172 7404
rect 28224 7392 28230 7404
rect 28353 7395 28411 7401
rect 28353 7392 28365 7395
rect 28224 7364 28365 7392
rect 28224 7352 28230 7364
rect 28353 7361 28365 7364
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 28997 7395 29055 7401
rect 28997 7361 29009 7395
rect 29043 7392 29055 7395
rect 29178 7392 29184 7404
rect 29043 7364 29184 7392
rect 29043 7361 29055 7364
rect 28997 7355 29055 7361
rect 29178 7352 29184 7364
rect 29236 7352 29242 7404
rect 29641 7395 29699 7401
rect 29641 7392 29653 7395
rect 29288 7364 29653 7392
rect 18414 7324 18420 7336
rect 17604 7296 18420 7324
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 22002 7324 22008 7336
rect 18800 7296 20024 7324
rect 21963 7296 22008 7324
rect 9401 7259 9459 7265
rect 9401 7225 9413 7259
rect 9447 7256 9459 7259
rect 11885 7259 11943 7265
rect 9447 7228 9674 7256
rect 9447 7225 9459 7228
rect 9401 7219 9459 7225
rect 9646 7188 9674 7228
rect 11885 7225 11897 7259
rect 11931 7256 11943 7259
rect 12066 7256 12072 7268
rect 11931 7228 12072 7256
rect 11931 7225 11943 7228
rect 11885 7219 11943 7225
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 15620 7228 15853 7256
rect 15620 7216 15626 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 15841 7219 15899 7225
rect 17497 7259 17555 7265
rect 17497 7225 17509 7259
rect 17543 7256 17555 7259
rect 18800 7256 18828 7296
rect 17543 7228 18828 7256
rect 19996 7256 20024 7296
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 26142 7324 26148 7336
rect 26103 7296 26148 7324
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 26513 7327 26571 7333
rect 26513 7293 26525 7327
rect 26559 7324 26571 7327
rect 27801 7327 27859 7333
rect 27801 7324 27813 7327
rect 26559 7296 27813 7324
rect 26559 7293 26571 7296
rect 26513 7287 26571 7293
rect 27801 7293 27813 7296
rect 27847 7324 27859 7327
rect 28902 7324 28908 7336
rect 27847 7296 28908 7324
rect 27847 7293 27859 7296
rect 27801 7287 27859 7293
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 21542 7256 21548 7268
rect 19996 7228 21548 7256
rect 17543 7225 17555 7228
rect 17497 7219 17555 7225
rect 21542 7216 21548 7228
rect 21600 7216 21606 7268
rect 23474 7216 23480 7268
rect 23532 7256 23538 7268
rect 23842 7256 23848 7268
rect 23532 7228 23848 7256
rect 23532 7216 23538 7228
rect 23842 7216 23848 7228
rect 23900 7256 23906 7268
rect 24762 7256 24768 7268
rect 23900 7228 24768 7256
rect 23900 7216 23906 7228
rect 24762 7216 24768 7228
rect 24820 7216 24826 7268
rect 27338 7216 27344 7268
rect 27396 7256 27402 7268
rect 29288 7256 29316 7364
rect 29641 7361 29653 7364
rect 29687 7361 29699 7395
rect 29641 7355 29699 7361
rect 30469 7395 30527 7401
rect 30469 7361 30481 7395
rect 30515 7392 30527 7395
rect 31110 7392 31116 7404
rect 30515 7364 31116 7392
rect 30515 7361 30527 7364
rect 30469 7355 30527 7361
rect 31110 7352 31116 7364
rect 31168 7352 31174 7404
rect 35894 7352 35900 7404
rect 35952 7392 35958 7404
rect 38013 7395 38071 7401
rect 38013 7392 38025 7395
rect 35952 7364 38025 7392
rect 35952 7352 35958 7364
rect 38013 7361 38025 7364
rect 38059 7361 38071 7395
rect 38013 7355 38071 7361
rect 38286 7324 38292 7336
rect 38247 7296 38292 7324
rect 38286 7284 38292 7296
rect 38344 7284 38350 7336
rect 31018 7256 31024 7268
rect 27396 7228 29316 7256
rect 30979 7228 31024 7256
rect 27396 7216 27402 7228
rect 31018 7216 31024 7228
rect 31076 7216 31082 7268
rect 31570 7216 31576 7268
rect 31628 7256 31634 7268
rect 31665 7259 31723 7265
rect 31665 7256 31677 7259
rect 31628 7228 31677 7256
rect 31628 7216 31634 7228
rect 31665 7225 31677 7228
rect 31711 7256 31723 7259
rect 32582 7256 32588 7268
rect 31711 7228 32588 7256
rect 31711 7225 31723 7228
rect 31665 7219 31723 7225
rect 32582 7216 32588 7228
rect 32640 7216 32646 7268
rect 10226 7188 10232 7200
rect 9646 7160 10232 7188
rect 10226 7148 10232 7160
rect 10284 7188 10290 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10284 7160 10425 7188
rect 10284 7148 10290 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 18598 7188 18604 7200
rect 12216 7160 18604 7188
rect 12216 7148 12222 7160
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19426 7188 19432 7200
rect 18748 7160 19432 7188
rect 18748 7148 18754 7160
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 21082 7188 21088 7200
rect 19576 7160 21088 7188
rect 19576 7148 19582 7160
rect 21082 7148 21088 7160
rect 21140 7188 21146 7200
rect 22370 7188 22376 7200
rect 21140 7160 22376 7188
rect 21140 7148 21146 7160
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 23382 7148 23388 7200
rect 23440 7188 23446 7200
rect 27890 7188 27896 7200
rect 23440 7160 27896 7188
rect 23440 7148 23446 7160
rect 27890 7148 27896 7160
rect 27948 7148 27954 7200
rect 28074 7148 28080 7200
rect 28132 7188 28138 7200
rect 28534 7188 28540 7200
rect 28132 7160 28540 7188
rect 28132 7148 28138 7160
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 32214 7148 32220 7200
rect 32272 7188 32278 7200
rect 32309 7191 32367 7197
rect 32309 7188 32321 7191
rect 32272 7160 32321 7188
rect 32272 7148 32278 7160
rect 32309 7157 32321 7160
rect 32355 7157 32367 7191
rect 32309 7151 32367 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 14642 6984 14648 6996
rect 14384 6956 14648 6984
rect 12529 6919 12587 6925
rect 12529 6885 12541 6919
rect 12575 6916 12587 6919
rect 14384 6916 14412 6956
rect 14642 6944 14648 6956
rect 14700 6984 14706 6996
rect 16390 6984 16396 6996
rect 14700 6956 16396 6984
rect 14700 6944 14706 6956
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 17402 6993 17408 6996
rect 17392 6987 17408 6993
rect 17392 6953 17404 6987
rect 17392 6947 17408 6953
rect 17402 6944 17408 6947
rect 17460 6944 17466 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 19518 6984 19524 6996
rect 18564 6956 19524 6984
rect 18564 6944 18570 6956
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 19692 6987 19750 6993
rect 19692 6953 19704 6987
rect 19738 6984 19750 6987
rect 20254 6984 20260 6996
rect 19738 6956 20260 6984
rect 19738 6953 19750 6956
rect 19692 6947 19750 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 21324 6956 21833 6984
rect 21324 6944 21330 6956
rect 21821 6953 21833 6956
rect 21867 6984 21879 6987
rect 21867 6956 24624 6984
rect 21867 6953 21879 6956
rect 21821 6947 21879 6953
rect 16298 6916 16304 6928
rect 12575 6888 12664 6916
rect 12575 6885 12587 6888
rect 12529 6879 12587 6885
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 12636 6848 12664 6888
rect 13464 6888 14412 6916
rect 15580 6888 16304 6916
rect 13464 6848 13492 6888
rect 13630 6848 13636 6860
rect 11471 6820 12572 6848
rect 12636 6820 13492 6848
rect 13591 6820 13636 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 12434 6780 12440 6792
rect 9815 6752 12440 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 12544 6780 12572 6820
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14148 6820 14289 6848
rect 14148 6808 14154 6820
rect 14277 6817 14289 6820
rect 14323 6848 14335 6851
rect 14550 6848 14556 6860
rect 14323 6820 14556 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15580 6848 15608 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 24596 6916 24624 6956
rect 24670 6944 24676 6996
rect 24728 6984 24734 6996
rect 27062 6984 27068 6996
rect 24728 6956 27068 6984
rect 24728 6944 24734 6956
rect 27062 6944 27068 6956
rect 27120 6944 27126 6996
rect 27154 6944 27160 6996
rect 27212 6984 27218 6996
rect 27212 6956 27568 6984
rect 27212 6944 27218 6956
rect 27246 6916 27252 6928
rect 24596 6888 27252 6916
rect 15068 6820 15608 6848
rect 15068 6808 15074 6820
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15896 6820 16037 6848
rect 15896 6808 15902 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16025 6811 16083 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6848 17187 6851
rect 19426 6848 19432 6860
rect 17175 6820 19432 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 23290 6848 23296 6860
rect 22112 6820 23296 6848
rect 13541 6783 13599 6789
rect 12544 6752 13124 6780
rect 9122 6712 9128 6724
rect 9035 6684 9128 6712
rect 9122 6672 9128 6684
rect 9180 6712 9186 6724
rect 10778 6712 10784 6724
rect 9180 6684 10784 6712
rect 9180 6672 9186 6684
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 13096 6712 13124 6752
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13587 6752 14136 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13998 6712 14004 6724
rect 13096 6684 14004 6712
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14108 6712 14136 6752
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 16448 6752 16497 6780
rect 16448 6740 16454 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 22112 6780 22140 6820
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 23569 6851 23627 6857
rect 23569 6817 23581 6851
rect 23615 6848 23627 6851
rect 23750 6848 23756 6860
rect 23615 6820 23756 6848
rect 23615 6817 23627 6820
rect 23569 6811 23627 6817
rect 23750 6808 23756 6820
rect 23808 6848 23814 6860
rect 24210 6848 24216 6860
rect 23808 6820 24216 6848
rect 23808 6808 23814 6820
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 24596 6848 24624 6888
rect 27246 6876 27252 6888
rect 27304 6876 27310 6928
rect 27540 6916 27568 6956
rect 27798 6944 27804 6996
rect 27856 6984 27862 6996
rect 28718 6984 28724 6996
rect 27856 6956 28724 6984
rect 27856 6944 27862 6956
rect 28718 6944 28724 6956
rect 28776 6944 28782 6996
rect 29178 6944 29184 6996
rect 29236 6984 29242 6996
rect 29825 6987 29883 6993
rect 29825 6984 29837 6987
rect 29236 6956 29837 6984
rect 29236 6944 29242 6956
rect 29825 6953 29837 6956
rect 29871 6953 29883 6987
rect 29825 6947 29883 6953
rect 28905 6919 28963 6925
rect 28905 6916 28917 6919
rect 27540 6888 28917 6916
rect 28905 6885 28917 6888
rect 28951 6885 28963 6919
rect 38286 6916 38292 6928
rect 28905 6879 28963 6885
rect 29288 6888 29408 6916
rect 38247 6888 38292 6916
rect 24596 6820 24716 6848
rect 20838 6752 22140 6780
rect 16485 6743 16543 6749
rect 23658 6740 23664 6792
rect 23716 6780 23722 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 23716 6752 24593 6780
rect 23716 6740 23722 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 24688 6780 24716 6820
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 27801 6851 27859 6857
rect 27801 6848 27813 6851
rect 24820 6820 27813 6848
rect 24820 6808 24826 6820
rect 27801 6817 27813 6820
rect 27847 6848 27859 6851
rect 29288 6848 29316 6888
rect 27847 6820 29316 6848
rect 29380 6848 29408 6888
rect 38286 6876 38292 6888
rect 38344 6876 38350 6928
rect 31570 6848 31576 6860
rect 29380 6820 31576 6848
rect 27847 6817 27859 6820
rect 27801 6811 27859 6817
rect 31570 6808 31576 6820
rect 31628 6808 31634 6860
rect 25314 6780 25320 6792
rect 24688 6752 25176 6780
rect 25275 6752 25320 6780
rect 24581 6743 24639 6749
rect 14108 6684 14412 6712
rect 14384 6656 14412 6684
rect 14458 6672 14464 6724
rect 14516 6712 14522 6724
rect 14553 6715 14611 6721
rect 14553 6712 14565 6715
rect 14516 6684 14565 6712
rect 14516 6672 14522 6684
rect 14553 6681 14565 6684
rect 14599 6712 14611 6715
rect 14826 6712 14832 6724
rect 14599 6684 14832 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 17310 6712 17316 6724
rect 15778 6684 17316 6712
rect 17310 6672 17316 6684
rect 17368 6672 17374 6724
rect 18630 6684 19656 6712
rect 10226 6644 10232 6656
rect 10187 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 11885 6647 11943 6653
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 12526 6644 12532 6656
rect 11931 6616 12532 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12526 6604 12532 6616
rect 12584 6644 12590 6656
rect 13078 6644 13084 6656
rect 12584 6616 13084 6644
rect 12584 6604 12590 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14366 6604 14372 6656
rect 14424 6604 14430 6656
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 18966 6644 18972 6656
rect 18923 6616 18972 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 19628 6644 19656 6684
rect 22830 6672 22836 6724
rect 22888 6672 22894 6724
rect 23198 6672 23204 6724
rect 23256 6712 23262 6724
rect 23293 6715 23351 6721
rect 23293 6712 23305 6715
rect 23256 6684 23305 6712
rect 23256 6672 23262 6684
rect 23293 6681 23305 6684
rect 23339 6681 23351 6715
rect 23293 6675 23351 6681
rect 24394 6672 24400 6724
rect 24452 6712 24458 6724
rect 24673 6715 24731 6721
rect 24673 6712 24685 6715
rect 24452 6684 24685 6712
rect 24452 6672 24458 6684
rect 24673 6681 24685 6684
rect 24719 6681 24731 6715
rect 25148 6712 25176 6752
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 25424 6712 25452 6743
rect 26694 6740 26700 6792
rect 26752 6780 26758 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 26752 6752 27169 6780
rect 26752 6740 26758 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 27246 6740 27252 6792
rect 27304 6780 27310 6792
rect 27304 6752 27349 6780
rect 27304 6740 27310 6752
rect 27706 6740 27712 6792
rect 27764 6780 27770 6792
rect 28074 6780 28080 6792
rect 27764 6752 28080 6780
rect 27764 6740 27770 6752
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 29178 6782 29184 6792
rect 29104 6780 29184 6782
rect 29012 6754 29184 6780
rect 29012 6752 29132 6754
rect 25148 6684 25452 6712
rect 25869 6715 25927 6721
rect 24673 6675 24731 6681
rect 25869 6681 25881 6715
rect 25915 6712 25927 6715
rect 26142 6712 26148 6724
rect 25915 6684 26148 6712
rect 25915 6681 25927 6684
rect 25869 6675 25927 6681
rect 26142 6672 26148 6684
rect 26200 6672 26206 6724
rect 26418 6712 26424 6724
rect 26379 6684 26424 6712
rect 26418 6672 26424 6684
rect 26476 6672 26482 6724
rect 26510 6672 26516 6724
rect 26568 6712 26574 6724
rect 28350 6712 28356 6724
rect 26568 6684 28356 6712
rect 26568 6672 26574 6684
rect 28350 6672 28356 6684
rect 28408 6672 28414 6724
rect 28442 6672 28448 6724
rect 28500 6712 28506 6724
rect 28500 6684 28545 6712
rect 28500 6672 28506 6684
rect 28810 6672 28816 6724
rect 28868 6712 28874 6724
rect 29012 6712 29040 6752
rect 29178 6740 29184 6754
rect 29236 6740 29242 6792
rect 29362 6740 29368 6792
rect 29420 6780 29426 6792
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 29420 6752 29929 6780
rect 29420 6740 29426 6752
rect 29917 6749 29929 6752
rect 29963 6780 29975 6783
rect 30561 6783 30619 6789
rect 30561 6780 30573 6783
rect 29963 6752 30573 6780
rect 29963 6749 29975 6752
rect 29917 6743 29975 6749
rect 30561 6749 30573 6752
rect 30607 6749 30619 6783
rect 30561 6743 30619 6749
rect 28868 6684 29040 6712
rect 30576 6712 30604 6743
rect 31110 6740 31116 6792
rect 31168 6740 31174 6792
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6780 31263 6783
rect 31294 6780 31300 6792
rect 31251 6752 31300 6780
rect 31251 6749 31263 6752
rect 31205 6743 31263 6749
rect 31294 6740 31300 6752
rect 31352 6780 31358 6792
rect 31849 6783 31907 6789
rect 31849 6780 31861 6783
rect 31352 6752 31861 6780
rect 31352 6740 31358 6752
rect 31849 6749 31861 6752
rect 31895 6780 31907 6783
rect 32490 6780 32496 6792
rect 31895 6752 32496 6780
rect 31895 6749 31907 6752
rect 31849 6743 31907 6749
rect 32490 6740 32496 6752
rect 32548 6740 32554 6792
rect 31128 6712 31156 6740
rect 30576 6684 31892 6712
rect 28868 6672 28874 6684
rect 31864 6656 31892 6684
rect 20714 6644 20720 6656
rect 19628 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 21174 6644 21180 6656
rect 21135 6616 21180 6644
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 22278 6604 22284 6656
rect 22336 6644 22342 6656
rect 29178 6644 29184 6656
rect 22336 6616 29184 6644
rect 22336 6604 22342 6616
rect 29178 6604 29184 6616
rect 29236 6604 29242 6656
rect 30466 6644 30472 6656
rect 30427 6616 30472 6644
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 31110 6644 31116 6656
rect 31071 6616 31116 6644
rect 31110 6604 31116 6616
rect 31168 6604 31174 6656
rect 31202 6604 31208 6656
rect 31260 6644 31266 6656
rect 31757 6647 31815 6653
rect 31757 6644 31769 6647
rect 31260 6616 31769 6644
rect 31260 6604 31266 6616
rect 31757 6613 31769 6616
rect 31803 6613 31815 6647
rect 31757 6607 31815 6613
rect 31846 6604 31852 6656
rect 31904 6604 31910 6656
rect 32401 6647 32459 6653
rect 32401 6613 32413 6647
rect 32447 6644 32459 6647
rect 32582 6644 32588 6656
rect 32447 6616 32588 6644
rect 32447 6613 32459 6616
rect 32401 6607 32459 6613
rect 32582 6604 32588 6616
rect 32640 6604 32646 6656
rect 32858 6644 32864 6656
rect 32819 6616 32864 6644
rect 32858 6604 32864 6616
rect 32916 6604 32922 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 33413 6647 33471 6653
rect 33413 6644 33425 6647
rect 33376 6616 33425 6644
rect 33376 6604 33382 6616
rect 33413 6613 33425 6616
rect 33459 6613 33471 6647
rect 33962 6644 33968 6656
rect 33923 6616 33968 6644
rect 33413 6607 33471 6613
rect 33962 6604 33968 6616
rect 34020 6604 34026 6656
rect 37642 6644 37648 6656
rect 37603 6616 37648 6644
rect 37642 6604 37648 6616
rect 37700 6604 37706 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 8294 6440 8300 6452
rect 4571 6412 8300 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10870 6440 10876 6452
rect 10643 6412 10876 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 13446 6440 13452 6452
rect 11756 6412 13452 6440
rect 11756 6400 11762 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 14056 6412 14964 6440
rect 14056 6400 14062 6412
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 13722 6372 13728 6384
rect 4672 6344 13728 6372
rect 4672 6332 4678 6344
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 14936 6372 14964 6412
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15804 6412 16221 6440
rect 15804 6400 15810 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16209 6403 16267 6409
rect 16482 6400 16488 6452
rect 16540 6440 16546 6452
rect 24026 6440 24032 6452
rect 16540 6412 24032 6440
rect 16540 6400 16546 6412
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 27706 6440 27712 6452
rect 24872 6412 27712 6440
rect 14936 6344 16252 6372
rect 16224 6316 16252 6344
rect 17862 6332 17868 6384
rect 17920 6332 17926 6384
rect 19426 6372 19432 6384
rect 19260 6344 19432 6372
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4120 6276 4445 6304
rect 4120 6264 4126 6276
rect 4433 6273 4445 6276
rect 4479 6304 4491 6307
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4479 6276 5181 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 5169 6273 5181 6276
rect 5215 6304 5227 6307
rect 8018 6304 8024 6316
rect 5215 6276 8024 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 8018 6264 8024 6276
rect 8076 6304 8082 6316
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 8076 6276 8125 6304
rect 8076 6264 8082 6276
rect 8113 6273 8125 6276
rect 8159 6304 8171 6307
rect 9122 6304 9128 6316
rect 8159 6276 9128 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9272 6276 14214 6304
rect 9272 6264 9278 6276
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 16117 6307 16175 6313
rect 16117 6304 16129 6307
rect 16080 6276 16129 6304
rect 16080 6264 16086 6276
rect 16117 6273 16129 6276
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 19260 6313 19288 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 19521 6375 19579 6381
rect 19521 6341 19533 6375
rect 19567 6372 19579 6375
rect 19794 6372 19800 6384
rect 19567 6344 19800 6372
rect 19567 6341 19579 6344
rect 19521 6335 19579 6341
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 22278 6372 22284 6384
rect 20746 6344 22284 6372
rect 22278 6332 22284 6344
rect 22336 6332 22342 6384
rect 24872 6372 24900 6412
rect 27706 6400 27712 6412
rect 27764 6400 27770 6452
rect 27890 6440 27896 6452
rect 27851 6412 27896 6440
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 28626 6440 28632 6452
rect 28587 6412 28632 6440
rect 28626 6400 28632 6412
rect 28684 6400 28690 6452
rect 28718 6400 28724 6452
rect 28776 6440 28782 6452
rect 30742 6440 30748 6452
rect 28776 6412 30748 6440
rect 28776 6400 28782 6412
rect 23506 6344 24900 6372
rect 26513 6375 26571 6381
rect 26513 6341 26525 6375
rect 26559 6372 26571 6375
rect 26878 6372 26884 6384
rect 26559 6344 26884 6372
rect 26559 6341 26571 6344
rect 26513 6335 26571 6341
rect 26878 6332 26884 6344
rect 26936 6332 26942 6384
rect 27062 6332 27068 6384
rect 27120 6372 27126 6384
rect 27249 6375 27307 6381
rect 27249 6372 27261 6375
rect 27120 6344 27261 6372
rect 27120 6332 27126 6344
rect 27249 6341 27261 6344
rect 27295 6341 27307 6375
rect 30116 6372 30144 6412
rect 30742 6400 30748 6412
rect 30800 6440 30806 6452
rect 32398 6440 32404 6452
rect 30800 6412 31340 6440
rect 32359 6412 32404 6440
rect 30800 6400 30806 6412
rect 30558 6372 30564 6384
rect 27249 6335 27307 6341
rect 28000 6344 29408 6372
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 18831 6276 19257 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 24210 6304 24216 6316
rect 24171 6276 24216 6304
rect 19245 6267 19303 6273
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 13630 6236 13636 6248
rect 10520 6208 13636 6236
rect 8573 6171 8631 6177
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 10520 6168 10548 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 14550 6236 14556 6248
rect 13740 6208 14556 6236
rect 8619 6140 10548 6168
rect 11149 6171 11207 6177
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 11149 6137 11161 6171
rect 11195 6168 11207 6171
rect 11974 6168 11980 6180
rect 11195 6140 11980 6168
rect 11195 6137 11207 6140
rect 11149 6131 11207 6137
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9766 6100 9772 6112
rect 9263 6072 9772 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10045 6103 10103 6109
rect 10045 6069 10057 6103
rect 10091 6100 10103 6103
rect 10226 6100 10232 6112
rect 10091 6072 10232 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10226 6060 10232 6072
rect 10284 6100 10290 6112
rect 11164 6100 11192 6131
rect 11974 6128 11980 6140
rect 12032 6168 12038 6180
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 12032 6140 12173 6168
rect 12032 6128 12038 6140
rect 12161 6137 12173 6140
rect 12207 6168 12219 6171
rect 12713 6171 12771 6177
rect 12713 6168 12725 6171
rect 12207 6140 12725 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12713 6137 12725 6140
rect 12759 6168 12771 6171
rect 13078 6168 13084 6180
rect 12759 6140 13084 6168
rect 12759 6137 12771 6140
rect 12713 6131 12771 6137
rect 13078 6128 13084 6140
rect 13136 6168 13142 6180
rect 13265 6171 13323 6177
rect 13265 6168 13277 6171
rect 13136 6140 13277 6168
rect 13136 6128 13142 6140
rect 13265 6137 13277 6140
rect 13311 6168 13323 6171
rect 13740 6168 13768 6208
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 14700 6208 15301 6236
rect 14700 6196 14706 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 15746 6236 15752 6248
rect 15611 6208 15752 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 17420 6208 18521 6236
rect 17420 6180 17448 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 18966 6196 18972 6248
rect 19024 6236 19030 6248
rect 21358 6236 21364 6248
rect 19024 6208 21364 6236
rect 19024 6196 19030 6208
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 22002 6236 22008 6248
rect 21963 6208 22008 6236
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 22278 6236 22284 6248
rect 22239 6208 22284 6236
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22370 6196 22376 6248
rect 22428 6236 22434 6248
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 22428 6208 24501 6236
rect 22428 6196 22434 6208
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 25608 6236 25636 6290
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 26292 6276 26433 6304
rect 26292 6264 26298 6276
rect 26421 6273 26433 6276
rect 26467 6304 26479 6307
rect 26694 6304 26700 6316
rect 26467 6276 26700 6304
rect 26467 6273 26479 6276
rect 26421 6267 26479 6273
rect 26694 6264 26700 6276
rect 26752 6264 26758 6316
rect 28000 6313 28028 6344
rect 29380 6316 29408 6344
rect 30024 6344 30144 6372
rect 30519 6344 30564 6372
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6304 27399 6307
rect 27985 6307 28043 6313
rect 27985 6304 27997 6307
rect 27387 6276 27997 6304
rect 27387 6273 27399 6276
rect 27341 6267 27399 6273
rect 27985 6273 27997 6276
rect 28031 6273 28043 6307
rect 28718 6304 28724 6316
rect 28679 6276 28724 6304
rect 27985 6267 28043 6273
rect 28718 6264 28724 6276
rect 28776 6264 28782 6316
rect 29362 6304 29368 6316
rect 29323 6276 29368 6304
rect 29362 6264 29368 6276
rect 29420 6264 29426 6316
rect 30024 6313 30052 6344
rect 30558 6332 30564 6344
rect 30616 6332 30622 6384
rect 30009 6307 30067 6313
rect 30009 6273 30021 6307
rect 30055 6273 30067 6307
rect 30009 6267 30067 6273
rect 30098 6264 30104 6316
rect 30156 6304 30162 6316
rect 30653 6307 30711 6313
rect 30653 6304 30665 6307
rect 30156 6276 30665 6304
rect 30156 6264 30162 6276
rect 30653 6273 30665 6276
rect 30699 6304 30711 6307
rect 31202 6304 31208 6316
rect 30699 6276 31208 6304
rect 30699 6273 30711 6276
rect 30653 6267 30711 6273
rect 31202 6264 31208 6276
rect 31260 6264 31266 6316
rect 31312 6313 31340 6412
rect 32398 6400 32404 6412
rect 32456 6400 32462 6452
rect 31297 6307 31355 6313
rect 31297 6273 31309 6307
rect 31343 6304 31355 6307
rect 31386 6304 31392 6316
rect 31343 6276 31392 6304
rect 31343 6273 31355 6276
rect 31297 6267 31355 6273
rect 31386 6264 31392 6276
rect 31444 6264 31450 6316
rect 32490 6304 32496 6316
rect 32451 6276 32496 6304
rect 32490 6264 32496 6276
rect 32548 6264 32554 6316
rect 27430 6236 27436 6248
rect 25608 6208 27436 6236
rect 24489 6199 24547 6205
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 31754 6236 31760 6248
rect 27764 6208 31760 6236
rect 27764 6196 27770 6208
rect 31754 6196 31760 6208
rect 31812 6196 31818 6248
rect 13311 6140 13768 6168
rect 13311 6137 13323 6140
rect 13265 6131 13323 6137
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 16482 6168 16488 6180
rect 15988 6140 16488 6168
rect 15988 6128 15994 6140
rect 16482 6128 16488 6140
rect 16540 6168 16546 6180
rect 17037 6171 17095 6177
rect 17037 6168 17049 6171
rect 16540 6140 17049 6168
rect 16540 6128 16546 6140
rect 17037 6137 17049 6140
rect 17083 6137 17095 6171
rect 17037 6131 17095 6137
rect 17402 6128 17408 6180
rect 17460 6128 17466 6180
rect 20993 6171 21051 6177
rect 20993 6137 21005 6171
rect 21039 6168 21051 6171
rect 21039 6140 22140 6168
rect 21039 6137 21051 6140
rect 20993 6131 21051 6137
rect 10284 6072 11192 6100
rect 10284 6060 10290 6072
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13504 6072 13829 6100
rect 13504 6060 13510 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 17310 6060 17316 6112
rect 17368 6100 17374 6112
rect 21726 6100 21732 6112
rect 17368 6072 21732 6100
rect 17368 6060 17374 6072
rect 21726 6060 21732 6072
rect 21784 6060 21790 6112
rect 22112 6100 22140 6140
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 23753 6171 23811 6177
rect 23753 6168 23765 6171
rect 23532 6140 23765 6168
rect 23532 6128 23538 6140
rect 23753 6137 23765 6140
rect 23799 6137 23811 6171
rect 29917 6171 29975 6177
rect 29917 6168 29929 6171
rect 23753 6131 23811 6137
rect 25792 6140 29929 6168
rect 22370 6100 22376 6112
rect 22112 6072 22376 6100
rect 22370 6060 22376 6072
rect 22428 6100 22434 6112
rect 23658 6100 23664 6112
rect 22428 6072 23664 6100
rect 22428 6060 22434 6072
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 25792 6100 25820 6140
rect 29917 6137 29929 6140
rect 29963 6137 29975 6171
rect 29917 6131 29975 6137
rect 32582 6128 32588 6180
rect 32640 6168 32646 6180
rect 33045 6171 33103 6177
rect 33045 6168 33057 6171
rect 32640 6140 33057 6168
rect 32640 6128 32646 6140
rect 33045 6137 33057 6140
rect 33091 6168 33103 6171
rect 33686 6168 33692 6180
rect 33091 6140 33692 6168
rect 33091 6137 33103 6140
rect 33045 6131 33103 6137
rect 33686 6128 33692 6140
rect 33744 6128 33750 6180
rect 25958 6100 25964 6112
rect 24084 6072 25820 6100
rect 25919 6072 25964 6100
rect 24084 6060 24090 6072
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 26050 6060 26056 6112
rect 26108 6100 26114 6112
rect 26510 6100 26516 6112
rect 26108 6072 26516 6100
rect 26108 6060 26114 6072
rect 26510 6060 26516 6072
rect 26568 6060 26574 6112
rect 26786 6060 26792 6112
rect 26844 6100 26850 6112
rect 29273 6103 29331 6109
rect 29273 6100 29285 6103
rect 26844 6072 29285 6100
rect 26844 6060 26850 6072
rect 29273 6069 29285 6072
rect 29319 6069 29331 6103
rect 29273 6063 29331 6069
rect 29638 6060 29644 6112
rect 29696 6100 29702 6112
rect 31205 6103 31263 6109
rect 31205 6100 31217 6103
rect 29696 6072 31217 6100
rect 29696 6060 29702 6072
rect 31205 6069 31217 6072
rect 31251 6069 31263 6103
rect 31205 6063 31263 6069
rect 33318 6060 33324 6112
rect 33376 6100 33382 6112
rect 33505 6103 33563 6109
rect 33505 6100 33517 6103
rect 33376 6072 33517 6100
rect 33376 6060 33382 6072
rect 33505 6069 33517 6072
rect 33551 6100 33563 6103
rect 34057 6103 34115 6109
rect 34057 6100 34069 6103
rect 33551 6072 34069 6100
rect 33551 6069 33563 6072
rect 33505 6063 33563 6069
rect 34057 6069 34069 6072
rect 34103 6069 34115 6103
rect 34057 6063 34115 6069
rect 36446 6060 36452 6112
rect 36504 6100 36510 6112
rect 37461 6103 37519 6109
rect 37461 6100 37473 6103
rect 36504 6072 37473 6100
rect 36504 6060 36510 6072
rect 37461 6069 37473 6072
rect 37507 6069 37519 6103
rect 38286 6100 38292 6112
rect 38247 6072 38292 6100
rect 37461 6063 37519 6069
rect 38286 6060 38292 6072
rect 38344 6060 38350 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5896 4215 5899
rect 4614 5896 4620 5908
rect 4203 5868 4620 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 10045 5899 10103 5905
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 10318 5896 10324 5908
rect 10091 5868 10324 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 10318 5856 10324 5868
rect 10376 5896 10382 5908
rect 14642 5896 14648 5908
rect 10376 5868 14648 5896
rect 10376 5856 10382 5868
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 16298 5896 16304 5908
rect 16259 5868 16304 5896
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17460 5868 19288 5896
rect 17460 5856 17466 5868
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 9214 5828 9220 5840
rect 3375 5800 9220 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5828 13783 5831
rect 13814 5828 13820 5840
rect 13771 5800 13820 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 18874 5828 18880 5840
rect 18835 5800 18880 5828
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 19260 5828 19288 5868
rect 19334 5856 19340 5908
rect 19392 5896 19398 5908
rect 19521 5899 19579 5905
rect 19521 5896 19533 5899
rect 19392 5868 19533 5896
rect 19392 5856 19398 5868
rect 19521 5865 19533 5868
rect 19567 5865 19579 5899
rect 19521 5859 19579 5865
rect 23311 5899 23369 5905
rect 23311 5865 23323 5899
rect 23357 5896 23369 5899
rect 26326 5896 26332 5908
rect 23357 5868 26188 5896
rect 26287 5868 26332 5896
rect 23357 5865 23369 5868
rect 23311 5859 23369 5865
rect 20165 5831 20223 5837
rect 19260 5800 20116 5828
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 11698 5760 11704 5772
rect 10643 5732 11704 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 11698 5720 11704 5732
rect 11756 5760 11762 5772
rect 11974 5760 11980 5772
rect 11756 5732 11980 5760
rect 11756 5720 11762 5732
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 13906 5760 13912 5772
rect 12299 5732 13912 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14826 5760 14832 5772
rect 14739 5732 14832 5760
rect 14826 5720 14832 5732
rect 14884 5760 14890 5772
rect 16390 5760 16396 5772
rect 14884 5732 16396 5760
rect 14884 5720 14890 5732
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 17126 5760 17132 5772
rect 17039 5732 17132 5760
rect 17126 5720 17132 5732
rect 17184 5760 17190 5772
rect 19518 5760 19524 5772
rect 17184 5732 19524 5760
rect 17184 5720 17190 5732
rect 19518 5720 19524 5732
rect 19576 5760 19582 5772
rect 19576 5732 20024 5760
rect 19576 5720 19582 5732
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3602 5692 3608 5704
rect 3467 5664 3608 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3602 5652 3608 5664
rect 3660 5692 3666 5704
rect 4062 5692 4068 5704
rect 3660 5664 4068 5692
rect 3660 5652 3666 5664
rect 4062 5652 4068 5664
rect 4120 5692 4126 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4120 5664 4721 5692
rect 4120 5652 4126 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 14550 5692 14556 5704
rect 14463 5664 14556 5692
rect 11057 5655 11115 5661
rect 9490 5624 9496 5636
rect 9451 5596 9496 5624
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 11072 5624 11100 5655
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 19058 5652 19064 5704
rect 19116 5692 19122 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19116 5664 19441 5692
rect 19116 5652 19122 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 13630 5624 13636 5636
rect 10836 5596 12572 5624
rect 13478 5596 13636 5624
rect 10836 5584 10842 5596
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 12434 5556 12440 5568
rect 11195 5528 12440 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12544 5556 12572 5596
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 14366 5556 14372 5568
rect 12544 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14568 5556 14596 5652
rect 16054 5596 16436 5624
rect 15746 5556 15752 5568
rect 14568 5528 15752 5556
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 16408 5556 16436 5596
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16540 5596 17417 5624
rect 16540 5584 16546 5596
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 19334 5624 19340 5636
rect 18630 5596 19340 5624
rect 17405 5587 17463 5593
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 19996 5624 20024 5732
rect 20088 5701 20116 5800
rect 20165 5797 20177 5831
rect 20211 5828 20223 5831
rect 26160 5828 26188 5868
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 26418 5856 26424 5908
rect 26476 5896 26482 5908
rect 27525 5899 27583 5905
rect 27525 5896 27537 5899
rect 26476 5868 27537 5896
rect 26476 5856 26482 5868
rect 27525 5865 27537 5868
rect 27571 5865 27583 5899
rect 27525 5859 27583 5865
rect 28169 5899 28227 5905
rect 28169 5865 28181 5899
rect 28215 5896 28227 5899
rect 28258 5896 28264 5908
rect 28215 5868 28264 5896
rect 28215 5865 28227 5868
rect 28169 5859 28227 5865
rect 28258 5856 28264 5868
rect 28316 5856 28322 5908
rect 29546 5856 29552 5908
rect 29604 5896 29610 5908
rect 29825 5899 29883 5905
rect 29825 5896 29837 5899
rect 29604 5868 29837 5896
rect 29604 5856 29610 5868
rect 29825 5865 29837 5868
rect 29871 5865 29883 5899
rect 29825 5859 29883 5865
rect 30282 5856 30288 5908
rect 30340 5896 30346 5908
rect 30469 5899 30527 5905
rect 30469 5896 30481 5899
rect 30340 5868 30481 5896
rect 30340 5856 30346 5868
rect 30469 5865 30481 5868
rect 30515 5865 30527 5899
rect 30469 5859 30527 5865
rect 31018 5856 31024 5908
rect 31076 5896 31082 5908
rect 31113 5899 31171 5905
rect 31113 5896 31125 5899
rect 31076 5868 31125 5896
rect 31076 5856 31082 5868
rect 31113 5865 31125 5868
rect 31159 5865 31171 5899
rect 31113 5859 31171 5865
rect 31754 5856 31760 5908
rect 31812 5896 31818 5908
rect 35434 5896 35440 5908
rect 31812 5868 31857 5896
rect 35395 5868 35440 5896
rect 31812 5856 31818 5868
rect 35434 5856 35440 5868
rect 35492 5856 35498 5908
rect 26602 5828 26608 5840
rect 20211 5800 22094 5828
rect 26160 5800 26608 5828
rect 20211 5797 20223 5800
rect 20165 5791 20223 5797
rect 22066 5760 22094 5800
rect 26602 5788 26608 5800
rect 26660 5788 26666 5840
rect 26881 5831 26939 5837
rect 26881 5797 26893 5831
rect 26927 5828 26939 5831
rect 26970 5828 26976 5840
rect 26927 5800 26976 5828
rect 26927 5797 26939 5800
rect 26881 5791 26939 5797
rect 26970 5788 26976 5800
rect 27028 5788 27034 5840
rect 28074 5788 28080 5840
rect 28132 5828 28138 5840
rect 28813 5831 28871 5837
rect 28813 5828 28825 5831
rect 28132 5800 28825 5828
rect 28132 5788 28138 5800
rect 28813 5797 28825 5800
rect 28859 5797 28871 5831
rect 30374 5828 30380 5840
rect 28813 5791 28871 5797
rect 28920 5800 30380 5828
rect 22554 5760 22560 5772
rect 22066 5732 22560 5760
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 22646 5720 22652 5772
rect 22704 5760 22710 5772
rect 28920 5760 28948 5800
rect 30374 5788 30380 5800
rect 30432 5788 30438 5840
rect 37458 5788 37464 5840
rect 37516 5828 37522 5840
rect 38013 5831 38071 5837
rect 38013 5828 38025 5831
rect 37516 5800 38025 5828
rect 37516 5788 37522 5800
rect 38013 5797 38025 5800
rect 38059 5797 38071 5831
rect 38013 5791 38071 5797
rect 31110 5760 31116 5772
rect 22704 5732 28948 5760
rect 22704 5720 22710 5732
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5661 20131 5695
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20073 5655 20131 5661
rect 20180 5664 20913 5692
rect 20180 5624 20208 5664
rect 20901 5661 20913 5664
rect 20947 5692 20959 5695
rect 22002 5692 22008 5704
rect 20947 5664 22008 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 22002 5652 22008 5664
rect 22060 5652 22066 5704
rect 23569 5695 23627 5701
rect 23569 5661 23581 5695
rect 23615 5692 23627 5695
rect 24210 5692 24216 5704
rect 23615 5664 24216 5692
rect 23615 5661 23627 5664
rect 23569 5655 23627 5661
rect 24210 5652 24216 5664
rect 24268 5692 24274 5704
rect 24578 5692 24584 5704
rect 24268 5664 24584 5692
rect 24268 5652 24274 5664
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26789 5695 26847 5701
rect 26789 5692 26801 5695
rect 26292 5664 26801 5692
rect 26292 5652 26298 5664
rect 26789 5661 26801 5664
rect 26835 5661 26847 5695
rect 26789 5655 26847 5661
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5692 27675 5695
rect 27798 5692 27804 5704
rect 27663 5664 27804 5692
rect 27663 5661 27675 5664
rect 27617 5655 27675 5661
rect 27798 5652 27804 5664
rect 27856 5652 27862 5704
rect 28074 5692 28080 5704
rect 28035 5664 28080 5692
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 28920 5701 28948 5732
rect 29012 5732 31116 5760
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5661 28963 5695
rect 28905 5655 28963 5661
rect 19996 5596 20208 5624
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 21545 5627 21603 5633
rect 21545 5624 21557 5627
rect 20312 5596 21557 5624
rect 20312 5584 20318 5596
rect 21545 5593 21557 5596
rect 21591 5593 21603 5627
rect 21545 5587 21603 5593
rect 21726 5584 21732 5636
rect 21784 5624 21790 5636
rect 24486 5624 24492 5636
rect 21784 5596 22048 5624
rect 22862 5596 24492 5624
rect 21784 5584 21790 5596
rect 21910 5556 21916 5568
rect 16408 5528 21916 5556
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 22020 5556 22048 5596
rect 24486 5584 24492 5596
rect 24544 5584 24550 5636
rect 24854 5584 24860 5636
rect 24912 5624 24918 5636
rect 26142 5624 26148 5636
rect 24912 5596 24957 5624
rect 26082 5596 26148 5624
rect 24912 5584 24918 5596
rect 26142 5584 26148 5596
rect 26200 5584 26206 5636
rect 29012 5624 29040 5732
rect 31110 5720 31116 5732
rect 31168 5720 31174 5772
rect 29917 5695 29975 5701
rect 29917 5661 29929 5695
rect 29963 5692 29975 5695
rect 30098 5692 30104 5704
rect 29963 5664 30104 5692
rect 29963 5661 29975 5664
rect 29917 5655 29975 5661
rect 30098 5652 30104 5664
rect 30156 5652 30162 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 30561 5695 30619 5701
rect 30561 5692 30573 5695
rect 30524 5664 30573 5692
rect 30524 5652 30530 5664
rect 30561 5661 30573 5664
rect 30607 5692 30619 5695
rect 31205 5695 31263 5701
rect 31205 5692 31217 5695
rect 30607 5664 31217 5692
rect 30607 5661 30619 5664
rect 30561 5655 30619 5661
rect 31205 5661 31217 5664
rect 31251 5692 31263 5695
rect 31849 5695 31907 5701
rect 31849 5692 31861 5695
rect 31251 5664 31861 5692
rect 31251 5661 31263 5664
rect 31205 5655 31263 5661
rect 31849 5661 31861 5664
rect 31895 5661 31907 5695
rect 32490 5692 32496 5704
rect 32403 5664 32496 5692
rect 31849 5655 31907 5661
rect 32490 5652 32496 5664
rect 32548 5692 32554 5704
rect 32858 5692 32864 5704
rect 32548 5664 32864 5692
rect 32548 5652 32554 5664
rect 32858 5652 32864 5664
rect 32916 5652 32922 5704
rect 33137 5695 33195 5701
rect 33137 5661 33149 5695
rect 33183 5692 33195 5695
rect 33318 5692 33324 5704
rect 33183 5664 33324 5692
rect 33183 5661 33195 5664
rect 33137 5655 33195 5661
rect 33318 5652 33324 5664
rect 33376 5692 33382 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 33376 5664 34897 5692
rect 33376 5652 33382 5664
rect 34885 5661 34897 5664
rect 34931 5692 34943 5695
rect 35250 5692 35256 5704
rect 34931 5664 35256 5692
rect 34931 5661 34943 5664
rect 34885 5655 34943 5661
rect 35250 5652 35256 5664
rect 35308 5652 35314 5704
rect 26252 5596 29040 5624
rect 26252 5556 26280 5596
rect 30374 5584 30380 5636
rect 30432 5624 30438 5636
rect 32401 5627 32459 5633
rect 32401 5624 32413 5627
rect 30432 5596 32413 5624
rect 30432 5584 30438 5596
rect 32401 5593 32413 5596
rect 32447 5593 32459 5627
rect 32401 5587 32459 5593
rect 37553 5627 37611 5633
rect 37553 5593 37565 5627
rect 37599 5624 37611 5627
rect 38194 5624 38200 5636
rect 37599 5596 38200 5624
rect 37599 5593 37611 5596
rect 37553 5587 37611 5593
rect 38194 5584 38200 5596
rect 38252 5584 38258 5636
rect 22020 5528 26280 5556
rect 27430 5516 27436 5568
rect 27488 5556 27494 5568
rect 29730 5556 29736 5568
rect 27488 5528 29736 5556
rect 27488 5516 27494 5528
rect 29730 5516 29736 5528
rect 29788 5516 29794 5568
rect 33042 5556 33048 5568
rect 33003 5528 33048 5556
rect 33042 5516 33048 5528
rect 33100 5516 33106 5568
rect 33594 5556 33600 5568
rect 33555 5528 33600 5556
rect 33594 5516 33600 5528
rect 33652 5556 33658 5568
rect 34149 5559 34207 5565
rect 34149 5556 34161 5559
rect 33652 5528 34161 5556
rect 33652 5516 33658 5528
rect 34149 5525 34161 5528
rect 34195 5525 34207 5559
rect 36078 5556 36084 5568
rect 36039 5528 36084 5556
rect 34149 5519 34207 5525
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 36446 5516 36452 5568
rect 36504 5556 36510 5568
rect 36633 5559 36691 5565
rect 36633 5556 36645 5559
rect 36504 5528 36645 5556
rect 36504 5516 36510 5528
rect 36633 5525 36645 5528
rect 36679 5525 36691 5559
rect 36633 5519 36691 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3602 5352 3608 5364
rect 3563 5324 3608 5352
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10468 5324 10517 5352
rect 10468 5312 10474 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 12342 5352 12348 5364
rect 10505 5315 10563 5321
rect 11348 5324 12348 5352
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 11348 5284 11376 5324
rect 12342 5312 12348 5324
rect 12400 5352 12406 5364
rect 13449 5355 13507 5361
rect 12400 5324 13400 5352
rect 12400 5312 12406 5324
rect 7883 5256 11376 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 11882 5244 11888 5296
rect 11940 5284 11946 5296
rect 11977 5287 12035 5293
rect 11977 5284 11989 5287
rect 11940 5256 11989 5284
rect 11940 5244 11946 5256
rect 11977 5253 11989 5256
rect 12023 5253 12035 5287
rect 11977 5247 12035 5253
rect 12434 5244 12440 5296
rect 12492 5244 12498 5296
rect 13372 5284 13400 5324
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 16022 5352 16028 5364
rect 13495 5324 16028 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 16022 5312 16028 5324
rect 16080 5312 16086 5364
rect 16298 5312 16304 5364
rect 16356 5312 16362 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 19705 5355 19763 5361
rect 17368 5324 19288 5352
rect 17368 5312 17374 5324
rect 13372 5256 14044 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 1946 5216 1952 5228
rect 1903 5188 1952 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 10134 5216 10140 5228
rect 7331 5188 10140 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11698 5216 11704 5228
rect 11195 5188 11704 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 14016 5157 14044 5256
rect 15010 5244 15016 5296
rect 15068 5244 15074 5296
rect 15470 5284 15476 5296
rect 15383 5256 15476 5284
rect 15470 5244 15476 5256
rect 15528 5284 15534 5296
rect 16316 5284 16344 5312
rect 19260 5296 19288 5324
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 19886 5352 19892 5364
rect 19751 5324 19892 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 23842 5352 23848 5364
rect 23803 5324 23848 5352
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 24581 5355 24639 5361
rect 24581 5352 24593 5355
rect 23992 5324 24593 5352
rect 23992 5312 23998 5324
rect 24581 5321 24593 5324
rect 24627 5321 24639 5355
rect 25682 5352 25688 5364
rect 25643 5324 25688 5352
rect 24581 5315 24639 5321
rect 25682 5312 25688 5324
rect 25740 5312 25746 5364
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 27706 5312 27712 5364
rect 27764 5352 27770 5364
rect 27985 5355 28043 5361
rect 27985 5352 27997 5355
rect 27764 5324 27997 5352
rect 27764 5312 27770 5324
rect 27985 5321 27997 5324
rect 28031 5321 28043 5355
rect 27985 5315 28043 5321
rect 28442 5312 28448 5364
rect 28500 5352 28506 5364
rect 28629 5355 28687 5361
rect 28629 5352 28641 5355
rect 28500 5324 28641 5352
rect 28500 5312 28506 5324
rect 28629 5321 28641 5324
rect 28675 5321 28687 5355
rect 29914 5352 29920 5364
rect 29875 5324 29920 5352
rect 28629 5315 28687 5321
rect 29914 5312 29920 5324
rect 29972 5312 29978 5364
rect 30558 5352 30564 5364
rect 30519 5324 30564 5352
rect 30558 5312 30564 5324
rect 30616 5312 30622 5364
rect 34146 5352 34152 5364
rect 34107 5324 34152 5352
rect 34146 5312 34152 5324
rect 34204 5312 34210 5364
rect 35250 5352 35256 5364
rect 35211 5324 35256 5352
rect 35250 5312 35256 5324
rect 35308 5312 35314 5364
rect 19242 5284 19248 5296
rect 15528 5256 16344 5284
rect 19155 5256 19248 5284
rect 15528 5244 15534 5256
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 22646 5284 22652 5296
rect 20746 5256 22652 5284
rect 22646 5244 22652 5256
rect 22704 5244 22710 5296
rect 30374 5284 30380 5296
rect 23598 5256 25636 5284
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 15804 5188 16313 5216
rect 15804 5176 15810 5188
rect 16301 5185 16313 5188
rect 16347 5216 16359 5219
rect 17126 5216 17132 5228
rect 16347 5188 17132 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 17126 5176 17132 5188
rect 17184 5216 17190 5228
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 17184 5188 17233 5216
rect 17184 5176 17190 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 19794 5216 19800 5228
rect 18630 5188 19800 5216
rect 17221 5179 17279 5185
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 24670 5216 24676 5228
rect 24228 5188 24676 5216
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 14001 5151 14059 5157
rect 9539 5120 10916 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 8496 5052 9674 5080
rect 8496 5024 8524 5052
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 8076 4984 8309 5012
rect 8076 4972 8082 4984
rect 8297 4981 8309 4984
rect 8343 5012 8355 5015
rect 8478 5012 8484 5024
rect 8343 4984 8484 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8938 5012 8944 5024
rect 8899 4984 8944 5012
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9646 5012 9674 5052
rect 10042 5012 10048 5024
rect 9646 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10888 5012 10916 5120
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14182 5148 14188 5160
rect 14047 5120 14188 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14182 5108 14188 5120
rect 14240 5148 14246 5160
rect 15102 5148 15108 5160
rect 14240 5120 15108 5148
rect 14240 5108 14246 5120
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 17497 5151 17555 5157
rect 17497 5148 17509 5151
rect 15436 5120 15700 5148
rect 15436 5108 15442 5120
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 14274 5080 14280 5092
rect 13320 5052 14280 5080
rect 13320 5040 13326 5052
rect 14274 5040 14280 5052
rect 14332 5040 14338 5092
rect 15672 5080 15700 5120
rect 17328 5120 17509 5148
rect 17328 5080 17356 5120
rect 17497 5117 17509 5120
rect 17543 5117 17555 5151
rect 17497 5111 17555 5117
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5148 21235 5151
rect 21453 5151 21511 5157
rect 21223 5120 21404 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 15672 5052 17356 5080
rect 15470 5012 15476 5024
rect 10888 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 17328 5012 17356 5052
rect 19242 5040 19248 5092
rect 19300 5080 19306 5092
rect 19978 5080 19984 5092
rect 19300 5052 19984 5080
rect 19300 5040 19306 5052
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 21376 5080 21404 5120
rect 21453 5117 21465 5151
rect 21499 5148 21511 5151
rect 22094 5148 22100 5160
rect 21499 5120 22100 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 22094 5108 22100 5120
rect 22152 5108 22158 5160
rect 22370 5148 22376 5160
rect 22331 5120 22376 5148
rect 22370 5108 22376 5120
rect 22428 5108 22434 5160
rect 23014 5108 23020 5160
rect 23072 5148 23078 5160
rect 24228 5148 24256 5188
rect 24670 5176 24676 5188
rect 24728 5176 24734 5228
rect 25608 5216 25636 5256
rect 25792 5256 30380 5284
rect 25792 5216 25820 5256
rect 30374 5244 30380 5256
rect 30432 5244 30438 5296
rect 33045 5287 33103 5293
rect 33045 5284 33057 5287
rect 30760 5256 33057 5284
rect 25608 5188 25820 5216
rect 25866 5176 25872 5228
rect 25924 5216 25930 5228
rect 26421 5219 26479 5225
rect 25924 5188 25969 5216
rect 25924 5176 25930 5188
rect 26421 5185 26433 5219
rect 26467 5185 26479 5219
rect 26421 5179 26479 5185
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 27982 5216 27988 5228
rect 27387 5188 27988 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 23072 5120 24256 5148
rect 23072 5108 23078 5120
rect 21818 5080 21824 5092
rect 21376 5052 21824 5080
rect 21818 5040 21824 5052
rect 21876 5040 21882 5092
rect 20070 5012 20076 5024
rect 17328 4984 20076 5012
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 23566 5012 23572 5024
rect 22520 4984 23572 5012
rect 22520 4972 22526 4984
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 24578 4972 24584 5024
rect 24636 5012 24642 5024
rect 25133 5015 25191 5021
rect 25133 5012 25145 5015
rect 24636 4984 25145 5012
rect 24636 4972 24642 4984
rect 25133 4981 25145 4984
rect 25179 4981 25191 5015
rect 25133 4975 25191 4981
rect 25314 4972 25320 5024
rect 25372 5012 25378 5024
rect 26436 5012 26464 5179
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28077 5219 28135 5225
rect 28077 5185 28089 5219
rect 28123 5216 28135 5219
rect 28626 5216 28632 5228
rect 28123 5188 28632 5216
rect 28123 5185 28135 5188
rect 28077 5179 28135 5185
rect 28626 5176 28632 5188
rect 28684 5176 28690 5228
rect 28718 5176 28724 5228
rect 28776 5216 28782 5228
rect 28776 5188 28821 5216
rect 28776 5176 28782 5188
rect 29178 5176 29184 5228
rect 29236 5216 29242 5228
rect 29365 5219 29423 5225
rect 29365 5216 29377 5219
rect 29236 5188 29377 5216
rect 29236 5176 29242 5188
rect 29365 5185 29377 5188
rect 29411 5185 29423 5219
rect 29822 5216 29828 5228
rect 29783 5188 29828 5216
rect 29365 5179 29423 5185
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 30524 5188 30665 5216
rect 30524 5176 30530 5188
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 27614 5108 27620 5160
rect 27672 5148 27678 5160
rect 30760 5148 30788 5256
rect 33045 5253 33057 5256
rect 33091 5253 33103 5287
rect 33045 5247 33103 5253
rect 31202 5176 31208 5228
rect 31260 5216 31266 5228
rect 31297 5219 31355 5225
rect 31297 5216 31309 5219
rect 31260 5188 31309 5216
rect 31260 5176 31266 5188
rect 31297 5185 31309 5188
rect 31343 5185 31355 5219
rect 31297 5179 31355 5185
rect 31386 5176 31392 5228
rect 31444 5216 31450 5228
rect 32493 5219 32551 5225
rect 32493 5216 32505 5219
rect 31444 5188 32505 5216
rect 31444 5176 31450 5188
rect 32493 5185 32505 5188
rect 32539 5216 32551 5219
rect 32582 5216 32588 5228
rect 32539 5188 32588 5216
rect 32539 5185 32551 5188
rect 32493 5179 32551 5185
rect 32582 5176 32588 5188
rect 32640 5176 32646 5228
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5216 33195 5219
rect 33226 5216 33232 5228
rect 33183 5188 33232 5216
rect 33183 5185 33195 5188
rect 33137 5179 33195 5185
rect 33226 5176 33232 5188
rect 33284 5176 33290 5228
rect 27672 5120 30788 5148
rect 27672 5108 27678 5120
rect 32306 5108 32312 5160
rect 32364 5148 32370 5160
rect 34701 5151 34759 5157
rect 34701 5148 34713 5151
rect 32364 5120 34713 5148
rect 32364 5108 32370 5120
rect 34701 5117 34713 5120
rect 34747 5117 34759 5151
rect 34701 5111 34759 5117
rect 26786 5040 26792 5092
rect 26844 5080 26850 5092
rect 29273 5083 29331 5089
rect 29273 5080 29285 5083
rect 26844 5052 29285 5080
rect 26844 5040 26850 5052
rect 29273 5049 29285 5052
rect 29319 5049 29331 5083
rect 29273 5043 29331 5049
rect 29730 5040 29736 5092
rect 29788 5080 29794 5092
rect 31205 5083 31263 5089
rect 31205 5080 31217 5083
rect 29788 5052 31217 5080
rect 29788 5040 29794 5052
rect 31205 5049 31217 5052
rect 31251 5049 31263 5083
rect 32398 5080 32404 5092
rect 32359 5052 32404 5080
rect 31205 5043 31263 5049
rect 32398 5040 32404 5052
rect 32456 5040 32462 5092
rect 25372 4984 26464 5012
rect 26513 5015 26571 5021
rect 25372 4972 25378 4984
rect 26513 4981 26525 5015
rect 26559 5012 26571 5015
rect 27890 5012 27896 5024
rect 26559 4984 27896 5012
rect 26559 4981 26571 4984
rect 26513 4975 26571 4981
rect 27890 4972 27896 4984
rect 27948 4972 27954 5024
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28810 5012 28816 5024
rect 28500 4984 28816 5012
rect 28500 4972 28506 4984
rect 28810 4972 28816 4984
rect 28868 4972 28874 5024
rect 29178 4972 29184 5024
rect 29236 5012 29242 5024
rect 30282 5012 30288 5024
rect 29236 4984 30288 5012
rect 29236 4972 29242 4984
rect 30282 4972 30288 4984
rect 30340 4972 30346 5024
rect 31662 4972 31668 5024
rect 31720 5012 31726 5024
rect 33594 5012 33600 5024
rect 31720 4984 33600 5012
rect 31720 4972 31726 4984
rect 33594 4972 33600 4984
rect 33652 5012 33658 5024
rect 35805 5015 35863 5021
rect 35805 5012 35817 5015
rect 33652 4984 35817 5012
rect 33652 4972 33658 4984
rect 35805 4981 35817 4984
rect 35851 5012 35863 5015
rect 36357 5015 36415 5021
rect 36357 5012 36369 5015
rect 35851 4984 36369 5012
rect 35851 4981 35863 4984
rect 35805 4975 35863 4981
rect 36357 4981 36369 4984
rect 36403 5012 36415 5015
rect 36446 5012 36452 5024
rect 36403 4984 36452 5012
rect 36403 4981 36415 4984
rect 36357 4975 36415 4981
rect 36446 4972 36452 4984
rect 36504 4972 36510 5024
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10042 4808 10048 4820
rect 9723 4780 10048 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10042 4768 10048 4780
rect 10100 4808 10106 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 10100 4780 10149 4808
rect 10100 4768 10106 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 10137 4771 10195 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 13538 4808 13544 4820
rect 11664 4780 13400 4808
rect 13499 4780 13544 4808
rect 11664 4768 11670 4780
rect 6917 4743 6975 4749
rect 6917 4709 6929 4743
rect 6963 4740 6975 4743
rect 9582 4740 9588 4752
rect 6963 4712 9588 4740
rect 6963 4709 6975 4712
rect 6917 4703 6975 4709
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4740 11391 4743
rect 13262 4740 13268 4752
rect 11379 4712 13268 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13372 4740 13400 4780
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14642 4808 14648 4820
rect 14415 4780 14648 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15859 4811 15917 4817
rect 15859 4808 15871 4811
rect 14884 4780 15871 4808
rect 14884 4768 14890 4780
rect 15859 4777 15871 4780
rect 15905 4808 15917 4811
rect 18322 4808 18328 4820
rect 15905 4780 18328 4808
rect 15905 4777 15917 4780
rect 15859 4771 15917 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 28721 4811 28779 4817
rect 28721 4808 28733 4811
rect 18432 4780 28733 4808
rect 14550 4740 14556 4752
rect 13372 4712 14556 4740
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 14274 4672 14280 4684
rect 8996 4644 14280 4672
rect 8996 4632 9002 4644
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4672 16175 4675
rect 17034 4672 17040 4684
rect 16163 4644 17040 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 8110 4604 8116 4616
rect 6411 4576 8116 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 18432 4590 18460 4780
rect 28721 4777 28733 4780
rect 28767 4777 28779 4811
rect 28721 4771 28779 4777
rect 29454 4768 29460 4820
rect 29512 4808 29518 4820
rect 29825 4811 29883 4817
rect 29825 4808 29837 4811
rect 29512 4780 29837 4808
rect 29512 4768 29518 4780
rect 29825 4777 29837 4780
rect 29871 4777 29883 4811
rect 29825 4771 29883 4777
rect 30190 4768 30196 4820
rect 30248 4808 30254 4820
rect 31202 4808 31208 4820
rect 30248 4780 31208 4808
rect 30248 4768 30254 4780
rect 31202 4768 31208 4780
rect 31260 4808 31266 4820
rect 31662 4808 31668 4820
rect 31260 4780 31668 4808
rect 31260 4768 31266 4780
rect 31662 4768 31668 4780
rect 31720 4768 31726 4820
rect 31754 4768 31760 4820
rect 31812 4808 31818 4820
rect 31812 4780 31857 4808
rect 31812 4768 31818 4780
rect 18506 4700 18512 4752
rect 18564 4740 18570 4752
rect 18785 4743 18843 4749
rect 18785 4740 18797 4743
rect 18564 4712 18797 4740
rect 18564 4700 18570 4712
rect 18785 4709 18797 4712
rect 18831 4740 18843 4743
rect 19334 4740 19340 4752
rect 18831 4712 19340 4740
rect 18831 4709 18843 4712
rect 18785 4703 18843 4709
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 21174 4740 21180 4752
rect 21087 4712 21180 4740
rect 21174 4700 21180 4712
rect 21232 4740 21238 4752
rect 21450 4740 21456 4752
rect 21232 4712 21456 4740
rect 21232 4700 21238 4712
rect 21450 4700 21456 4712
rect 21508 4700 21514 4752
rect 24486 4700 24492 4752
rect 24544 4740 24550 4752
rect 27706 4740 27712 4752
rect 24544 4712 27712 4740
rect 24544 4700 24550 4712
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 28258 4700 28264 4752
rect 28316 4740 28322 4752
rect 30006 4740 30012 4752
rect 28316 4712 30012 4740
rect 28316 4700 28322 4712
rect 30006 4700 30012 4712
rect 30064 4700 30070 4752
rect 31478 4700 31484 4752
rect 31536 4740 31542 4752
rect 35437 4743 35495 4749
rect 35437 4740 35449 4743
rect 31536 4712 35449 4740
rect 31536 4700 31542 4712
rect 35437 4709 35449 4712
rect 35483 4709 35495 4743
rect 35437 4703 35495 4709
rect 19426 4672 19432 4684
rect 19387 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19794 4632 19800 4684
rect 19852 4672 19858 4684
rect 28077 4675 28135 4681
rect 28077 4672 28089 4675
rect 19852 4644 28089 4672
rect 19852 4632 19858 4644
rect 28077 4641 28089 4644
rect 28123 4641 28135 4675
rect 30190 4672 30196 4684
rect 28077 4635 28135 4641
rect 28828 4644 30196 4672
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 7469 4539 7527 4545
rect 7469 4505 7481 4539
rect 7515 4536 7527 4539
rect 13630 4536 13636 4548
rect 7515 4508 13636 4536
rect 7515 4505 7527 4508
rect 7469 4499 7527 4505
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 19705 4539 19763 4545
rect 13780 4508 14674 4536
rect 13780 4496 13786 4508
rect 19705 4505 19717 4539
rect 19751 4505 19763 4539
rect 22020 4536 22048 4567
rect 23566 4564 23572 4616
rect 23624 4604 23630 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 23624 4576 24685 4604
rect 23624 4564 23630 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 25774 4604 25780 4616
rect 25735 4576 25780 4604
rect 24673 4567 24731 4573
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4604 26019 4607
rect 26050 4604 26056 4616
rect 26007 4576 26056 4604
rect 26007 4573 26019 4576
rect 25961 4567 26019 4573
rect 26050 4564 26056 4576
rect 26108 4564 26114 4616
rect 26160 4576 26556 4604
rect 22186 4536 22192 4548
rect 20930 4508 21312 4536
rect 22020 4508 22192 4536
rect 19705 4499 19763 4505
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4468 8082 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8076 4440 8493 4468
rect 8076 4428 8082 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 11882 4468 11888 4480
rect 11795 4440 11888 4468
rect 8481 4431 8539 4437
rect 11882 4428 11888 4440
rect 11940 4468 11946 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 11940 4440 12449 4468
rect 11940 4428 11946 4440
rect 12437 4437 12449 4440
rect 12483 4468 12495 4471
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12483 4440 13001 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 12989 4437 13001 4440
rect 13035 4468 13047 4471
rect 14090 4468 14096 4480
rect 13035 4440 14096 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 19720 4468 19748 4499
rect 14608 4440 19748 4468
rect 21284 4468 21312 4508
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 22278 4496 22284 4548
rect 22336 4536 22342 4548
rect 22554 4536 22560 4548
rect 22336 4508 22560 4536
rect 22336 4496 22342 4508
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 26160 4536 26188 4576
rect 26418 4536 26424 4548
rect 23506 4508 26188 4536
rect 26379 4508 26424 4536
rect 26418 4496 26424 4508
rect 26476 4496 26482 4548
rect 26528 4536 26556 4576
rect 27890 4564 27896 4616
rect 27948 4604 27954 4616
rect 28828 4613 28856 4644
rect 30190 4632 30196 4644
rect 30248 4632 30254 4684
rect 33226 4672 33232 4684
rect 30484 4644 33232 4672
rect 30484 4616 30512 4644
rect 28169 4607 28227 4613
rect 28169 4604 28181 4607
rect 27948 4576 28181 4604
rect 27948 4564 27954 4576
rect 28169 4573 28181 4576
rect 28215 4604 28227 4607
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 28215 4576 28825 4604
rect 28215 4573 28227 4576
rect 28169 4567 28227 4573
rect 28813 4573 28825 4576
rect 28859 4573 28871 4607
rect 28813 4567 28871 4573
rect 28902 4564 28908 4616
rect 28960 4604 28966 4616
rect 29546 4604 29552 4616
rect 28960 4576 29552 4604
rect 28960 4564 28966 4576
rect 29546 4564 29552 4576
rect 29604 4564 29610 4616
rect 29917 4607 29975 4613
rect 29917 4573 29929 4607
rect 29963 4604 29975 4607
rect 30466 4604 30472 4616
rect 29963 4576 30472 4604
rect 29963 4573 29975 4576
rect 29917 4567 29975 4573
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 30561 4607 30619 4613
rect 30561 4573 30573 4607
rect 30607 4604 30619 4607
rect 30650 4604 30656 4616
rect 30607 4576 30656 4604
rect 30607 4573 30619 4576
rect 30561 4567 30619 4573
rect 30650 4564 30656 4576
rect 30708 4564 30714 4616
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4604 31263 4607
rect 31294 4604 31300 4616
rect 31251 4576 31300 4604
rect 31251 4573 31263 4576
rect 31205 4567 31263 4573
rect 31294 4564 31300 4576
rect 31352 4564 31358 4616
rect 31846 4604 31852 4616
rect 31807 4576 31852 4604
rect 31846 4564 31852 4576
rect 31904 4564 31910 4616
rect 32508 4613 32536 4644
rect 33226 4632 33232 4644
rect 33284 4632 33290 4684
rect 33686 4672 33692 4684
rect 33599 4644 33692 4672
rect 33686 4632 33692 4644
rect 33744 4672 33750 4684
rect 34330 4672 34336 4684
rect 33744 4644 34336 4672
rect 33744 4632 33750 4644
rect 34330 4632 34336 4644
rect 34388 4632 34394 4684
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4573 32551 4607
rect 32493 4567 32551 4573
rect 32953 4607 33011 4613
rect 32953 4573 32965 4607
rect 32999 4604 33011 4607
rect 32999 4576 35020 4604
rect 32999 4573 33011 4576
rect 32953 4567 33011 4573
rect 26786 4536 26792 4548
rect 26528 4508 26792 4536
rect 26786 4496 26792 4508
rect 26844 4496 26850 4548
rect 27338 4536 27344 4548
rect 27299 4508 27344 4536
rect 27338 4496 27344 4508
rect 27396 4496 27402 4548
rect 27433 4539 27491 4545
rect 27433 4505 27445 4539
rect 27479 4505 27491 4539
rect 27433 4499 27491 4505
rect 23658 4468 23664 4480
rect 21284 4440 23664 4468
rect 14608 4428 14614 4440
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 23750 4428 23756 4480
rect 23808 4468 23814 4480
rect 24302 4468 24308 4480
rect 23808 4440 24308 4468
rect 23808 4428 23814 4440
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 24486 4428 24492 4480
rect 24544 4468 24550 4480
rect 24765 4471 24823 4477
rect 24765 4468 24777 4471
rect 24544 4440 24777 4468
rect 24544 4428 24550 4440
rect 24765 4437 24777 4440
rect 24811 4437 24823 4471
rect 24765 4431 24823 4437
rect 25038 4428 25044 4480
rect 25096 4468 25102 4480
rect 25317 4471 25375 4477
rect 25317 4468 25329 4471
rect 25096 4440 25329 4468
rect 25096 4428 25102 4440
rect 25317 4437 25329 4440
rect 25363 4468 25375 4471
rect 27448 4468 27476 4499
rect 27706 4496 27712 4548
rect 27764 4536 27770 4548
rect 31113 4539 31171 4545
rect 31113 4536 31125 4539
rect 27764 4508 29776 4536
rect 27764 4496 27770 4508
rect 25363 4440 27476 4468
rect 25363 4437 25375 4440
rect 25317 4431 25375 4437
rect 27614 4428 27620 4480
rect 27672 4468 27678 4480
rect 29638 4468 29644 4480
rect 27672 4440 29644 4468
rect 27672 4428 27678 4440
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 29748 4468 29776 4508
rect 29932 4508 31125 4536
rect 29932 4468 29960 4508
rect 31113 4505 31125 4508
rect 31159 4505 31171 4539
rect 31113 4499 31171 4505
rect 31478 4496 31484 4548
rect 31536 4536 31542 4548
rect 32398 4536 32404 4548
rect 31536 4508 31892 4536
rect 32359 4508 32404 4536
rect 31536 4496 31542 4508
rect 29748 4440 29960 4468
rect 30006 4428 30012 4480
rect 30064 4468 30070 4480
rect 30377 4471 30435 4477
rect 30377 4468 30389 4471
rect 30064 4440 30389 4468
rect 30064 4428 30070 4440
rect 30377 4437 30389 4440
rect 30423 4437 30435 4471
rect 31864 4468 31892 4508
rect 32398 4496 32404 4508
rect 32456 4496 32462 4548
rect 32968 4468 32996 4567
rect 34790 4536 34796 4548
rect 33152 4508 34796 4536
rect 33152 4477 33180 4508
rect 34790 4496 34796 4508
rect 34848 4496 34854 4548
rect 34992 4545 35020 4576
rect 38010 4564 38016 4616
rect 38068 4604 38074 4616
rect 38289 4607 38347 4613
rect 38289 4604 38301 4607
rect 38068 4576 38301 4604
rect 38068 4564 38074 4576
rect 38289 4573 38301 4576
rect 38335 4573 38347 4607
rect 38289 4567 38347 4573
rect 34977 4539 35035 4545
rect 34977 4505 34989 4539
rect 35023 4536 35035 4539
rect 35989 4539 36047 4545
rect 35989 4536 36001 4539
rect 35023 4508 36001 4536
rect 35023 4505 35035 4508
rect 34977 4499 35035 4505
rect 35989 4505 36001 4508
rect 36035 4505 36047 4539
rect 35989 4499 36047 4505
rect 36446 4496 36452 4548
rect 36504 4536 36510 4548
rect 37093 4539 37151 4545
rect 37093 4536 37105 4539
rect 36504 4508 37105 4536
rect 36504 4496 36510 4508
rect 37093 4505 37105 4508
rect 37139 4505 37151 4539
rect 37093 4499 37151 4505
rect 31864 4440 32996 4468
rect 33137 4471 33195 4477
rect 30377 4431 30435 4437
rect 33137 4437 33149 4471
rect 33183 4437 33195 4471
rect 33137 4431 33195 4437
rect 33594 4428 33600 4480
rect 33652 4468 33658 4480
rect 34149 4471 34207 4477
rect 34149 4468 34161 4471
rect 33652 4440 34161 4468
rect 33652 4428 33658 4440
rect 34149 4437 34161 4440
rect 34195 4437 34207 4471
rect 34149 4431 34207 4437
rect 35710 4428 35716 4480
rect 35768 4468 35774 4480
rect 36541 4471 36599 4477
rect 36541 4468 36553 4471
rect 35768 4440 36553 4468
rect 35768 4428 35774 4440
rect 36541 4437 36553 4440
rect 36587 4437 36599 4471
rect 38102 4468 38108 4480
rect 38063 4440 38108 4468
rect 36541 4431 36599 4437
rect 38102 4428 38108 4440
rect 38160 4428 38166 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 10042 4264 10048 4276
rect 9955 4236 10048 4264
rect 10042 4224 10048 4236
rect 10100 4264 10106 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10100 4236 10609 4264
rect 10100 4224 10106 4236
rect 10597 4233 10609 4236
rect 10643 4264 10655 4267
rect 11882 4264 11888 4276
rect 10643 4236 11888 4264
rect 10643 4233 10655 4236
rect 10597 4227 10655 4233
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12345 4267 12403 4273
rect 12345 4264 12357 4267
rect 12032 4236 12357 4264
rect 12032 4224 12038 4236
rect 12345 4233 12357 4236
rect 12391 4233 12403 4267
rect 12345 4227 12403 4233
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 19242 4264 19248 4276
rect 14424 4236 19248 4264
rect 14424 4224 14430 4236
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 22278 4264 22284 4276
rect 21284 4236 22284 4264
rect 13354 4156 13360 4208
rect 13412 4156 13418 4208
rect 14734 4156 14740 4208
rect 14792 4196 14798 4208
rect 21174 4196 21180 4208
rect 14792 4168 14858 4196
rect 16316 4168 17080 4196
rect 14792 4156 14798 4168
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 12526 4128 12532 4140
rect 7331 4100 12532 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 16316 4137 16344 4168
rect 17052 4140 17080 4168
rect 19168 4168 21180 4196
rect 16301 4131 16359 4137
rect 14148 4100 14193 4128
rect 14148 4088 14154 4100
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6043 4032 9444 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 7745 3995 7803 4001
rect 7745 3992 7757 3995
rect 6932 3964 7757 3992
rect 6932 3936 6960 3964
rect 7745 3961 7757 3964
rect 7791 3992 7803 3995
rect 8018 3992 8024 4004
rect 7791 3964 8024 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 8018 3952 8024 3964
rect 8076 3992 8082 4004
rect 8297 3995 8355 4001
rect 8297 3992 8309 3995
rect 8076 3964 8309 3992
rect 8076 3952 8082 3964
rect 8297 3961 8309 3964
rect 8343 3992 8355 3995
rect 8849 3995 8907 4001
rect 8849 3992 8861 3995
rect 8343 3964 8861 3992
rect 8343 3961 8355 3964
rect 8297 3955 8355 3961
rect 8849 3961 8861 3964
rect 8895 3961 8907 3995
rect 8849 3955 8907 3961
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4120 3896 4445 3924
rect 4120 3884 4126 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6914 3924 6920 3936
rect 6779 3896 6920 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 8662 3924 8668 3936
rect 7064 3896 8668 3924
rect 7064 3884 7070 3896
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9416 3924 9444 4032
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 13817 4063 13875 4069
rect 10376 4032 12848 4060
rect 10376 4020 10382 4032
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3992 9551 3995
rect 12710 3992 12716 4004
rect 9539 3964 12716 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 11054 3924 11060 3936
rect 9416 3896 11060 3924
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11238 3924 11244 3936
rect 11195 3896 11244 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12820 3924 12848 4032
rect 13817 4029 13829 4063
rect 13863 4060 13875 4063
rect 14182 4060 14188 4072
rect 13863 4032 14188 4060
rect 13863 4029 13875 4032
rect 13817 4023 13875 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16868 3992 16896 4091
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 17092 4100 17601 4128
rect 17092 4088 17098 4100
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 17862 4060 17868 4072
rect 17823 4032 17868 4060
rect 17862 4020 17868 4032
rect 17920 4060 17926 4072
rect 19168 4060 19196 4168
rect 21174 4156 21180 4168
rect 21232 4156 21238 4208
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19300 4100 19901 4128
rect 19300 4088 19306 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20772 4100 20817 4128
rect 20772 4088 20778 4100
rect 17920 4032 19196 4060
rect 19337 4063 19395 4069
rect 17920 4020 17926 4032
rect 19337 4029 19349 4063
rect 19383 4060 19395 4063
rect 21284 4060 21312 4236
rect 22278 4224 22284 4236
rect 22336 4224 22342 4276
rect 23753 4267 23811 4273
rect 23753 4233 23765 4267
rect 23799 4264 23811 4267
rect 24854 4264 24860 4276
rect 23799 4236 24860 4264
rect 23799 4233 23811 4236
rect 23753 4227 23811 4233
rect 24854 4224 24860 4236
rect 24912 4224 24918 4276
rect 25498 4224 25504 4276
rect 25556 4264 25562 4276
rect 25961 4267 26019 4273
rect 25961 4264 25973 4267
rect 25556 4236 25973 4264
rect 25556 4224 25562 4236
rect 25961 4233 25973 4236
rect 26007 4264 26019 4267
rect 29822 4264 29828 4276
rect 26007 4236 29828 4264
rect 26007 4233 26019 4236
rect 25961 4227 26019 4233
rect 29822 4224 29828 4236
rect 29880 4224 29886 4276
rect 34793 4267 34851 4273
rect 34793 4264 34805 4267
rect 30208 4236 34805 4264
rect 21453 4199 21511 4205
rect 21453 4165 21465 4199
rect 21499 4196 21511 4199
rect 22186 4196 22192 4208
rect 21499 4168 22192 4196
rect 21499 4165 21511 4168
rect 21453 4159 21511 4165
rect 22020 4137 22048 4168
rect 22186 4156 22192 4168
rect 22244 4156 22250 4208
rect 24118 4196 24124 4208
rect 23506 4168 24124 4196
rect 24118 4156 24124 4168
rect 24176 4156 24182 4208
rect 24578 4196 24584 4208
rect 24228 4168 24584 4196
rect 24228 4137 24256 4168
rect 24578 4156 24584 4168
rect 24636 4156 24642 4208
rect 27430 4196 27436 4208
rect 25714 4168 27436 4196
rect 27430 4156 27436 4168
rect 27488 4156 27494 4208
rect 27709 4199 27767 4205
rect 27709 4165 27721 4199
rect 27755 4196 27767 4199
rect 30101 4199 30159 4205
rect 30101 4196 30113 4199
rect 27755 4168 30113 4196
rect 27755 4165 27767 4168
rect 27709 4159 27767 4165
rect 30101 4165 30113 4168
rect 30147 4165 30159 4199
rect 30101 4159 30159 4165
rect 30208 4140 30236 4236
rect 34793 4233 34805 4236
rect 34839 4233 34851 4267
rect 36446 4264 36452 4276
rect 36407 4236 36452 4264
rect 34793 4227 34851 4233
rect 36446 4224 36452 4236
rect 36504 4224 36510 4276
rect 33318 4196 33324 4208
rect 32508 4168 33324 4196
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4097 24271 4131
rect 26234 4128 26240 4140
rect 24213 4091 24271 4097
rect 25700 4100 26240 4128
rect 19383 4032 21312 4060
rect 19383 4029 19395 4032
rect 19337 4023 19395 4029
rect 21358 4020 21364 4072
rect 21416 4060 21422 4072
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 21416 4032 22293 4060
rect 21416 4020 21422 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 22428 4032 23336 4060
rect 22428 4020 22434 4032
rect 14016 3964 14688 3992
rect 14016 3924 14044 3964
rect 12820 3896 14044 3924
rect 14660 3924 14688 3964
rect 16224 3964 16896 3992
rect 16224 3924 16252 3964
rect 19150 3952 19156 4004
rect 19208 3992 19214 4004
rect 20625 3995 20683 4001
rect 20625 3992 20637 3995
rect 19208 3964 20637 3992
rect 19208 3952 19214 3964
rect 20625 3961 20637 3964
rect 20671 3961 20683 3995
rect 20625 3955 20683 3961
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 22002 3992 22008 4004
rect 20772 3964 22008 3992
rect 20772 3952 20778 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 14660 3896 16252 3924
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 16816 3896 17049 3924
rect 16816 3884 16822 3896
rect 17037 3893 17049 3896
rect 17083 3893 17095 3927
rect 19978 3924 19984 3936
rect 19939 3896 19984 3924
rect 17037 3887 17095 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 21726 3884 21732 3936
rect 21784 3924 21790 3936
rect 23014 3924 23020 3936
rect 21784 3896 23020 3924
rect 21784 3884 21790 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23308 3924 23336 4032
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24176 4032 24501 4060
rect 24176 4020 24182 4032
rect 24489 4029 24501 4032
rect 24535 4060 24547 4063
rect 25700 4060 25728 4100
rect 26234 4088 26240 4100
rect 26292 4088 26298 4140
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 26694 4128 26700 4140
rect 26467 4100 26700 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 26694 4088 26700 4100
rect 26752 4088 26758 4140
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 28905 4131 28963 4137
rect 28905 4128 28917 4131
rect 28868 4100 28917 4128
rect 28868 4088 28874 4100
rect 28905 4097 28917 4100
rect 28951 4097 28963 4131
rect 28905 4091 28963 4097
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 29549 4131 29607 4137
rect 29052 4100 29132 4128
rect 29052 4088 29058 4100
rect 24535 4032 25728 4060
rect 24535 4029 24547 4032
rect 24489 4023 24547 4029
rect 26142 4020 26148 4072
rect 26200 4060 26206 4072
rect 27522 4060 27528 4072
rect 26200 4032 27384 4060
rect 27483 4032 27528 4060
rect 26200 4020 26206 4032
rect 26418 3992 26424 4004
rect 25516 3964 26424 3992
rect 25516 3924 25544 3964
rect 26418 3952 26424 3964
rect 26476 3952 26482 4004
rect 26602 3952 26608 4004
rect 26660 3992 26666 4004
rect 27356 3992 27384 4032
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 27798 4060 27804 4072
rect 27759 4032 27804 4060
rect 27798 4020 27804 4032
rect 27856 4020 27862 4072
rect 28534 4020 28540 4072
rect 28592 4060 28598 4072
rect 28592 4032 28994 4060
rect 28592 4020 28598 4032
rect 28813 3995 28871 4001
rect 28813 3992 28825 3995
rect 26660 3964 27108 3992
rect 27356 3964 28825 3992
rect 26660 3952 26666 3964
rect 23308 3896 25544 3924
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26142 3924 26148 3936
rect 26016 3896 26148 3924
rect 26016 3884 26022 3896
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 26513 3927 26571 3933
rect 26513 3893 26525 3927
rect 26559 3924 26571 3927
rect 26970 3924 26976 3936
rect 26559 3896 26976 3924
rect 26559 3893 26571 3896
rect 26513 3887 26571 3893
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 27080 3924 27108 3964
rect 28813 3961 28825 3964
rect 28859 3961 28871 3995
rect 28813 3955 28871 3961
rect 28074 3924 28080 3936
rect 27080 3896 28080 3924
rect 28074 3884 28080 3896
rect 28132 3884 28138 3936
rect 28966 3924 28994 4032
rect 29104 3992 29132 4100
rect 29549 4097 29561 4131
rect 29595 4128 29607 4131
rect 30190 4128 30196 4140
rect 29595 4100 29684 4128
rect 30103 4100 30196 4128
rect 29595 4097 29607 4100
rect 29549 4091 29607 4097
rect 29270 4020 29276 4072
rect 29328 4060 29334 4072
rect 29457 4063 29515 4069
rect 29457 4060 29469 4063
rect 29328 4032 29469 4060
rect 29328 4020 29334 4032
rect 29457 4029 29469 4032
rect 29503 4029 29515 4063
rect 29656 4060 29684 4100
rect 30190 4088 30196 4100
rect 30248 4088 30254 4140
rect 30282 4088 30288 4140
rect 30340 4128 30346 4140
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30340 4100 30849 4128
rect 30340 4088 30346 4100
rect 30837 4097 30849 4100
rect 30883 4128 30895 4131
rect 31478 4128 31484 4140
rect 30883 4100 31340 4128
rect 31439 4100 31484 4128
rect 30883 4097 30895 4100
rect 30837 4091 30895 4097
rect 30098 4060 30104 4072
rect 29656 4032 30104 4060
rect 29457 4023 29515 4029
rect 30098 4020 30104 4032
rect 30156 4020 30162 4072
rect 31312 4060 31340 4100
rect 31478 4088 31484 4100
rect 31536 4088 31542 4140
rect 32122 4088 32128 4140
rect 32180 4128 32186 4140
rect 32508 4137 32536 4168
rect 33318 4156 33324 4168
rect 33376 4196 33382 4208
rect 38197 4199 38255 4205
rect 33376 4168 33824 4196
rect 33376 4156 33382 4168
rect 32493 4131 32551 4137
rect 32493 4128 32505 4131
rect 32180 4100 32505 4128
rect 32180 4088 32186 4100
rect 32493 4097 32505 4100
rect 32539 4097 32551 4131
rect 32493 4091 32551 4097
rect 32582 4088 32588 4140
rect 32640 4128 32646 4140
rect 33796 4137 33824 4168
rect 38197 4165 38209 4199
rect 38243 4196 38255 4199
rect 38286 4196 38292 4208
rect 38243 4168 38292 4196
rect 38243 4165 38255 4168
rect 38197 4159 38255 4165
rect 38286 4156 38292 4168
rect 38344 4156 38350 4208
rect 33137 4131 33195 4137
rect 33137 4128 33149 4131
rect 32640 4100 33149 4128
rect 32640 4088 32646 4100
rect 33137 4097 33149 4100
rect 33183 4097 33195 4131
rect 33137 4091 33195 4097
rect 33781 4131 33839 4137
rect 33781 4097 33793 4131
rect 33827 4128 33839 4131
rect 35345 4131 35403 4137
rect 35345 4128 35357 4131
rect 33827 4100 35357 4128
rect 33827 4097 33839 4100
rect 33781 4091 33839 4097
rect 35345 4097 35357 4100
rect 35391 4128 35403 4131
rect 35710 4128 35716 4140
rect 35391 4100 35716 4128
rect 35391 4097 35403 4100
rect 35345 4091 35403 4097
rect 33152 4060 33180 4091
rect 35710 4088 35716 4100
rect 35768 4128 35774 4140
rect 35897 4131 35955 4137
rect 35897 4128 35909 4131
rect 35768 4100 35909 4128
rect 35768 4088 35774 4100
rect 35897 4097 35909 4100
rect 35943 4097 35955 4131
rect 35897 4091 35955 4097
rect 37918 4088 37924 4140
rect 37976 4128 37982 4140
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 37976 4100 38025 4128
rect 37976 4088 37982 4100
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 38013 4091 38071 4097
rect 36262 4060 36268 4072
rect 31312 4032 31524 4060
rect 33152 4032 36268 4060
rect 31389 3995 31447 4001
rect 31389 3992 31401 3995
rect 29104 3964 31401 3992
rect 31389 3961 31401 3964
rect 31435 3961 31447 3995
rect 31389 3955 31447 3961
rect 30190 3924 30196 3936
rect 28966 3896 30196 3924
rect 30190 3884 30196 3896
rect 30248 3884 30254 3936
rect 30742 3924 30748 3936
rect 30703 3896 30748 3924
rect 30742 3884 30748 3896
rect 30800 3884 30806 3936
rect 31496 3924 31524 4032
rect 36262 4020 36268 4032
rect 36320 4020 36326 4072
rect 31570 3952 31576 4004
rect 31628 3992 31634 4004
rect 34241 3995 34299 4001
rect 34241 3992 34253 3995
rect 31628 3964 34253 3992
rect 31628 3952 31634 3964
rect 34241 3961 34253 3964
rect 34287 3961 34299 3995
rect 37461 3995 37519 4001
rect 37461 3992 37473 3995
rect 34241 3955 34299 3961
rect 34348 3964 37473 3992
rect 32122 3924 32128 3936
rect 31496 3896 32128 3924
rect 32122 3884 32128 3896
rect 32180 3884 32186 3936
rect 32398 3924 32404 3936
rect 32359 3896 32404 3924
rect 32398 3884 32404 3896
rect 32456 3884 32462 3936
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 33045 3927 33103 3933
rect 33045 3924 33057 3927
rect 32732 3896 33057 3924
rect 32732 3884 32738 3896
rect 33045 3893 33057 3896
rect 33091 3893 33103 3927
rect 33686 3924 33692 3936
rect 33647 3896 33692 3924
rect 33045 3887 33103 3893
rect 33686 3884 33692 3896
rect 33744 3884 33750 3936
rect 33778 3884 33784 3936
rect 33836 3924 33842 3936
rect 34348 3924 34376 3964
rect 37461 3961 37473 3964
rect 37507 3961 37519 3995
rect 37461 3955 37519 3961
rect 33836 3896 34376 3924
rect 33836 3884 33842 3896
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 9677 3723 9735 3729
rect 5583 3692 9628 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 7653 3655 7711 3661
rect 7653 3652 7665 3655
rect 5500 3624 7665 3652
rect 5500 3612 5506 3624
rect 7653 3621 7665 3624
rect 7699 3621 7711 3655
rect 9600 3652 9628 3692
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9766 3720 9772 3732
rect 9723 3692 9772 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9766 3680 9772 3692
rect 9824 3720 9830 3732
rect 10042 3720 10048 3732
rect 9824 3692 10048 3720
rect 9824 3680 9830 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 12434 3720 12440 3732
rect 10376 3692 10421 3720
rect 11256 3692 12440 3720
rect 10376 3680 10382 3692
rect 11256 3652 11284 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12676 3692 16988 3720
rect 12676 3680 12682 3692
rect 7653 3615 7711 3621
rect 7760 3624 9536 3652
rect 9600 3624 11284 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 4249 3587 4307 3593
rect 1903 3556 2774 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2746 3448 2774 3556
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 7760 3584 7788 3624
rect 8110 3584 8116 3596
rect 4295 3556 7788 3584
rect 7860 3556 8116 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 7860 3525 7888 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 9508 3584 9536 3624
rect 10962 3584 10968 3596
rect 9508 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4120 3488 4169 3516
rect 4120 3476 4126 3488
rect 4157 3485 4169 3488
rect 4203 3516 4215 3519
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4203 3488 4905 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8260 3488 8309 3516
rect 8260 3476 8266 3488
rect 8297 3485 8309 3488
rect 8343 3516 8355 3519
rect 10042 3516 10048 3528
rect 8343 3488 10048 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 11256 3525 11284 3624
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13320 3624 13584 3652
rect 13320 3612 13326 3624
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11882 3584 11888 3596
rect 11388 3556 11888 3584
rect 11388 3544 11394 3556
rect 11882 3544 11888 3556
rect 11940 3584 11946 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11940 3556 11989 3584
rect 11940 3544 11946 3556
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 13556 3584 13584 3624
rect 13630 3612 13636 3664
rect 13688 3652 13694 3664
rect 14274 3652 14280 3664
rect 13688 3624 14280 3652
rect 13688 3612 13694 3624
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 13722 3584 13728 3596
rect 12768 3556 13492 3584
rect 13556 3556 13728 3584
rect 12768 3544 12774 3556
rect 11241 3519 11299 3525
rect 10192 3488 10237 3516
rect 10192 3476 10198 3488
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 13464 3516 13492 3556
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 16114 3584 16120 3596
rect 13832 3556 16120 3584
rect 13832 3516 13860 3556
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16776 3556 16865 3584
rect 13464 3488 13860 3516
rect 11241 3479 11299 3485
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14148 3488 14381 3516
rect 14148 3476 14154 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 14369 3479 14427 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 7193 3451 7251 3457
rect 2746 3420 7144 3448
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3329 3383 3387 3389
rect 3329 3380 3341 3383
rect 3292 3352 3341 3380
rect 3292 3340 3298 3352
rect 3329 3349 3341 3352
rect 3375 3349 3387 3383
rect 5994 3380 6000 3392
rect 5955 3352 6000 3380
rect 3329 3343 3387 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 7006 3380 7012 3392
rect 6687 3352 7012 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7116 3380 7144 3420
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 7239 3420 11284 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 8386 3380 8392 3392
rect 7116 3352 8392 3380
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8938 3380 8944 3392
rect 8527 3352 8944 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 11146 3380 11152 3392
rect 11107 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11256 3380 11284 3420
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 12250 3448 12256 3460
rect 11572 3420 12256 3448
rect 11572 3408 11578 3420
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12584 3420 12742 3448
rect 12584 3408 12590 3420
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 14645 3451 14703 3457
rect 14645 3448 14657 3451
rect 13596 3420 14657 3448
rect 13596 3408 13602 3420
rect 14645 3417 14657 3420
rect 14691 3417 14703 3451
rect 16206 3448 16212 3460
rect 15870 3420 16212 3448
rect 14645 3411 14703 3417
rect 15948 3380 15976 3420
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 11256 3352 15976 3380
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 16776 3380 16804 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 16960 3584 16988 3692
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 21726 3720 21732 3732
rect 17276 3692 21732 3720
rect 17276 3680 17282 3692
rect 21726 3680 21732 3692
rect 21784 3680 21790 3732
rect 21818 3680 21824 3732
rect 21876 3720 21882 3732
rect 21876 3692 26740 3720
rect 21876 3680 21882 3692
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 19613 3655 19671 3661
rect 19613 3652 19625 3655
rect 18196 3624 19625 3652
rect 18196 3612 18202 3624
rect 19613 3621 19625 3624
rect 19659 3621 19671 3655
rect 19613 3615 19671 3621
rect 23308 3624 24716 3652
rect 16960 3556 19472 3584
rect 16853 3547 16911 3553
rect 19444 3525 19472 3556
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22244 3556 22600 3584
rect 22244 3544 22250 3556
rect 22572 3525 22600 3556
rect 23308 3525 23336 3624
rect 24688 3584 24716 3624
rect 24946 3584 24952 3596
rect 23400 3556 24624 3584
rect 24688 3556 24952 3584
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 17129 3451 17187 3457
rect 17129 3448 17141 3451
rect 16908 3420 17141 3448
rect 16908 3408 16914 3420
rect 17129 3417 17141 3420
rect 17175 3417 17187 3451
rect 19978 3448 19984 3460
rect 18354 3420 19984 3448
rect 17129 3411 17187 3417
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 20070 3408 20076 3460
rect 20128 3448 20134 3460
rect 20530 3448 20536 3460
rect 20128 3420 20536 3448
rect 20128 3408 20134 3420
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 21818 3408 21824 3460
rect 21876 3408 21882 3460
rect 22281 3451 22339 3457
rect 22281 3417 22293 3451
rect 22327 3448 22339 3451
rect 22370 3448 22376 3460
rect 22327 3420 22376 3448
rect 22327 3417 22339 3420
rect 22281 3411 22339 3417
rect 22370 3408 22376 3420
rect 22428 3408 22434 3460
rect 22572 3448 22600 3479
rect 23400 3448 23428 3556
rect 24596 3528 24624 3556
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 25222 3544 25228 3596
rect 25280 3584 25286 3596
rect 26602 3584 26608 3596
rect 25280 3556 26608 3584
rect 25280 3544 25286 3556
rect 26602 3544 26608 3556
rect 26660 3544 26666 3596
rect 26712 3584 26740 3692
rect 27338 3680 27344 3732
rect 27396 3720 27402 3732
rect 29825 3723 29883 3729
rect 29825 3720 29837 3723
rect 27396 3692 29837 3720
rect 27396 3680 27402 3692
rect 29825 3689 29837 3692
rect 29871 3689 29883 3723
rect 29825 3683 29883 3689
rect 32582 3680 32588 3732
rect 32640 3720 32646 3732
rect 33778 3720 33784 3732
rect 32640 3692 33784 3720
rect 32640 3680 32646 3692
rect 33778 3680 33784 3692
rect 33836 3680 33842 3732
rect 34330 3720 34336 3732
rect 34243 3692 34336 3720
rect 34330 3680 34336 3692
rect 34388 3720 34394 3732
rect 34885 3723 34943 3729
rect 34885 3720 34897 3723
rect 34388 3692 34897 3720
rect 34388 3680 34394 3692
rect 34885 3689 34897 3692
rect 34931 3689 34943 3723
rect 34885 3683 34943 3689
rect 35710 3680 35716 3732
rect 35768 3720 35774 3732
rect 35989 3723 36047 3729
rect 35989 3720 36001 3723
rect 35768 3692 36001 3720
rect 35768 3680 35774 3692
rect 35989 3689 36001 3692
rect 36035 3689 36047 3723
rect 35989 3683 36047 3689
rect 27430 3612 27436 3664
rect 27488 3652 27494 3664
rect 30926 3652 30932 3664
rect 27488 3624 30932 3652
rect 27488 3612 27494 3624
rect 30926 3612 30932 3624
rect 30984 3612 30990 3664
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 33870 3652 33876 3664
rect 31904 3624 33876 3652
rect 31904 3612 31910 3624
rect 31757 3587 31815 3593
rect 31757 3584 31769 3587
rect 26712 3556 31769 3584
rect 31757 3553 31769 3556
rect 31803 3553 31815 3587
rect 31757 3547 31815 3553
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3485 24087 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24029 3479 24087 3485
rect 22572 3420 23428 3448
rect 17034 3380 17040 3392
rect 16632 3352 17040 3380
rect 16632 3340 16638 3352
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 18414 3340 18420 3392
rect 18472 3380 18478 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18472 3352 18613 3380
rect 18472 3340 18478 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20714 3380 20720 3392
rect 19484 3352 20720 3380
rect 19484 3340 19490 3352
rect 20714 3340 20720 3352
rect 20772 3340 20778 3392
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 23109 3383 23167 3389
rect 23109 3380 23121 3383
rect 21324 3352 23121 3380
rect 21324 3340 21330 3352
rect 23109 3349 23121 3352
rect 23155 3349 23167 3383
rect 23109 3343 23167 3349
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 23845 3383 23903 3389
rect 23845 3380 23857 3383
rect 23256 3352 23857 3380
rect 23256 3340 23262 3352
rect 23845 3349 23857 3352
rect 23891 3349 23903 3383
rect 24044 3380 24072 3479
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27580 3488 27625 3516
rect 27580 3476 27586 3488
rect 27982 3476 27988 3528
rect 28040 3516 28046 3528
rect 28166 3516 28172 3528
rect 28040 3488 28172 3516
rect 28040 3476 28046 3488
rect 28166 3476 28172 3488
rect 28224 3476 28230 3528
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28408 3488 28733 3516
rect 28408 3476 28414 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3516 28871 3519
rect 28902 3516 28908 3528
rect 28859 3488 28908 3516
rect 28859 3485 28871 3488
rect 28813 3479 28871 3485
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 29733 3519 29791 3525
rect 29733 3485 29745 3519
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 24857 3451 24915 3457
rect 24857 3448 24869 3451
rect 24268 3420 24869 3448
rect 24268 3408 24274 3420
rect 24857 3417 24869 3420
rect 24903 3448 24915 3451
rect 25130 3448 25136 3460
rect 24903 3420 25136 3448
rect 24903 3417 24915 3420
rect 24857 3411 24915 3417
rect 25130 3408 25136 3420
rect 25188 3408 25194 3460
rect 26510 3448 26516 3460
rect 26344 3420 26516 3448
rect 25682 3380 25688 3392
rect 24044 3352 25688 3380
rect 23845 3343 23903 3349
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 26344 3389 26372 3420
rect 26510 3408 26516 3420
rect 26568 3408 26574 3460
rect 26881 3451 26939 3457
rect 26881 3417 26893 3451
rect 26927 3417 26939 3451
rect 26881 3411 26939 3417
rect 26329 3383 26387 3389
rect 26329 3349 26341 3383
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26418 3340 26424 3392
rect 26476 3380 26482 3392
rect 26896 3380 26924 3411
rect 26970 3408 26976 3460
rect 27028 3448 27034 3460
rect 27028 3420 27073 3448
rect 27028 3408 27034 3420
rect 27706 3408 27712 3460
rect 27764 3448 27770 3460
rect 29748 3448 29776 3479
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30561 3519 30619 3525
rect 30561 3516 30573 3519
rect 30340 3488 30573 3516
rect 30340 3476 30346 3488
rect 30561 3485 30573 3488
rect 30607 3516 30619 3519
rect 31018 3516 31024 3528
rect 30607 3488 31024 3516
rect 30607 3485 30619 3488
rect 30561 3479 30619 3485
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 31202 3516 31208 3528
rect 31163 3488 31208 3516
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 31846 3516 31852 3528
rect 31807 3488 31852 3516
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32508 3525 32536 3624
rect 33870 3612 33876 3624
rect 33928 3612 33934 3664
rect 34790 3612 34796 3664
rect 34848 3652 34854 3664
rect 34848 3624 38056 3652
rect 34848 3612 34854 3624
rect 33318 3544 33324 3596
rect 33376 3584 33382 3596
rect 35437 3587 35495 3593
rect 35437 3584 35449 3587
rect 33376 3556 35449 3584
rect 33376 3544 33382 3556
rect 35437 3553 35449 3556
rect 35483 3553 35495 3587
rect 35437 3547 35495 3553
rect 32493 3519 32551 3525
rect 32493 3485 32505 3519
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 32858 3476 32864 3528
rect 32916 3516 32922 3528
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 32916 3488 33149 3516
rect 32916 3476 32922 3488
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 31113 3451 31171 3457
rect 31113 3448 31125 3451
rect 27764 3420 29776 3448
rect 29840 3420 31125 3448
rect 27764 3408 27770 3420
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 26476 3352 28089 3380
rect 26476 3340 26482 3352
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 28077 3343 28135 3349
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 29840 3380 29868 3420
rect 31113 3417 31125 3420
rect 31159 3417 31171 3451
rect 31113 3411 31171 3417
rect 31662 3408 31668 3460
rect 31720 3448 31726 3460
rect 33045 3451 33103 3457
rect 33045 3448 33057 3451
rect 31720 3420 33057 3448
rect 31720 3408 31726 3420
rect 33045 3417 33057 3420
rect 33091 3417 33103 3451
rect 33152 3448 33180 3479
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 33781 3519 33839 3525
rect 33781 3516 33793 3519
rect 33284 3488 33793 3516
rect 33284 3476 33290 3488
rect 33781 3485 33793 3488
rect 33827 3516 33839 3519
rect 34422 3516 34428 3528
rect 33827 3488 34428 3516
rect 33827 3485 33839 3488
rect 33781 3479 33839 3485
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 36446 3476 36452 3528
rect 36504 3516 36510 3528
rect 38028 3525 38056 3624
rect 37277 3519 37335 3525
rect 37277 3516 37289 3519
rect 36504 3488 37289 3516
rect 36504 3476 36510 3488
rect 37277 3485 37289 3488
rect 37323 3485 37335 3519
rect 37277 3479 37335 3485
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 37001 3451 37059 3457
rect 37001 3448 37013 3451
rect 33152 3420 37013 3448
rect 33045 3411 33103 3417
rect 37001 3417 37013 3420
rect 37047 3417 37059 3451
rect 37001 3411 37059 3417
rect 30466 3380 30472 3392
rect 29420 3352 29868 3380
rect 30427 3352 30472 3380
rect 29420 3340 29426 3352
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 31754 3340 31760 3392
rect 31812 3380 31818 3392
rect 32401 3383 32459 3389
rect 32401 3380 32413 3383
rect 31812 3352 32413 3380
rect 31812 3340 31818 3352
rect 32401 3349 32413 3352
rect 32447 3349 32459 3383
rect 32401 3343 32459 3349
rect 33226 3340 33232 3392
rect 33284 3380 33290 3392
rect 33689 3383 33747 3389
rect 33689 3380 33701 3383
rect 33284 3352 33701 3380
rect 33284 3340 33290 3352
rect 33689 3349 33701 3352
rect 33735 3349 33747 3383
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 33689 3343 33747 3349
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2406 3176 2412 3188
rect 2319 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3176 2470 3188
rect 3418 3176 3424 3188
rect 2464 3148 3424 3176
rect 2464 3136 2470 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 9766 3176 9772 3188
rect 8076 3148 8524 3176
rect 9727 3148 9772 3176
rect 8076 3136 8082 3148
rect 4249 3111 4307 3117
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 8496 3108 8524 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 11701 3179 11759 3185
rect 11701 3176 11713 3179
rect 9876 3148 11713 3176
rect 9876 3108 9904 3148
rect 11701 3145 11713 3148
rect 11747 3145 11759 3179
rect 11701 3139 11759 3145
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 12345 3179 12403 3185
rect 12345 3176 12357 3179
rect 11848 3148 12357 3176
rect 11848 3136 11854 3148
rect 12345 3145 12357 3148
rect 12391 3176 12403 3179
rect 13538 3176 13544 3188
rect 12391 3148 13544 3176
rect 12391 3145 12403 3148
rect 12345 3139 12403 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 16574 3176 16580 3188
rect 14568 3148 16580 3176
rect 4295 3080 8432 3108
rect 8496 3080 9904 3108
rect 10321 3111 10379 3117
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 4062 3040 4068 3052
rect 3743 3012 4068 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 4062 3000 4068 3012
rect 4120 3040 4126 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 4120 3012 4169 3040
rect 4120 3000 4126 3012
rect 4157 3009 4169 3012
rect 4203 3040 4215 3043
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4203 3012 4813 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8018 3040 8024 3052
rect 7607 3012 8024 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 4816 2972 4844 3003
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 4816 2944 7389 2972
rect 7377 2941 7389 2944
rect 7423 2972 7435 2975
rect 7926 2972 7932 2984
rect 7423 2944 7932 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8297 2975 8355 2981
rect 8297 2941 8309 2975
rect 8343 2941 8355 2975
rect 8404 2972 8432 3080
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 10502 3108 10508 3120
rect 10367 3080 10508 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 10873 3111 10931 3117
rect 10873 3108 10885 3111
rect 10744 3080 10885 3108
rect 10744 3068 10750 3080
rect 10873 3077 10885 3080
rect 10919 3077 10931 3111
rect 10873 3071 10931 3077
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 11020 3080 12650 3108
rect 11020 3068 11026 3080
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 13817 3111 13875 3117
rect 13817 3108 13829 3111
rect 13780 3080 13829 3108
rect 13780 3068 13786 3080
rect 13817 3077 13829 3080
rect 13863 3077 13875 3111
rect 13817 3071 13875 3077
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 10100 3012 10241 3040
rect 10100 3000 10106 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10229 3003 10287 3009
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 11606 3040 11612 3052
rect 11112 3012 11612 3040
rect 11112 3000 11118 3012
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11882 3000 11888 3012
rect 11940 3040 11946 3052
rect 12434 3040 12440 3052
rect 11940 3012 12440 3040
rect 11940 3000 11946 3012
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14568 3049 14596 3148
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 19426 3176 19432 3188
rect 16724 3148 19432 3176
rect 16724 3136 16730 3148
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 22922 3176 22928 3188
rect 19720 3148 22048 3176
rect 16114 3108 16120 3120
rect 16054 3080 16120 3108
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 17218 3108 17224 3120
rect 16224 3080 17224 3108
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14148 3012 14565 3040
rect 14148 3000 14154 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 12526 2972 12532 2984
rect 8404 2944 12532 2972
rect 8297 2935 8355 2941
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 4706 2904 4712 2916
rect 3191 2876 4712 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 4893 2907 4951 2913
rect 4893 2873 4905 2907
rect 4939 2904 4951 2907
rect 5902 2904 5908 2916
rect 4939 2876 5908 2904
rect 4939 2873 4951 2876
rect 4893 2867 4951 2873
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 8202 2904 8208 2916
rect 6788 2876 8208 2904
rect 6788 2864 6794 2876
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8312 2904 8340 2935
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 13872 2944 14841 2972
rect 13872 2932 13878 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 8312 2876 12434 2904
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 5994 2836 6000 2848
rect 5955 2808 6000 2836
rect 5994 2796 6000 2808
rect 6052 2836 6058 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6052 2808 6561 2836
rect 6052 2796 6058 2808
rect 6549 2805 6561 2808
rect 6595 2836 6607 2839
rect 6914 2836 6920 2848
rect 6595 2808 6920 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8444 2808 9137 2836
rect 8444 2796 8450 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 11882 2836 11888 2848
rect 9640 2808 11888 2836
rect 9640 2796 9646 2808
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12406 2836 12434 2876
rect 16224 2836 16252 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 19150 3108 19156 3120
rect 18354 3080 19156 3108
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 16574 3000 16580 3052
rect 16632 3040 16638 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16632 3012 16865 3040
rect 16632 3000 16638 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 19245 3043 19303 3049
rect 19245 3009 19257 3043
rect 19291 3040 19303 3043
rect 19426 3040 19432 3052
rect 19291 3012 19432 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 19426 3000 19432 3012
rect 19484 3040 19490 3052
rect 19720 3049 19748 3148
rect 19981 3111 20039 3117
rect 19981 3077 19993 3111
rect 20027 3108 20039 3111
rect 20070 3108 20076 3120
rect 20027 3080 20076 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 22020 3108 22048 3148
rect 22296 3148 22928 3176
rect 22296 3120 22324 3148
rect 22922 3136 22928 3148
rect 22980 3136 22986 3188
rect 23753 3179 23811 3185
rect 23753 3145 23765 3179
rect 23799 3176 23811 3179
rect 24210 3176 24216 3188
rect 23799 3148 24216 3176
rect 23799 3145 23811 3148
rect 23753 3139 23811 3145
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 26142 3176 26148 3188
rect 24728 3148 26148 3176
rect 24728 3136 24734 3148
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 31573 3179 31631 3185
rect 31573 3176 31585 3179
rect 27264 3148 31585 3176
rect 22186 3108 22192 3120
rect 22020 3080 22192 3108
rect 22020 3049 22048 3080
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22278 3068 22284 3120
rect 22336 3108 22342 3120
rect 24394 3108 24400 3120
rect 22336 3080 22429 3108
rect 23506 3080 24400 3108
rect 22336 3068 22342 3080
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 27264 3108 27292 3148
rect 31573 3145 31585 3148
rect 31619 3145 31631 3179
rect 38102 3176 38108 3188
rect 31573 3139 31631 3145
rect 31726 3148 38108 3176
rect 31726 3108 31754 3148
rect 38102 3136 38108 3148
rect 38160 3136 38166 3188
rect 25254 3080 27292 3108
rect 28276 3080 31754 3108
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19484 3012 19717 3040
rect 19484 3000 19490 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 22005 3043 22063 3049
rect 19705 3003 19763 3009
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 18874 2972 18880 2984
rect 17175 2944 18880 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 19058 2904 19064 2916
rect 18248 2876 19064 2904
rect 12406 2808 16252 2836
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 18248 2836 18276 2876
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 21100 2904 21128 3026
rect 22005 3009 22017 3043
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 25961 3043 26019 3049
rect 25961 3009 25973 3043
rect 26007 3040 26019 3043
rect 26142 3040 26148 3052
rect 26007 3012 26148 3040
rect 26007 3009 26019 3012
rect 25961 3003 26019 3009
rect 26142 3000 26148 3012
rect 26200 3000 26206 3052
rect 26602 3040 26608 3052
rect 26563 3012 26608 3040
rect 26602 3000 26608 3012
rect 26660 3000 26666 3052
rect 27706 3040 27712 3052
rect 26712 3012 27712 3040
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 22278 2972 22284 2984
rect 21499 2944 22284 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 22370 2932 22376 2984
rect 22428 2972 22434 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 22428 2944 24225 2972
rect 22428 2932 22434 2944
rect 24213 2941 24225 2944
rect 24259 2972 24271 2975
rect 25314 2972 25320 2984
rect 24259 2944 25320 2972
rect 24259 2941 24271 2944
rect 24213 2935 24271 2941
rect 25314 2932 25320 2944
rect 25372 2932 25378 2984
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 25648 2944 25697 2972
rect 25648 2932 25654 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 25685 2935 25743 2941
rect 26050 2932 26056 2984
rect 26108 2972 26114 2984
rect 26712 2972 26740 3012
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 28276 3049 28304 3080
rect 28261 3043 28319 3049
rect 28261 3009 28273 3043
rect 28307 3009 28319 3043
rect 28261 3003 28319 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 29089 3041 29147 3047
rect 28868 3038 28948 3040
rect 29089 3038 29101 3041
rect 28868 3012 29101 3038
rect 28868 3000 28874 3012
rect 28920 3010 29101 3012
rect 29089 3007 29101 3010
rect 29135 3007 29147 3041
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 29089 3001 29147 3007
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 30392 3049 30420 3080
rect 31846 3068 31852 3120
rect 31904 3108 31910 3120
rect 33686 3108 33692 3120
rect 31904 3080 33088 3108
rect 33647 3080 33692 3108
rect 31904 3068 31910 3080
rect 30377 3043 30435 3049
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30926 3040 30932 3052
rect 30887 3012 30932 3040
rect 30377 3003 30435 3009
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31665 3043 31723 3049
rect 31665 3040 31677 3043
rect 31076 3012 31677 3040
rect 31076 3000 31082 3012
rect 31665 3009 31677 3012
rect 31711 3040 31723 3043
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 31711 3012 32505 3040
rect 31711 3009 31723 3012
rect 31665 3003 31723 3009
rect 32493 3009 32505 3012
rect 32539 3009 32551 3043
rect 33060 3040 33088 3080
rect 33686 3068 33692 3080
rect 33744 3068 33750 3120
rect 36262 3108 36268 3120
rect 36223 3080 36268 3108
rect 36262 3068 36268 3080
rect 36320 3068 36326 3120
rect 33129 3043 33187 3049
rect 33129 3040 33141 3043
rect 33060 3012 33141 3040
rect 32493 3003 32551 3009
rect 33129 3009 33141 3012
rect 33175 3009 33187 3043
rect 33129 3003 33187 3009
rect 33781 3043 33839 3049
rect 33781 3009 33793 3043
rect 33827 3040 33839 3043
rect 33870 3040 33876 3052
rect 33827 3012 33876 3040
rect 33827 3009 33839 3012
rect 33781 3003 33839 3009
rect 33870 3000 33876 3012
rect 33928 3000 33934 3052
rect 34422 3040 34428 3052
rect 34335 3012 34428 3040
rect 34422 3000 34428 3012
rect 34480 3040 34486 3052
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34480 3012 35081 3040
rect 34480 3000 34486 3012
rect 35069 3009 35081 3012
rect 35115 3040 35127 3043
rect 35115 3012 35664 3040
rect 35115 3009 35127 3012
rect 35069 3003 35127 3009
rect 26108 2944 26740 2972
rect 27617 2975 27675 2981
rect 26108 2932 26114 2944
rect 27617 2941 27629 2975
rect 27663 2941 27675 2975
rect 27617 2935 27675 2941
rect 21100 2876 22048 2904
rect 16347 2808 18276 2836
rect 18601 2839 18659 2845
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 18601 2805 18613 2839
rect 18647 2836 18659 2839
rect 21910 2836 21916 2848
rect 18647 2808 21916 2836
rect 18647 2805 18659 2808
rect 18601 2799 18659 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22020 2836 22048 2876
rect 24118 2864 24124 2916
rect 24176 2904 24182 2916
rect 27157 2907 27215 2913
rect 27157 2904 27169 2907
rect 24176 2876 24532 2904
rect 24176 2864 24182 2876
rect 24504 2848 24532 2876
rect 26252 2876 27169 2904
rect 23658 2836 23664 2848
rect 22020 2808 23664 2836
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 24486 2796 24492 2848
rect 24544 2796 24550 2848
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 26252 2836 26280 2876
rect 27157 2873 27169 2876
rect 27203 2873 27215 2907
rect 27632 2904 27660 2935
rect 27798 2932 27804 2984
rect 27856 2972 27862 2984
rect 30285 2975 30343 2981
rect 30285 2972 30297 2975
rect 27856 2944 30297 2972
rect 27856 2932 27862 2944
rect 30285 2941 30297 2944
rect 30331 2941 30343 2975
rect 30285 2935 30343 2941
rect 30558 2932 30564 2984
rect 30616 2972 30622 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 30616 2944 35541 2972
rect 30616 2932 30622 2944
rect 35529 2941 35541 2944
rect 35575 2941 35587 2975
rect 35636 2972 35664 3012
rect 36446 3000 36452 3052
rect 36504 3040 36510 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36504 3012 36553 3040
rect 36504 3000 36510 3012
rect 36541 3009 36553 3012
rect 36587 3040 36599 3043
rect 36906 3040 36912 3052
rect 36587 3012 36912 3040
rect 36587 3009 36599 3012
rect 36541 3003 36599 3009
rect 36906 3000 36912 3012
rect 36964 3040 36970 3052
rect 37461 3043 37519 3049
rect 37461 3040 37473 3043
rect 36964 3012 37473 3040
rect 36964 3000 36970 3012
rect 37461 3009 37473 3012
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 37645 2975 37703 2981
rect 37645 2972 37657 2975
rect 35636 2944 37657 2972
rect 35529 2935 35587 2941
rect 37645 2941 37657 2944
rect 37691 2941 37703 2975
rect 37645 2935 37703 2941
rect 29641 2907 29699 2913
rect 29641 2904 29653 2907
rect 27632 2876 29653 2904
rect 27157 2867 27215 2873
rect 29641 2873 29653 2876
rect 29687 2873 29699 2907
rect 32398 2904 32404 2916
rect 32359 2876 32404 2904
rect 29641 2867 29699 2873
rect 32398 2864 32404 2876
rect 32456 2864 32462 2916
rect 32490 2864 32496 2916
rect 32548 2904 32554 2916
rect 34333 2907 34391 2913
rect 34333 2904 34345 2907
rect 32548 2876 34345 2904
rect 32548 2864 32554 2876
rect 34333 2873 34345 2876
rect 34379 2873 34391 2907
rect 34333 2867 34391 2873
rect 26510 2836 26516 2848
rect 25096 2808 26280 2836
rect 26471 2808 26516 2836
rect 25096 2796 25102 2808
rect 26510 2796 26516 2808
rect 26568 2796 26574 2848
rect 26602 2796 26608 2848
rect 26660 2836 26666 2848
rect 28074 2836 28080 2848
rect 26660 2808 28080 2836
rect 26660 2796 26666 2808
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28445 2839 28503 2845
rect 28445 2805 28457 2839
rect 28491 2836 28503 2839
rect 28810 2836 28816 2848
rect 28491 2808 28816 2836
rect 28491 2805 28503 2808
rect 28445 2799 28503 2805
rect 28810 2796 28816 2808
rect 28868 2796 28874 2848
rect 28994 2796 29000 2848
rect 29052 2836 29058 2848
rect 29052 2808 29097 2836
rect 29052 2796 29058 2808
rect 31202 2796 31208 2848
rect 31260 2836 31266 2848
rect 32306 2836 32312 2848
rect 31260 2808 32312 2836
rect 31260 2796 31266 2808
rect 32306 2796 32312 2808
rect 32364 2796 32370 2848
rect 33042 2836 33048 2848
rect 33003 2808 33048 2836
rect 33042 2796 33048 2808
rect 33100 2796 33106 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34977 2839 35035 2845
rect 34977 2836 34989 2839
rect 34572 2808 34989 2836
rect 34572 2796 34578 2808
rect 34977 2805 34989 2808
rect 35023 2805 35035 2839
rect 34977 2799 35035 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 5994 2632 6000 2644
rect 5955 2604 6000 2632
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 6972 2604 7481 2632
rect 6972 2592 6978 2604
rect 7469 2601 7481 2604
rect 7515 2632 7527 2635
rect 9217 2635 9275 2641
rect 9217 2632 9229 2635
rect 7515 2604 9229 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 9217 2601 9229 2604
rect 9263 2601 9275 2635
rect 31478 2632 31484 2644
rect 9217 2595 9275 2601
rect 10060 2604 31484 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 4203 2536 5856 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 5442 2496 5448 2508
rect 2608 2468 5448 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2406 2428 2412 2440
rect 1903 2400 2412 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2608 2437 2636 2468
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5828 2496 5856 2536
rect 5902 2524 5908 2576
rect 5960 2564 5966 2576
rect 5960 2536 9904 2564
rect 5960 2524 5966 2536
rect 6730 2496 6736 2508
rect 5828 2468 6736 2496
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 6840 2468 9076 2496
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3292 2400 3985 2428
rect 3292 2388 3298 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 3973 2391 4031 2397
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 6840 2437 6868 2468
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 8018 2428 8024 2440
rect 7979 2400 8024 2428
rect 6825 2391 6883 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2360 4951 2363
rect 8202 2360 8208 2372
rect 4939 2332 8208 2360
rect 4939 2329 4951 2332
rect 4893 2323 4951 2329
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 8297 2363 8355 2369
rect 8297 2329 8309 2363
rect 8343 2329 8355 2363
rect 9048 2360 9076 2468
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9876 2428 9904 2536
rect 10060 2505 10088 2604
rect 31478 2592 31484 2604
rect 31536 2592 31542 2644
rect 33137 2635 33195 2641
rect 33137 2601 33149 2635
rect 33183 2632 33195 2635
rect 34330 2632 34336 2644
rect 33183 2604 34336 2632
rect 33183 2601 33195 2604
rect 33137 2595 33195 2601
rect 34330 2592 34336 2604
rect 34388 2592 34394 2644
rect 35802 2632 35808 2644
rect 35763 2604 35808 2632
rect 35802 2592 35808 2604
rect 35860 2592 35866 2644
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11330 2564 11336 2576
rect 11195 2536 11336 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 11977 2567 12035 2573
rect 11977 2533 11989 2567
rect 12023 2564 12035 2567
rect 12250 2564 12256 2576
rect 12023 2536 12256 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 16850 2524 16856 2576
rect 16908 2564 16914 2576
rect 17129 2567 17187 2573
rect 17129 2564 17141 2567
rect 16908 2536 17141 2564
rect 16908 2524 16914 2536
rect 17129 2533 17141 2536
rect 17175 2533 17187 2567
rect 17129 2527 17187 2533
rect 21174 2524 21180 2576
rect 21232 2564 21238 2576
rect 21269 2567 21327 2573
rect 21269 2564 21281 2567
rect 21232 2536 21281 2564
rect 21232 2524 21238 2536
rect 21269 2533 21281 2536
rect 21315 2533 21327 2567
rect 30466 2564 30472 2576
rect 21269 2527 21327 2533
rect 23492 2536 30472 2564
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 14090 2496 14096 2508
rect 13771 2468 14096 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14090 2456 14096 2468
rect 14148 2496 14154 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 14148 2468 14565 2496
rect 14148 2456 14154 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15838 2496 15844 2508
rect 14875 2468 15844 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 17310 2496 17316 2508
rect 16347 2468 17316 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 19426 2496 19432 2508
rect 18923 2468 19432 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 19426 2456 19432 2468
rect 19484 2496 19490 2508
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 19484 2468 19533 2496
rect 19484 2456 19490 2468
rect 19521 2465 19533 2468
rect 19567 2496 19579 2499
rect 19886 2496 19892 2508
rect 19567 2468 19892 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 22094 2496 22100 2508
rect 22055 2468 22100 2496
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 22373 2499 22431 2505
rect 22373 2465 22385 2499
rect 22419 2496 22431 2499
rect 23382 2496 23388 2508
rect 22419 2468 23388 2496
rect 22419 2465 22431 2468
rect 22373 2459 22431 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 9876 2400 12374 2428
rect 23492 2414 23520 2536
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 32306 2564 32312 2576
rect 32267 2536 32312 2564
rect 32306 2524 32312 2536
rect 32364 2524 32370 2576
rect 33502 2524 33508 2576
rect 33560 2564 33566 2576
rect 33597 2567 33655 2573
rect 33597 2564 33609 2567
rect 33560 2536 33609 2564
rect 33560 2524 33566 2536
rect 33597 2533 33609 2536
rect 33643 2533 33655 2567
rect 33597 2527 33655 2533
rect 23845 2499 23903 2505
rect 23845 2465 23857 2499
rect 23891 2496 23903 2499
rect 24486 2496 24492 2508
rect 23891 2468 24492 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 24486 2456 24492 2468
rect 24544 2456 24550 2508
rect 25038 2496 25044 2508
rect 24999 2468 25044 2496
rect 25038 2456 25044 2468
rect 25096 2456 25102 2508
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2496 25559 2499
rect 26510 2496 26516 2508
rect 25547 2468 26516 2496
rect 25547 2465 25559 2468
rect 25501 2459 25559 2465
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 28258 2496 28264 2508
rect 26988 2468 28264 2496
rect 25685 2431 25743 2437
rect 9769 2391 9827 2397
rect 25685 2397 25697 2431
rect 25731 2428 25743 2431
rect 26326 2428 26332 2440
rect 25731 2400 26332 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 26988 2428 27016 2468
rect 28258 2456 28264 2468
rect 28316 2456 28322 2508
rect 30558 2496 30564 2508
rect 28736 2468 30564 2496
rect 27154 2428 27160 2440
rect 26467 2400 27016 2428
rect 27115 2400 27160 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27154 2388 27160 2400
rect 27212 2388 27218 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28736 2437 28764 2468
rect 30558 2456 30564 2468
rect 30616 2456 30622 2508
rect 31386 2496 31392 2508
rect 30668 2468 31392 2496
rect 28721 2431 28779 2437
rect 28721 2428 28733 2431
rect 28408 2400 28733 2428
rect 28408 2388 28414 2400
rect 28721 2397 28733 2400
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 30668 2437 30696 2468
rect 31386 2456 31392 2468
rect 31444 2456 31450 2508
rect 32214 2496 32220 2508
rect 31496 2468 32220 2496
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 28960 2400 29745 2428
rect 28960 2388 28966 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2428 31355 2431
rect 31496 2428 31524 2468
rect 32214 2456 32220 2468
rect 32272 2456 32278 2508
rect 33870 2456 33876 2508
rect 33928 2496 33934 2508
rect 36633 2499 36691 2505
rect 36633 2496 36645 2499
rect 33928 2468 36645 2496
rect 33928 2456 33934 2468
rect 36633 2465 36645 2468
rect 36679 2465 36691 2499
rect 36633 2459 36691 2465
rect 37461 2499 37519 2505
rect 37461 2465 37473 2499
rect 37507 2496 37519 2499
rect 37642 2496 37648 2508
rect 37507 2468 37648 2496
rect 37507 2465 37519 2468
rect 37461 2459 37519 2465
rect 37642 2456 37648 2468
rect 37700 2456 37706 2508
rect 31343 2400 31524 2428
rect 31343 2397 31355 2400
rect 31297 2391 31355 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 31628 2400 32505 2428
rect 31628 2388 31634 2400
rect 32493 2397 32505 2400
rect 32539 2428 32551 2431
rect 32582 2428 32588 2440
rect 32539 2400 32588 2428
rect 32539 2397 32551 2400
rect 32493 2391 32551 2397
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 33560 2400 33793 2428
rect 33560 2388 33566 2400
rect 33781 2397 33793 2400
rect 33827 2428 33839 2431
rect 33962 2428 33968 2440
rect 33827 2400 33968 2428
rect 33827 2397 33839 2400
rect 33781 2391 33839 2397
rect 33962 2388 33968 2400
rect 34020 2388 34026 2440
rect 35161 2431 35219 2437
rect 35161 2397 35173 2431
rect 35207 2428 35219 2431
rect 35434 2428 35440 2440
rect 35207 2400 35440 2428
rect 35207 2397 35219 2400
rect 35161 2391 35219 2397
rect 35434 2388 35440 2400
rect 35492 2388 35498 2440
rect 35897 2431 35955 2437
rect 35897 2397 35909 2431
rect 35943 2428 35955 2431
rect 36078 2428 36084 2440
rect 35943 2400 36084 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 36078 2388 36084 2400
rect 36136 2428 36142 2440
rect 36722 2428 36728 2440
rect 36136 2400 36728 2428
rect 36136 2388 36142 2400
rect 36722 2388 36728 2400
rect 36780 2388 36786 2440
rect 36906 2428 36912 2440
rect 36867 2400 36912 2428
rect 36906 2388 36912 2400
rect 36964 2388 36970 2440
rect 37734 2428 37740 2440
rect 37695 2400 37740 2428
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 11146 2360 11152 2372
rect 9048 2332 11152 2360
rect 8297 2323 8355 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 1673 2255 1731 2261
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 8312 2292 8340 2323
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 13446 2360 13452 2372
rect 13407 2332 13452 2360
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 15286 2320 15292 2372
rect 15344 2320 15350 2372
rect 17862 2320 17868 2372
rect 17920 2320 17926 2372
rect 18601 2363 18659 2369
rect 18601 2329 18613 2363
rect 18647 2360 18659 2363
rect 19058 2360 19064 2372
rect 18647 2332 19064 2360
rect 18647 2329 18659 2332
rect 18601 2323 18659 2329
rect 19058 2320 19064 2332
rect 19116 2320 19122 2372
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 19797 2363 19855 2369
rect 19797 2360 19809 2363
rect 19392 2332 19809 2360
rect 19392 2320 19398 2332
rect 19797 2329 19809 2332
rect 19843 2329 19855 2363
rect 22278 2360 22284 2372
rect 21022 2332 22284 2360
rect 19797 2323 19855 2329
rect 11238 2292 11244 2304
rect 8312 2264 11244 2292
rect 6641 2255 6699 2261
rect 11238 2252 11244 2264
rect 11296 2292 11302 2304
rect 16666 2292 16672 2304
rect 11296 2264 16672 2292
rect 11296 2252 11302 2264
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 19812 2292 19840 2323
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 26142 2320 26148 2372
rect 26200 2360 26206 2372
rect 27893 2363 27951 2369
rect 27893 2360 27905 2363
rect 26200 2332 27905 2360
rect 26200 2320 26206 2332
rect 27893 2329 27905 2332
rect 27939 2329 27951 2363
rect 27893 2323 27951 2329
rect 20622 2292 20628 2304
rect 19812 2264 20628 2292
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 25188 2264 26249 2292
rect 25188 2252 25194 2264
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 26237 2255 26295 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 26476 2264 27353 2292
rect 26476 2252 26482 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 28442 2252 28448 2304
rect 28500 2292 28506 2304
rect 28537 2295 28595 2301
rect 28537 2292 28549 2295
rect 28500 2264 28549 2292
rect 28500 2252 28506 2264
rect 28537 2261 28549 2264
rect 28583 2261 28595 2295
rect 28537 2255 28595 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 30558 2292 30564 2304
rect 30519 2264 30564 2292
rect 29917 2255 29975 2261
rect 30558 2252 30564 2264
rect 30616 2252 30622 2304
rect 31202 2292 31208 2304
rect 31163 2264 31208 2292
rect 31202 2252 31208 2264
rect 31260 2252 31266 2304
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 34977 2295 35035 2301
rect 34977 2292 34989 2295
rect 34848 2264 34989 2292
rect 34848 2252 34854 2264
rect 34977 2261 34989 2264
rect 35023 2261 35035 2295
rect 34977 2255 35035 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 9674 2088 9680 2100
rect 3476 2060 9680 2088
rect 3476 2048 3482 2060
rect 9674 2048 9680 2060
rect 9732 2048 9738 2100
rect 24578 2048 24584 2100
rect 24636 2088 24642 2100
rect 27154 2088 27160 2100
rect 24636 2060 27160 2088
rect 24636 2048 24642 2060
rect 27154 2048 27160 2060
rect 27212 2048 27218 2100
rect 28166 2048 28172 2100
rect 28224 2088 28230 2100
rect 28224 2060 35894 2088
rect 28224 2048 28230 2060
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 10594 2020 10600 2032
rect 8260 1992 10600 2020
rect 8260 1980 8266 1992
rect 10594 1980 10600 1992
rect 10652 1980 10658 2032
rect 24946 1980 24952 2032
rect 25004 2020 25010 2032
rect 30558 2020 30564 2032
rect 25004 1992 30564 2020
rect 25004 1980 25010 1992
rect 30558 1980 30564 1992
rect 30616 1980 30622 2032
rect 5442 1912 5448 1964
rect 5500 1952 5506 1964
rect 15286 1952 15292 1964
rect 5500 1924 15292 1952
rect 5500 1912 5506 1924
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 25774 1912 25780 1964
rect 25832 1952 25838 1964
rect 31202 1952 31208 1964
rect 25832 1924 31208 1952
rect 25832 1912 25838 1924
rect 31202 1912 31208 1924
rect 31260 1912 31266 1964
rect 35866 1952 35894 2060
rect 37734 1952 37740 1964
rect 35866 1924 37740 1952
rect 37734 1912 37740 1924
rect 37792 1912 37798 1964
rect 22278 1844 22284 1896
rect 22336 1884 22342 1896
rect 33042 1884 33048 1896
rect 22336 1856 33048 1884
rect 22336 1844 22342 1856
rect 33042 1844 33048 1856
rect 33100 1844 33106 1896
rect 20530 1776 20536 1828
rect 20588 1816 20594 1828
rect 24302 1816 24308 1828
rect 20588 1788 24308 1816
rect 20588 1776 20594 1788
rect 24302 1776 24308 1788
rect 24360 1816 24366 1828
rect 32214 1816 32220 1828
rect 24360 1788 32220 1816
rect 24360 1776 24366 1788
rect 32214 1776 32220 1788
rect 32272 1776 32278 1828
<< via1 >>
rect 2964 37612 3016 37664
rect 21824 37612 21876 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2964 37451 3016 37460
rect 2964 37417 2973 37451
rect 2973 37417 3007 37451
rect 3007 37417 3016 37451
rect 2964 37408 3016 37417
rect 13544 37408 13596 37460
rect 23020 37408 23072 37460
rect 35440 37408 35492 37460
rect 36728 37451 36780 37460
rect 36728 37417 36737 37451
rect 36737 37417 36771 37451
rect 36771 37417 36780 37451
rect 36728 37408 36780 37417
rect 20536 37340 20588 37392
rect 7104 37272 7156 37324
rect 1952 37204 2004 37256
rect 2872 37247 2924 37256
rect 2872 37213 2881 37247
rect 2881 37213 2915 37247
rect 2915 37213 2924 37247
rect 2872 37204 2924 37213
rect 5264 37247 5316 37256
rect 5264 37213 5273 37247
rect 5273 37213 5307 37247
rect 5307 37213 5316 37247
rect 5264 37204 5316 37213
rect 13544 37272 13596 37324
rect 20628 37315 20680 37324
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 10692 37247 10744 37256
rect 10692 37213 10701 37247
rect 10701 37213 10735 37247
rect 10735 37213 10744 37247
rect 10692 37204 10744 37213
rect 14280 37204 14332 37256
rect 20628 37281 20637 37315
rect 20637 37281 20671 37315
rect 20671 37281 20680 37315
rect 20628 37272 20680 37281
rect 15844 37247 15896 37256
rect 15844 37213 15853 37247
rect 15853 37213 15887 37247
rect 15887 37213 15896 37247
rect 15844 37204 15896 37213
rect 17132 37247 17184 37256
rect 17132 37213 17141 37247
rect 17141 37213 17175 37247
rect 17175 37213 17184 37247
rect 17132 37204 17184 37213
rect 18420 37204 18472 37256
rect 9496 37136 9548 37188
rect 19340 37136 19392 37188
rect 21272 37204 21324 37256
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 25228 37136 25280 37188
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 30748 37247 30800 37256
rect 30748 37213 30757 37247
rect 30757 37213 30791 37247
rect 30791 37213 30800 37247
rect 30748 37204 30800 37213
rect 33600 37247 33652 37256
rect 30656 37136 30708 37188
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 35440 37204 35492 37256
rect 36912 37247 36964 37256
rect 36912 37213 36921 37247
rect 36921 37213 36955 37247
rect 36955 37213 36964 37247
rect 36912 37204 36964 37213
rect 37464 37247 37516 37256
rect 37464 37213 37473 37247
rect 37473 37213 37507 37247
rect 37507 37213 37516 37247
rect 37464 37204 37516 37213
rect 35532 37179 35584 37188
rect 35532 37145 35541 37179
rect 35541 37145 35575 37179
rect 35575 37145 35584 37179
rect 35532 37136 35584 37145
rect 3884 37068 3936 37120
rect 5172 37068 5224 37120
rect 7380 37111 7432 37120
rect 7380 37077 7389 37111
rect 7389 37077 7423 37111
rect 7423 37077 7432 37111
rect 7380 37068 7432 37077
rect 8392 37068 8444 37120
rect 10324 37068 10376 37120
rect 12440 37111 12492 37120
rect 12440 37077 12449 37111
rect 12449 37077 12483 37111
rect 12483 37077 12492 37111
rect 12440 37068 12492 37077
rect 15476 37068 15528 37120
rect 16764 37068 16816 37120
rect 19432 37068 19484 37120
rect 22100 37068 22152 37120
rect 23848 37068 23900 37120
rect 25136 37068 25188 37120
rect 27068 37068 27120 37120
rect 29000 37068 29052 37120
rect 30380 37068 30432 37120
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2872 36864 2924 36916
rect 10692 36864 10744 36916
rect 14280 36864 14332 36916
rect 20536 36907 20588 36916
rect 20536 36873 20545 36907
rect 20545 36873 20579 36907
rect 20579 36873 20588 36907
rect 20536 36864 20588 36873
rect 21272 36907 21324 36916
rect 21272 36873 21281 36907
rect 21281 36873 21315 36907
rect 21315 36873 21324 36907
rect 21272 36864 21324 36873
rect 1676 36771 1728 36780
rect 1676 36737 1685 36771
rect 1685 36737 1719 36771
rect 1719 36737 1728 36771
rect 1676 36728 1728 36737
rect 19340 36728 19392 36780
rect 23020 36796 23072 36848
rect 21824 36728 21876 36780
rect 22008 36771 22060 36780
rect 22008 36737 22017 36771
rect 22017 36737 22051 36771
rect 22051 36737 22060 36771
rect 22008 36728 22060 36737
rect 38660 36796 38712 36848
rect 18788 36660 18840 36712
rect 25320 36660 25372 36712
rect 35532 36660 35584 36712
rect 1768 36567 1820 36576
rect 1768 36533 1777 36567
rect 1777 36533 1811 36567
rect 1811 36533 1820 36567
rect 1768 36524 1820 36533
rect 37464 36660 37516 36712
rect 37924 36592 37976 36644
rect 29736 36524 29788 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 20 36320 72 36372
rect 1768 36320 1820 36372
rect 13820 36320 13872 36372
rect 38200 36363 38252 36372
rect 38200 36329 38209 36363
rect 38209 36329 38243 36363
rect 38243 36329 38252 36363
rect 38200 36320 38252 36329
rect 1952 36252 2004 36304
rect 5448 36116 5500 36168
rect 37740 36116 37792 36168
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 18696 35776 18748 35828
rect 19432 35776 19484 35828
rect 27896 35436 27948 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 18420 34187 18472 34196
rect 18420 34153 18429 34187
rect 18429 34153 18463 34187
rect 18463 34153 18472 34187
rect 18420 34144 18472 34153
rect 17684 33847 17736 33856
rect 17684 33813 17693 33847
rect 17693 33813 17727 33847
rect 17727 33813 17736 33847
rect 17684 33804 17736 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 38200 33507 38252 33516
rect 38200 33473 38209 33507
rect 38209 33473 38243 33507
rect 38243 33473 38252 33507
rect 38200 33464 38252 33473
rect 9312 33328 9364 33380
rect 26148 33260 26200 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1676 33099 1728 33108
rect 1676 33065 1685 33099
rect 1685 33065 1719 33099
rect 1719 33065 1728 33099
rect 1676 33056 1728 33065
rect 5264 33056 5316 33108
rect 5448 32784 5500 32836
rect 9220 32716 9272 32768
rect 25504 32716 25556 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15844 32172 15896 32224
rect 38108 32376 38160 32428
rect 28632 32172 28684 32224
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 9496 31968 9548 32020
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 10508 31807 10560 31816
rect 10508 31773 10517 31807
rect 10517 31773 10551 31807
rect 10551 31773 10560 31807
rect 10508 31764 10560 31773
rect 30104 31764 30156 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31399 1636 31408
rect 1584 31365 1593 31399
rect 1593 31365 1627 31399
rect 1627 31365 1636 31399
rect 1584 31356 1636 31365
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 38016 30812 38068 30864
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19340 30200 19392 30252
rect 38016 30243 38068 30252
rect 38016 30209 38025 30243
rect 38025 30209 38059 30243
rect 38059 30209 38068 30243
rect 38016 30200 38068 30209
rect 1584 30175 1636 30184
rect 1584 30141 1593 30175
rect 1593 30141 1627 30175
rect 1627 30141 1636 30175
rect 1584 30132 1636 30141
rect 2504 30132 2556 30184
rect 19340 29996 19392 30048
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 24584 29248 24636 29300
rect 30748 29248 30800 29300
rect 12072 29112 12124 29164
rect 30932 29155 30984 29164
rect 30932 29121 30941 29155
rect 30941 29121 30975 29155
rect 30975 29121 30984 29155
rect 30932 29112 30984 29121
rect 34152 29112 34204 29164
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 30656 28203 30708 28212
rect 30656 28169 30665 28203
rect 30665 28169 30699 28203
rect 30699 28169 30708 28203
rect 30656 28160 30708 28169
rect 1860 28067 1912 28076
rect 1860 28033 1869 28067
rect 1869 28033 1903 28067
rect 1903 28033 1912 28067
rect 1860 28024 1912 28033
rect 31208 28024 31260 28076
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 31208 27863 31260 27872
rect 31208 27829 31217 27863
rect 31217 27829 31251 27863
rect 31251 27829 31260 27863
rect 31208 27820 31260 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 23020 27591 23072 27600
rect 23020 27557 23029 27591
rect 23029 27557 23063 27591
rect 23063 27557 23072 27591
rect 23020 27548 23072 27557
rect 22100 27276 22152 27328
rect 38292 27319 38344 27328
rect 38292 27285 38301 27319
rect 38301 27285 38335 27319
rect 38335 27285 38344 27319
rect 38292 27276 38344 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 18788 27115 18840 27124
rect 18788 27081 18797 27115
rect 18797 27081 18831 27115
rect 18831 27081 18840 27115
rect 18788 27072 18840 27081
rect 6828 26936 6880 26988
rect 20536 26868 20588 26920
rect 37372 26868 37424 26920
rect 38292 26911 38344 26920
rect 38292 26877 38301 26911
rect 38301 26877 38335 26911
rect 38335 26877 38344 26911
rect 38292 26868 38344 26877
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 15660 26732 15712 26784
rect 18328 26732 18380 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9404 26528 9456 26580
rect 22008 26528 22060 26580
rect 36912 26528 36964 26580
rect 38016 26367 38068 26376
rect 38016 26333 38025 26367
rect 38025 26333 38059 26367
rect 38059 26333 38068 26367
rect 38016 26324 38068 26333
rect 18144 26256 18196 26308
rect 20076 26256 20128 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 33600 26027 33652 26036
rect 33600 25993 33609 26027
rect 33609 25993 33643 26027
rect 33643 25993 33652 26027
rect 33600 25984 33652 25993
rect 34244 25848 34296 25900
rect 34244 25687 34296 25696
rect 34244 25653 34253 25687
rect 34253 25653 34287 25687
rect 34287 25653 34296 25687
rect 34244 25644 34296 25653
rect 38016 25644 38068 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 38200 25440 38252 25492
rect 37832 25279 37884 25288
rect 37832 25245 37841 25279
rect 37841 25245 37875 25279
rect 37875 25245 37884 25279
rect 37832 25236 37884 25245
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 37464 24896 37516 24948
rect 38016 24896 38068 24948
rect 25504 24828 25556 24880
rect 26700 24828 26752 24880
rect 21640 24760 21692 24812
rect 37924 24760 37976 24812
rect 38108 24760 38160 24812
rect 1676 24599 1728 24608
rect 1676 24565 1685 24599
rect 1685 24565 1719 24599
rect 1719 24565 1728 24599
rect 1676 24556 1728 24565
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 25228 24395 25280 24404
rect 25228 24361 25237 24395
rect 25237 24361 25271 24395
rect 25271 24361 25280 24395
rect 25228 24352 25280 24361
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 24952 24148 25004 24200
rect 33416 24055 33468 24064
rect 33416 24021 33425 24055
rect 33425 24021 33459 24055
rect 33459 24021 33468 24055
rect 33416 24012 33468 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 38016 23715 38068 23724
rect 38016 23681 38025 23715
rect 38025 23681 38059 23715
rect 38059 23681 38068 23715
rect 38016 23672 38068 23681
rect 38200 23511 38252 23520
rect 38200 23477 38209 23511
rect 38209 23477 38243 23511
rect 38243 23477 38252 23511
rect 38200 23468 38252 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1860 23264 1912 23316
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 38016 22720 38068 22772
rect 1768 22584 1820 22636
rect 37280 22584 37332 22636
rect 1676 22491 1728 22500
rect 1676 22457 1685 22491
rect 1685 22457 1719 22491
rect 1719 22457 1728 22491
rect 1676 22448 1728 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6828 21836 6880 21888
rect 9864 21836 9916 21888
rect 37280 21836 37332 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21496 1636 21548
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 1860 21403 1912 21412
rect 1860 21369 1869 21403
rect 1869 21369 1903 21403
rect 1903 21369 1912 21403
rect 1860 21360 1912 21369
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 38108 21088 38160 21140
rect 38108 20884 38160 20936
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1860 20408 1912 20460
rect 20260 20247 20312 20256
rect 20260 20213 20269 20247
rect 20269 20213 20303 20247
rect 20303 20213 20312 20247
rect 20260 20204 20312 20213
rect 33416 20204 33468 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 27896 20043 27948 20052
rect 27896 20009 27905 20043
rect 27905 20009 27939 20043
rect 27939 20009 27948 20043
rect 27896 20000 27948 20009
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 29276 19728 29328 19780
rect 38108 19703 38160 19712
rect 38108 19669 38117 19703
rect 38117 19669 38151 19703
rect 38151 19669 38160 19703
rect 38108 19660 38160 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1952 19320 2004 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 26148 18955 26200 18964
rect 26148 18921 26157 18955
rect 26157 18921 26191 18955
rect 26191 18921 26200 18955
rect 26148 18912 26200 18921
rect 25688 18751 25740 18760
rect 25688 18717 25697 18751
rect 25697 18717 25731 18751
rect 25731 18717 25740 18751
rect 25688 18708 25740 18717
rect 26148 18708 26200 18760
rect 38108 18708 38160 18760
rect 25596 18615 25648 18624
rect 25596 18581 25605 18615
rect 25605 18581 25639 18615
rect 25639 18581 25648 18615
rect 25596 18572 25648 18581
rect 33048 18615 33100 18624
rect 33048 18581 33057 18615
rect 33057 18581 33091 18615
rect 33091 18581 33100 18615
rect 33048 18572 33100 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 19432 18300 19484 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 19340 18232 19392 18284
rect 19340 18096 19392 18148
rect 24860 18207 24912 18216
rect 24860 18173 24869 18207
rect 24869 18173 24903 18207
rect 24903 18173 24912 18207
rect 24860 18164 24912 18173
rect 33048 18164 33100 18216
rect 30104 18096 30156 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 25136 18028 25188 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19248 17824 19300 17876
rect 21640 17867 21692 17876
rect 21640 17833 21649 17867
rect 21649 17833 21683 17867
rect 21683 17833 21692 17867
rect 21640 17824 21692 17833
rect 25688 17867 25740 17876
rect 25688 17833 25697 17867
rect 25697 17833 25731 17867
rect 25731 17833 25740 17867
rect 25688 17824 25740 17833
rect 23940 17756 23992 17808
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 22100 17688 22152 17740
rect 19524 17620 19576 17672
rect 23204 17620 23256 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 18144 17484 18196 17536
rect 23664 17552 23716 17604
rect 23112 17484 23164 17536
rect 25136 17484 25188 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3424 17280 3476 17332
rect 23112 17280 23164 17332
rect 18604 17255 18656 17264
rect 18604 17221 18613 17255
rect 18613 17221 18647 17255
rect 18647 17221 18656 17255
rect 18604 17212 18656 17221
rect 19248 17212 19300 17264
rect 22284 17212 22336 17264
rect 23940 17255 23992 17264
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 17316 17144 17368 17196
rect 21640 17144 21692 17196
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 15476 17076 15528 17128
rect 20812 17076 20864 17128
rect 22100 17119 22152 17128
rect 22100 17085 22109 17119
rect 22109 17085 22143 17119
rect 22143 17085 22152 17119
rect 22100 17076 22152 17085
rect 23664 17119 23716 17128
rect 18144 17051 18196 17060
rect 18144 17017 18153 17051
rect 18153 17017 18187 17051
rect 18187 17017 18196 17051
rect 18144 17008 18196 17017
rect 21732 17008 21784 17060
rect 23664 17085 23673 17119
rect 23673 17085 23707 17119
rect 23707 17085 23716 17119
rect 23664 17076 23716 17085
rect 24952 17280 25004 17332
rect 25872 17076 25924 17128
rect 23112 17008 23164 17060
rect 32956 17076 33008 17128
rect 15384 16940 15436 16992
rect 16028 16940 16080 16992
rect 16580 16940 16632 16992
rect 19248 16940 19300 16992
rect 21456 16940 21508 16992
rect 22376 16940 22428 16992
rect 24584 16983 24636 16992
rect 24584 16949 24593 16983
rect 24593 16949 24627 16983
rect 24627 16949 24636 16983
rect 24584 16940 24636 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16736 2096 16788
rect 14280 16736 14332 16788
rect 17592 16736 17644 16788
rect 19432 16736 19484 16788
rect 24952 16736 25004 16788
rect 23664 16668 23716 16720
rect 14832 16643 14884 16652
rect 14832 16609 14841 16643
rect 14841 16609 14875 16643
rect 14875 16609 14884 16643
rect 14832 16600 14884 16609
rect 15568 16600 15620 16652
rect 16212 16600 16264 16652
rect 17316 16532 17368 16584
rect 22100 16600 22152 16652
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 25136 16600 25188 16652
rect 13636 16464 13688 16516
rect 16120 16507 16172 16516
rect 16120 16473 16129 16507
rect 16129 16473 16163 16507
rect 16163 16473 16172 16507
rect 16120 16464 16172 16473
rect 16580 16464 16632 16516
rect 16764 16507 16816 16516
rect 16764 16473 16773 16507
rect 16773 16473 16807 16507
rect 16807 16473 16816 16507
rect 16764 16464 16816 16473
rect 10876 16396 10928 16448
rect 18420 16464 18472 16516
rect 21272 16464 21324 16516
rect 21732 16507 21784 16516
rect 21732 16473 21741 16507
rect 21741 16473 21775 16507
rect 21775 16473 21784 16507
rect 21732 16464 21784 16473
rect 21916 16464 21968 16516
rect 24952 16464 25004 16516
rect 25228 16507 25280 16516
rect 25228 16473 25237 16507
rect 25237 16473 25271 16507
rect 25271 16473 25280 16507
rect 25228 16464 25280 16473
rect 17224 16396 17276 16448
rect 22192 16396 22244 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 16120 16192 16172 16244
rect 4068 16056 4120 16108
rect 10692 15988 10744 16040
rect 14648 16124 14700 16176
rect 15752 16167 15804 16176
rect 15752 16133 15761 16167
rect 15761 16133 15795 16167
rect 15795 16133 15804 16167
rect 15752 16124 15804 16133
rect 13820 15988 13872 16040
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 16396 15988 16448 16040
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 15108 15920 15160 15972
rect 19432 16124 19484 16176
rect 20076 16124 20128 16176
rect 23296 16192 23348 16244
rect 24768 16192 24820 16244
rect 24860 16192 24912 16244
rect 32956 16235 33008 16244
rect 32956 16201 32965 16235
rect 32965 16201 32999 16235
rect 32999 16201 33008 16235
rect 32956 16192 33008 16201
rect 16580 16056 16632 16108
rect 18420 16099 18472 16108
rect 16856 15988 16908 16040
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 19984 16056 20036 16108
rect 20260 16056 20312 16108
rect 22100 16056 22152 16108
rect 24492 16099 24544 16108
rect 24492 16065 24501 16099
rect 24501 16065 24535 16099
rect 24535 16065 24544 16099
rect 24492 16056 24544 16065
rect 24768 16056 24820 16108
rect 37832 16056 37884 16108
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 19524 15988 19576 16040
rect 20720 16031 20772 16040
rect 20720 15997 20729 16031
rect 20729 15997 20763 16031
rect 20763 15997 20772 16031
rect 20720 15988 20772 15997
rect 23204 16031 23256 16040
rect 23204 15997 23213 16031
rect 23213 15997 23247 16031
rect 23247 15997 23256 16031
rect 23204 15988 23256 15997
rect 38292 16031 38344 16040
rect 38292 15997 38301 16031
rect 38301 15997 38335 16031
rect 38335 15997 38344 16031
rect 38292 15988 38344 15997
rect 16304 15852 16356 15904
rect 18236 15852 18288 15904
rect 19616 15852 19668 15904
rect 22008 15852 22060 15904
rect 23940 15895 23992 15904
rect 23940 15861 23949 15895
rect 23949 15861 23983 15895
rect 23983 15861 23992 15895
rect 23940 15852 23992 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 14740 15648 14792 15700
rect 16580 15648 16632 15700
rect 19524 15648 19576 15700
rect 20812 15648 20864 15700
rect 21824 15648 21876 15700
rect 22008 15691 22060 15700
rect 22008 15657 22017 15691
rect 22017 15657 22051 15691
rect 22051 15657 22060 15691
rect 22008 15648 22060 15657
rect 23848 15648 23900 15700
rect 38016 15648 38068 15700
rect 38292 15691 38344 15700
rect 38292 15657 38301 15691
rect 38301 15657 38335 15691
rect 38335 15657 38344 15691
rect 38292 15648 38344 15657
rect 15016 15580 15068 15632
rect 13912 15512 13964 15564
rect 15108 15512 15160 15564
rect 2412 15444 2464 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 13820 15444 13872 15496
rect 14648 15444 14700 15496
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 15660 15512 15712 15564
rect 16764 15580 16816 15632
rect 17684 15580 17736 15632
rect 18328 15512 18380 15564
rect 19432 15580 19484 15632
rect 14740 15444 14792 15453
rect 17316 15444 17368 15496
rect 23480 15580 23532 15632
rect 23940 15580 23992 15632
rect 35440 15580 35492 15632
rect 16028 15419 16080 15428
rect 16028 15385 16037 15419
rect 16037 15385 16071 15419
rect 16071 15385 16080 15419
rect 16028 15376 16080 15385
rect 18328 15419 18380 15428
rect 18328 15385 18337 15419
rect 18337 15385 18371 15419
rect 18371 15385 18380 15419
rect 18328 15376 18380 15385
rect 19616 15419 19668 15428
rect 19616 15385 19625 15419
rect 19625 15385 19659 15419
rect 19659 15385 19668 15419
rect 19616 15376 19668 15385
rect 21272 15376 21324 15428
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 14556 15308 14608 15360
rect 15936 15308 15988 15360
rect 16856 15308 16908 15360
rect 21456 15444 21508 15496
rect 25320 15512 25372 15564
rect 25596 15512 25648 15564
rect 22744 15444 22796 15496
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 25136 15444 25188 15496
rect 29828 15444 29880 15496
rect 24676 15376 24728 15428
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 15476 15104 15528 15156
rect 15752 15104 15804 15156
rect 16488 15104 16540 15156
rect 19340 15147 19392 15156
rect 2136 14968 2188 15020
rect 7380 14968 7432 15020
rect 11704 14968 11756 15020
rect 14372 15036 14424 15088
rect 13728 14968 13780 15020
rect 14556 14968 14608 15020
rect 15384 15036 15436 15088
rect 16948 15036 17000 15088
rect 17224 15036 17276 15088
rect 18236 15079 18288 15088
rect 18236 15045 18245 15079
rect 18245 15045 18279 15079
rect 18279 15045 18288 15079
rect 18236 15036 18288 15045
rect 19340 15113 19349 15147
rect 19349 15113 19383 15147
rect 19383 15113 19392 15147
rect 19340 15104 19392 15113
rect 20720 15104 20772 15156
rect 21548 15104 21600 15156
rect 22008 15104 22060 15156
rect 23480 15104 23532 15156
rect 24768 15104 24820 15156
rect 25044 15104 25096 15156
rect 20812 15079 20864 15088
rect 20812 15045 20821 15079
rect 20821 15045 20855 15079
rect 20855 15045 20864 15079
rect 20812 15036 20864 15045
rect 22284 15036 22336 15088
rect 24124 15079 24176 15088
rect 24124 15045 24133 15079
rect 24133 15045 24167 15079
rect 24167 15045 24176 15079
rect 24124 15036 24176 15045
rect 10784 14900 10836 14952
rect 15292 14968 15344 15020
rect 16028 14968 16080 15020
rect 16212 14968 16264 15020
rect 19156 14968 19208 15020
rect 19892 15011 19944 15020
rect 17040 14900 17092 14952
rect 1860 14832 1912 14884
rect 15200 14832 15252 14884
rect 16396 14832 16448 14884
rect 17500 14875 17552 14884
rect 17500 14841 17509 14875
rect 17509 14841 17543 14875
rect 17543 14841 17552 14875
rect 17500 14832 17552 14841
rect 18420 14900 18472 14952
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 18512 14832 18564 14884
rect 11244 14764 11296 14816
rect 13544 14764 13596 14816
rect 14004 14764 14056 14816
rect 15108 14764 15160 14816
rect 16304 14764 16356 14816
rect 19064 14764 19116 14816
rect 22744 14900 22796 14952
rect 23112 14943 23164 14952
rect 23112 14909 23121 14943
rect 23121 14909 23155 14943
rect 23155 14909 23164 14943
rect 23112 14900 23164 14909
rect 23204 14900 23256 14952
rect 25228 14900 25280 14952
rect 21548 14832 21600 14884
rect 27160 14832 27212 14884
rect 24492 14764 24544 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 11704 14492 11756 14544
rect 12256 14492 12308 14544
rect 14188 14560 14240 14612
rect 14740 14560 14792 14612
rect 15660 14560 15712 14612
rect 17868 14560 17920 14612
rect 18328 14560 18380 14612
rect 18512 14560 18564 14612
rect 14372 14492 14424 14544
rect 15752 14492 15804 14544
rect 16488 14492 16540 14544
rect 15016 14467 15068 14476
rect 12164 14356 12216 14408
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 17500 14492 17552 14544
rect 17684 14467 17736 14476
rect 17684 14433 17693 14467
rect 17693 14433 17727 14467
rect 17727 14433 17736 14467
rect 17684 14424 17736 14433
rect 19892 14424 19944 14476
rect 20260 14424 20312 14476
rect 21548 14492 21600 14544
rect 20812 14399 20864 14408
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 12532 14288 12584 14340
rect 14464 14331 14516 14340
rect 14464 14297 14473 14331
rect 14473 14297 14507 14331
rect 14507 14297 14516 14331
rect 14464 14288 14516 14297
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 13360 14220 13412 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 14924 14220 14976 14272
rect 16580 14288 16632 14340
rect 15936 14220 15988 14272
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 19432 14331 19484 14340
rect 19432 14297 19441 14331
rect 19441 14297 19475 14331
rect 19475 14297 19484 14331
rect 19432 14288 19484 14297
rect 19984 14331 20036 14340
rect 19984 14297 19993 14331
rect 19993 14297 20027 14331
rect 20027 14297 20036 14331
rect 19984 14288 20036 14297
rect 18788 14220 18840 14272
rect 21548 14288 21600 14340
rect 23204 14467 23256 14476
rect 23204 14433 23213 14467
rect 23213 14433 23247 14467
rect 23247 14433 23256 14467
rect 23204 14424 23256 14433
rect 31300 14492 31352 14544
rect 24676 14467 24728 14476
rect 24676 14433 24685 14467
rect 24685 14433 24719 14467
rect 24719 14433 24728 14467
rect 25228 14467 25280 14476
rect 24676 14424 24728 14433
rect 25228 14433 25237 14467
rect 25237 14433 25271 14467
rect 25271 14433 25280 14467
rect 25228 14424 25280 14433
rect 26332 14356 26384 14408
rect 38016 14399 38068 14408
rect 22376 14331 22428 14340
rect 22376 14297 22385 14331
rect 22385 14297 22419 14331
rect 22419 14297 22428 14331
rect 22376 14288 22428 14297
rect 23020 14331 23072 14340
rect 23020 14297 23029 14331
rect 23029 14297 23063 14331
rect 23063 14297 23072 14331
rect 23020 14288 23072 14297
rect 23388 14220 23440 14272
rect 25964 14263 26016 14272
rect 25964 14229 25973 14263
rect 25973 14229 26007 14263
rect 26007 14229 26016 14263
rect 25964 14220 26016 14229
rect 26608 14263 26660 14272
rect 26608 14229 26617 14263
rect 26617 14229 26651 14263
rect 26651 14229 26660 14263
rect 26608 14220 26660 14229
rect 38016 14365 38025 14399
rect 38025 14365 38059 14399
rect 38059 14365 38068 14399
rect 38016 14356 38068 14365
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 34244 14220 34296 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 10876 14016 10928 14068
rect 14464 14016 14516 14068
rect 15568 14016 15620 14068
rect 11060 13948 11112 14000
rect 13544 13948 13596 14000
rect 15200 13948 15252 14000
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 16488 13948 16540 14000
rect 18604 14016 18656 14068
rect 17684 13948 17736 14000
rect 19340 13948 19392 14000
rect 21456 13948 21508 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 12164 13880 12216 13932
rect 12256 13923 12308 13932
rect 12256 13889 12265 13923
rect 12265 13889 12299 13923
rect 12299 13889 12308 13923
rect 12256 13880 12308 13889
rect 12532 13812 12584 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13912 13880 13964 13932
rect 18052 13923 18104 13932
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 20260 13880 20312 13932
rect 13360 13812 13412 13821
rect 13636 13812 13688 13864
rect 15660 13855 15712 13864
rect 7748 13744 7800 13796
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 15476 13744 15528 13796
rect 16304 13812 16356 13864
rect 17040 13812 17092 13864
rect 19432 13812 19484 13864
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 22192 13991 22244 14000
rect 22192 13957 22201 13991
rect 22201 13957 22235 13991
rect 22235 13957 22244 13991
rect 22192 13948 22244 13957
rect 22376 13948 22428 14000
rect 23112 13991 23164 14000
rect 23112 13957 23121 13991
rect 23121 13957 23155 13991
rect 23155 13957 23164 13991
rect 37280 14016 37332 14068
rect 38292 14059 38344 14068
rect 38292 14025 38301 14059
rect 38301 14025 38335 14059
rect 38335 14025 38344 14059
rect 38292 14016 38344 14025
rect 23112 13948 23164 13957
rect 25044 13948 25096 14000
rect 27528 13948 27580 14000
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 28816 13812 28868 13864
rect 34244 13812 34296 13864
rect 35808 13812 35860 13864
rect 10508 13676 10560 13728
rect 12900 13676 12952 13728
rect 13820 13676 13872 13728
rect 15200 13676 15252 13728
rect 15292 13676 15344 13728
rect 21548 13744 21600 13796
rect 24308 13744 24360 13796
rect 21180 13676 21232 13728
rect 22192 13676 22244 13728
rect 24216 13676 24268 13728
rect 27988 13676 28040 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 11060 13515 11112 13524
rect 11060 13481 11069 13515
rect 11069 13481 11103 13515
rect 11103 13481 11112 13515
rect 11060 13472 11112 13481
rect 14924 13472 14976 13524
rect 15476 13472 15528 13524
rect 1952 13404 2004 13456
rect 9864 13404 9916 13456
rect 13544 13404 13596 13456
rect 13728 13404 13780 13456
rect 20628 13472 20680 13524
rect 23020 13472 23072 13524
rect 26424 13472 26476 13524
rect 10324 13268 10376 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 21732 13404 21784 13456
rect 23848 13404 23900 13456
rect 15292 13336 15344 13388
rect 16672 13336 16724 13388
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 19248 13336 19300 13388
rect 20168 13336 20220 13388
rect 23204 13336 23256 13388
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 12900 13268 12952 13277
rect 13820 13268 13872 13320
rect 14280 13311 14332 13320
rect 9312 13200 9364 13252
rect 10232 13200 10284 13252
rect 10692 13200 10744 13252
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 16028 13268 16080 13320
rect 16304 13268 16356 13320
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 24400 13404 24452 13456
rect 25136 13336 25188 13388
rect 26148 13336 26200 13388
rect 31208 13404 31260 13456
rect 24492 13268 24544 13320
rect 15108 13243 15160 13252
rect 15108 13209 15117 13243
rect 15117 13209 15151 13243
rect 15151 13209 15160 13243
rect 15660 13243 15712 13252
rect 15108 13200 15160 13209
rect 15660 13209 15669 13243
rect 15669 13209 15703 13243
rect 15703 13209 15712 13243
rect 15660 13200 15712 13209
rect 17224 13243 17276 13252
rect 17224 13209 17233 13243
rect 17233 13209 17267 13243
rect 17267 13209 17276 13243
rect 17224 13200 17276 13209
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 2504 13175 2556 13184
rect 2504 13141 2513 13175
rect 2513 13141 2547 13175
rect 2547 13141 2556 13175
rect 2504 13132 2556 13141
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 15200 13132 15252 13184
rect 18420 13200 18472 13252
rect 17776 13132 17828 13184
rect 20720 13243 20772 13252
rect 20720 13209 20729 13243
rect 20729 13209 20763 13243
rect 20763 13209 20772 13243
rect 20720 13200 20772 13209
rect 21364 13200 21416 13252
rect 22284 13200 22336 13252
rect 24584 13243 24636 13252
rect 21732 13132 21784 13184
rect 24584 13209 24593 13243
rect 24593 13209 24627 13243
rect 24627 13209 24636 13243
rect 24584 13200 24636 13209
rect 25136 13243 25188 13252
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 26056 13200 26108 13252
rect 27344 13200 27396 13252
rect 24400 13132 24452 13184
rect 24492 13132 24544 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2136 12928 2188 12980
rect 2504 12860 2556 12912
rect 7748 12903 7800 12912
rect 5540 12792 5592 12844
rect 7748 12869 7757 12903
rect 7757 12869 7791 12903
rect 7791 12869 7800 12903
rect 7748 12860 7800 12869
rect 10416 12860 10468 12912
rect 14004 12903 14056 12912
rect 14004 12869 14013 12903
rect 14013 12869 14047 12903
rect 14047 12869 14056 12903
rect 14004 12860 14056 12869
rect 14372 12928 14424 12980
rect 13544 12792 13596 12844
rect 12256 12724 12308 12776
rect 13912 12767 13964 12776
rect 12532 12699 12584 12708
rect 12532 12665 12541 12699
rect 12541 12665 12575 12699
rect 12575 12665 12584 12699
rect 12532 12656 12584 12665
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 14280 12724 14332 12776
rect 15384 12860 15436 12912
rect 16028 12860 16080 12912
rect 17684 12860 17736 12912
rect 18604 12860 18656 12912
rect 18788 12903 18840 12912
rect 18788 12869 18797 12903
rect 18797 12869 18831 12903
rect 18831 12869 18840 12903
rect 18788 12860 18840 12869
rect 20076 12903 20128 12912
rect 20076 12869 20085 12903
rect 20085 12869 20119 12903
rect 20119 12869 20128 12903
rect 20076 12860 20128 12869
rect 20168 12903 20220 12912
rect 20168 12869 20177 12903
rect 20177 12869 20211 12903
rect 20211 12869 20220 12903
rect 20168 12860 20220 12869
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 15660 12724 15712 12776
rect 14096 12656 14148 12708
rect 14740 12656 14792 12708
rect 16764 12724 16816 12776
rect 17040 12724 17092 12776
rect 20168 12724 20220 12776
rect 22284 12860 22336 12912
rect 21456 12792 21508 12844
rect 24676 12928 24728 12980
rect 25136 12928 25188 12980
rect 27528 12928 27580 12980
rect 28448 12928 28500 12980
rect 28816 12971 28868 12980
rect 28816 12937 28825 12971
rect 28825 12937 28859 12971
rect 28859 12937 28868 12971
rect 28816 12928 28868 12937
rect 26608 12860 26660 12912
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 21824 12724 21876 12776
rect 25964 12792 26016 12844
rect 23756 12724 23808 12776
rect 23940 12767 23992 12776
rect 23940 12733 23949 12767
rect 23949 12733 23983 12767
rect 23983 12733 23992 12767
rect 23940 12724 23992 12733
rect 21180 12699 21232 12708
rect 21180 12665 21189 12699
rect 21189 12665 21223 12699
rect 21223 12665 21232 12699
rect 21180 12656 21232 12665
rect 25688 12724 25740 12776
rect 26792 12792 26844 12844
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 38016 12860 38068 12912
rect 26056 12699 26108 12708
rect 26056 12665 26065 12699
rect 26065 12665 26099 12699
rect 26099 12665 26108 12699
rect 26056 12656 26108 12665
rect 27068 12724 27120 12776
rect 34152 12724 34204 12776
rect 38292 12767 38344 12776
rect 38292 12733 38301 12767
rect 38301 12733 38335 12767
rect 38335 12733 38344 12767
rect 38292 12724 38344 12733
rect 27528 12656 27580 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 13176 12588 13228 12640
rect 24676 12588 24728 12640
rect 30104 12631 30156 12640
rect 30104 12597 30113 12631
rect 30113 12597 30147 12631
rect 30147 12597 30156 12631
rect 30104 12588 30156 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5540 12384 5592 12436
rect 15752 12384 15804 12436
rect 15844 12384 15896 12436
rect 13452 12316 13504 12368
rect 19340 12384 19392 12436
rect 20720 12384 20772 12436
rect 23756 12427 23808 12436
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 12624 12248 12676 12300
rect 12716 12291 12768 12300
rect 12716 12257 12725 12291
rect 12725 12257 12759 12291
rect 12759 12257 12768 12291
rect 12716 12248 12768 12257
rect 14188 12248 14240 12300
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 17684 12248 17736 12300
rect 20996 12316 21048 12368
rect 20904 12248 20956 12300
rect 10140 12180 10192 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 9772 12155 9824 12164
rect 9772 12121 9781 12155
rect 9781 12121 9815 12155
rect 9815 12121 9824 12155
rect 9772 12112 9824 12121
rect 9864 12112 9916 12164
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 13452 12180 13504 12232
rect 14004 12180 14056 12232
rect 14280 12180 14332 12232
rect 14556 12180 14608 12232
rect 18420 12180 18472 12232
rect 20352 12180 20404 12232
rect 20812 12180 20864 12232
rect 12072 12112 12124 12164
rect 12394 12112 12446 12164
rect 10968 12087 11020 12096
rect 8576 12044 8628 12053
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 14648 12044 14700 12096
rect 15660 12112 15712 12164
rect 16488 12155 16540 12164
rect 16488 12121 16497 12155
rect 16497 12121 16531 12155
rect 16531 12121 16540 12155
rect 16488 12112 16540 12121
rect 18236 12155 18288 12164
rect 18236 12121 18245 12155
rect 18245 12121 18279 12155
rect 18279 12121 18288 12155
rect 18236 12112 18288 12121
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 21640 12155 21692 12164
rect 21640 12121 21649 12155
rect 21649 12121 21683 12155
rect 21683 12121 21692 12155
rect 21640 12112 21692 12121
rect 21824 12112 21876 12164
rect 18604 12044 18656 12096
rect 24308 12316 24360 12368
rect 22652 12291 22704 12300
rect 22652 12257 22661 12291
rect 22661 12257 22695 12291
rect 22695 12257 22704 12291
rect 22652 12248 22704 12257
rect 25688 12384 25740 12436
rect 26056 12427 26108 12436
rect 26056 12393 26065 12427
rect 26065 12393 26099 12427
rect 26099 12393 26108 12427
rect 26056 12384 26108 12393
rect 27528 12384 27580 12436
rect 25320 12316 25372 12368
rect 26424 12316 26476 12368
rect 26792 12316 26844 12368
rect 28172 12316 28224 12368
rect 30104 12316 30156 12368
rect 37464 12316 37516 12368
rect 38292 12359 38344 12368
rect 38292 12325 38301 12359
rect 38301 12325 38335 12359
rect 38335 12325 38344 12359
rect 38292 12316 38344 12325
rect 24032 12180 24084 12232
rect 26608 12180 26660 12232
rect 27436 12248 27488 12300
rect 26884 12180 26936 12232
rect 27068 12223 27120 12232
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 27528 12223 27580 12232
rect 27528 12189 27537 12223
rect 27537 12189 27571 12223
rect 27571 12189 27580 12223
rect 27528 12180 27580 12189
rect 28080 12180 28132 12232
rect 29000 12223 29052 12232
rect 29000 12189 29009 12223
rect 29009 12189 29043 12223
rect 29043 12189 29052 12223
rect 29000 12180 29052 12189
rect 24308 12112 24360 12164
rect 25412 12044 25464 12096
rect 25504 12044 25556 12096
rect 28356 12044 28408 12096
rect 29276 12044 29328 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 10968 11840 11020 11892
rect 15568 11883 15620 11892
rect 8392 11704 8444 11756
rect 9220 11704 9272 11756
rect 9956 11772 10008 11824
rect 14096 11815 14148 11824
rect 14096 11781 14105 11815
rect 14105 11781 14139 11815
rect 14139 11781 14148 11815
rect 14096 11772 14148 11781
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 17684 11840 17736 11892
rect 14740 11815 14792 11824
rect 14740 11781 14749 11815
rect 14749 11781 14783 11815
rect 14783 11781 14792 11815
rect 14740 11772 14792 11781
rect 15844 11772 15896 11824
rect 17040 11815 17092 11824
rect 10508 11704 10560 11756
rect 10784 11636 10836 11688
rect 11152 11704 11204 11756
rect 12256 11704 12308 11756
rect 12624 11704 12676 11756
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 15936 11704 15988 11756
rect 17040 11781 17049 11815
rect 17049 11781 17083 11815
rect 17083 11781 17092 11815
rect 17040 11772 17092 11781
rect 17132 11772 17184 11824
rect 17868 11772 17920 11824
rect 21180 11840 21232 11892
rect 23940 11883 23992 11892
rect 21088 11772 21140 11824
rect 21732 11772 21784 11824
rect 23940 11849 23949 11883
rect 23949 11849 23983 11883
rect 23983 11849 23992 11883
rect 23940 11840 23992 11849
rect 26056 11840 26108 11892
rect 27252 11883 27304 11892
rect 27252 11849 27261 11883
rect 27261 11849 27295 11883
rect 27295 11849 27304 11883
rect 27252 11840 27304 11849
rect 27436 11840 27488 11892
rect 30380 11840 30432 11892
rect 33232 11840 33284 11892
rect 34152 11840 34204 11892
rect 22560 11772 22612 11824
rect 24768 11815 24820 11824
rect 24768 11781 24777 11815
rect 24777 11781 24811 11815
rect 24811 11781 24820 11815
rect 24768 11772 24820 11781
rect 16396 11704 16448 11756
rect 23848 11747 23900 11756
rect 16672 11636 16724 11688
rect 17868 11679 17920 11688
rect 13728 11568 13780 11620
rect 14188 11568 14240 11620
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 20076 11679 20128 11688
rect 20076 11645 20085 11679
rect 20085 11645 20119 11679
rect 20119 11645 20128 11679
rect 20076 11636 20128 11645
rect 12164 11500 12216 11552
rect 16028 11500 16080 11552
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 26332 11704 26384 11756
rect 30932 11772 30984 11824
rect 28632 11747 28684 11756
rect 22468 11636 22520 11688
rect 25320 11679 25372 11688
rect 25320 11645 25329 11679
rect 25329 11645 25363 11679
rect 25363 11645 25372 11679
rect 25320 11636 25372 11645
rect 25872 11636 25924 11688
rect 22744 11568 22796 11620
rect 23848 11568 23900 11620
rect 27436 11636 27488 11688
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 35900 11636 35952 11688
rect 27252 11568 27304 11620
rect 21640 11500 21692 11552
rect 26240 11500 26292 11552
rect 27436 11500 27488 11552
rect 27988 11568 28040 11620
rect 30380 11611 30432 11620
rect 30380 11577 30389 11611
rect 30389 11577 30423 11611
rect 30423 11577 30432 11611
rect 30380 11568 30432 11577
rect 29736 11543 29788 11552
rect 29736 11509 29745 11543
rect 29745 11509 29779 11543
rect 29779 11509 29788 11543
rect 29736 11500 29788 11509
rect 30932 11543 30984 11552
rect 30932 11509 30941 11543
rect 30941 11509 30975 11543
rect 30975 11509 30984 11543
rect 30932 11500 30984 11509
rect 33508 11500 33560 11552
rect 38292 11543 38344 11552
rect 38292 11509 38301 11543
rect 38301 11509 38335 11543
rect 38335 11509 38344 11543
rect 38292 11500 38344 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 12348 11296 12400 11348
rect 11060 11228 11112 11280
rect 15384 11296 15436 11348
rect 15568 11296 15620 11348
rect 15752 11296 15804 11348
rect 16028 11296 16080 11348
rect 16212 11296 16264 11348
rect 16488 11296 16540 11348
rect 14648 11228 14700 11280
rect 9864 11160 9916 11212
rect 12164 11160 12216 11212
rect 12808 11160 12860 11212
rect 8392 11092 8444 11144
rect 11152 11092 11204 11144
rect 11612 11092 11664 11144
rect 12624 11092 12676 11144
rect 12992 11092 13044 11144
rect 1860 10956 1912 11008
rect 11520 11024 11572 11076
rect 9588 10956 9640 11008
rect 11152 10956 11204 11008
rect 12348 10956 12400 11008
rect 13820 11024 13872 11076
rect 14280 11092 14332 11144
rect 16396 11160 16448 11212
rect 16948 11160 17000 11212
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 16028 11092 16080 11144
rect 15752 11067 15804 11076
rect 15752 11033 15761 11067
rect 15761 11033 15795 11067
rect 15795 11033 15804 11067
rect 15752 11024 15804 11033
rect 15844 11067 15896 11076
rect 15844 11033 15853 11067
rect 15853 11033 15887 11067
rect 15887 11033 15896 11067
rect 15844 11024 15896 11033
rect 18604 11228 18656 11280
rect 20076 11296 20128 11348
rect 21180 11296 21232 11348
rect 23848 11296 23900 11348
rect 24124 11296 24176 11348
rect 24492 11296 24544 11348
rect 24676 11296 24728 11348
rect 25412 11296 25464 11348
rect 22192 11228 22244 11280
rect 19064 11160 19116 11212
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 21272 11160 21324 11212
rect 21732 11160 21784 11212
rect 22468 11160 22520 11212
rect 23112 11160 23164 11212
rect 23756 11160 23808 11212
rect 24492 11160 24544 11212
rect 29736 11296 29788 11348
rect 28080 11228 28132 11280
rect 29644 11228 29696 11280
rect 29828 11228 29880 11280
rect 30472 11228 30524 11280
rect 19432 11092 19484 11144
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 17592 11024 17644 11076
rect 20628 11024 20680 11076
rect 13176 10956 13228 11008
rect 16028 10956 16080 11008
rect 16672 10956 16724 11008
rect 22468 11024 22520 11076
rect 23572 11092 23624 11144
rect 31024 11160 31076 11212
rect 25780 11092 25832 11144
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 26516 11135 26568 11144
rect 25872 11092 25924 11101
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27988 11092 28040 11144
rect 29828 11092 29880 11144
rect 30012 11092 30064 11144
rect 30656 11092 30708 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 26976 11024 27028 11076
rect 28264 11067 28316 11076
rect 21824 10956 21876 11008
rect 25136 10956 25188 11008
rect 25228 10999 25280 11008
rect 25228 10965 25237 10999
rect 25237 10965 25271 10999
rect 25271 10965 25280 10999
rect 25228 10956 25280 10965
rect 25504 10956 25556 11008
rect 27988 10956 28040 11008
rect 28264 11033 28273 11067
rect 28273 11033 28307 11067
rect 28307 11033 28316 11067
rect 28264 11024 28316 11033
rect 28540 10956 28592 11008
rect 31392 11024 31444 11076
rect 29644 10956 29696 11008
rect 31300 10956 31352 11008
rect 37924 10956 37976 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 10876 10752 10928 10804
rect 11152 10684 11204 10736
rect 11244 10684 11296 10736
rect 12716 10727 12768 10736
rect 12716 10693 12725 10727
rect 12725 10693 12759 10727
rect 12759 10693 12768 10727
rect 12716 10684 12768 10693
rect 12900 10684 12952 10736
rect 13452 10684 13504 10736
rect 16580 10684 16632 10736
rect 17408 10684 17460 10736
rect 20076 10752 20128 10804
rect 21548 10752 21600 10804
rect 23572 10795 23624 10804
rect 23572 10761 23581 10795
rect 23581 10761 23615 10795
rect 23615 10761 23624 10795
rect 24768 10795 24820 10804
rect 23572 10752 23624 10761
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 25228 10752 25280 10804
rect 28264 10752 28316 10804
rect 28632 10752 28684 10804
rect 19064 10684 19116 10736
rect 9404 10616 9456 10668
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 10968 10659 11020 10668
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 16764 10616 16816 10668
rect 10876 10548 10928 10600
rect 12164 10548 12216 10600
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 8668 10412 8720 10464
rect 10968 10480 11020 10532
rect 13912 10480 13964 10532
rect 16948 10548 17000 10600
rect 18328 10591 18380 10600
rect 15016 10523 15068 10532
rect 15016 10489 15025 10523
rect 15025 10489 15059 10523
rect 15059 10489 15068 10523
rect 15016 10480 15068 10489
rect 15844 10480 15896 10532
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 20076 10548 20128 10600
rect 22652 10684 22704 10736
rect 24860 10684 24912 10736
rect 25136 10684 25188 10736
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 21916 10616 21968 10668
rect 23204 10616 23256 10668
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 22744 10548 22796 10600
rect 24032 10591 24084 10600
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 24492 10616 24544 10668
rect 25504 10616 25556 10668
rect 25780 10616 25832 10668
rect 28080 10659 28132 10668
rect 25320 10548 25372 10600
rect 26424 10591 26476 10600
rect 20444 10480 20496 10532
rect 21824 10480 21876 10532
rect 21916 10480 21968 10532
rect 23940 10480 23992 10532
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 26608 10591 26660 10600
rect 26608 10557 26617 10591
rect 26617 10557 26651 10591
rect 26651 10557 26660 10591
rect 26608 10548 26660 10557
rect 28080 10625 28089 10659
rect 28089 10625 28123 10659
rect 28123 10625 28132 10659
rect 28080 10616 28132 10625
rect 28172 10616 28224 10668
rect 31392 10616 31444 10668
rect 38016 10616 38068 10668
rect 27068 10480 27120 10532
rect 12992 10412 13044 10464
rect 17408 10412 17460 10464
rect 18880 10412 18932 10464
rect 20260 10412 20312 10464
rect 26332 10412 26384 10464
rect 26792 10412 26844 10464
rect 27252 10412 27304 10464
rect 27344 10412 27396 10464
rect 30104 10455 30156 10464
rect 30104 10421 30113 10455
rect 30113 10421 30147 10455
rect 30147 10421 30156 10455
rect 30104 10412 30156 10421
rect 31392 10455 31444 10464
rect 31392 10421 31401 10455
rect 31401 10421 31435 10455
rect 31435 10421 31444 10455
rect 31392 10412 31444 10421
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 12808 10208 12860 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 19432 10208 19484 10260
rect 9588 10140 9640 10192
rect 10140 10072 10192 10124
rect 12532 10072 12584 10124
rect 16120 10140 16172 10192
rect 16672 10140 16724 10192
rect 18880 10183 18932 10192
rect 18880 10149 18889 10183
rect 18889 10149 18923 10183
rect 18923 10149 18932 10183
rect 18880 10140 18932 10149
rect 22100 10208 22152 10260
rect 24584 10208 24636 10260
rect 26424 10208 26476 10260
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13360 10004 13412 10056
rect 22744 10140 22796 10192
rect 22652 10072 22704 10124
rect 24768 10072 24820 10124
rect 26240 10140 26292 10192
rect 30104 10140 30156 10192
rect 26792 10072 26844 10124
rect 27160 10072 27212 10124
rect 28540 10115 28592 10124
rect 16304 10004 16356 10056
rect 11060 9936 11112 9988
rect 12164 9979 12216 9988
rect 12164 9945 12173 9979
rect 12173 9945 12207 9979
rect 12207 9945 12216 9979
rect 12164 9936 12216 9945
rect 12624 9936 12676 9988
rect 13912 9936 13964 9988
rect 14372 9936 14424 9988
rect 15108 9936 15160 9988
rect 15844 9936 15896 9988
rect 13820 9868 13872 9920
rect 18972 10004 19024 10056
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 19984 10004 20036 10056
rect 20444 10004 20496 10056
rect 19248 9936 19300 9988
rect 19340 9936 19392 9988
rect 19892 9936 19944 9988
rect 21272 9979 21324 9988
rect 21272 9945 21281 9979
rect 21281 9945 21315 9979
rect 21315 9945 21324 9979
rect 21272 9936 21324 9945
rect 18880 9868 18932 9920
rect 19432 9868 19484 9920
rect 19708 9868 19760 9920
rect 22192 9936 22244 9988
rect 26240 10004 26292 10056
rect 28540 10081 28549 10115
rect 28549 10081 28583 10115
rect 28583 10081 28592 10115
rect 28540 10072 28592 10081
rect 25688 9979 25740 9988
rect 25688 9945 25697 9979
rect 25697 9945 25731 9979
rect 25731 9945 25740 9979
rect 25688 9936 25740 9945
rect 26148 9936 26200 9988
rect 29828 10004 29880 10056
rect 30288 10004 30340 10056
rect 27068 9979 27120 9988
rect 27068 9945 27077 9979
rect 27077 9945 27111 9979
rect 27111 9945 27120 9979
rect 27068 9936 27120 9945
rect 27712 9868 27764 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 13084 9664 13136 9716
rect 16856 9664 16908 9716
rect 20076 9664 20128 9716
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 11244 9596 11296 9648
rect 11336 9596 11388 9648
rect 14188 9596 14240 9648
rect 14740 9596 14792 9648
rect 15200 9596 15252 9648
rect 21548 9664 21600 9716
rect 22192 9664 22244 9716
rect 8668 9528 8720 9580
rect 11888 9528 11940 9580
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 12348 9460 12400 9512
rect 9312 9435 9364 9444
rect 9312 9401 9321 9435
rect 9321 9401 9355 9435
rect 9355 9401 9364 9435
rect 9312 9392 9364 9401
rect 16212 9528 16264 9580
rect 16672 9528 16724 9580
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 13636 9460 13688 9512
rect 13728 9460 13780 9512
rect 13084 9392 13136 9444
rect 16304 9503 16356 9512
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 16764 9460 16816 9512
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 19616 9460 19668 9512
rect 20168 9460 20220 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 13912 9324 13964 9376
rect 17132 9392 17184 9444
rect 22192 9528 22244 9580
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 22100 9503 22152 9512
rect 22100 9469 22109 9503
rect 22109 9469 22143 9503
rect 22143 9469 22152 9503
rect 23480 9596 23532 9648
rect 24584 9664 24636 9716
rect 27252 9664 27304 9716
rect 24676 9596 24728 9648
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 27620 9596 27672 9648
rect 28356 9596 28408 9648
rect 25872 9528 25924 9580
rect 26884 9528 26936 9580
rect 27988 9528 28040 9580
rect 30472 9596 30524 9648
rect 30380 9571 30432 9580
rect 30380 9537 30389 9571
rect 30389 9537 30423 9571
rect 30423 9537 30432 9571
rect 30380 9528 30432 9537
rect 22100 9460 22152 9469
rect 23848 9503 23900 9512
rect 23848 9469 23857 9503
rect 23857 9469 23891 9503
rect 23891 9469 23900 9503
rect 23848 9460 23900 9469
rect 24952 9460 25004 9512
rect 26240 9460 26292 9512
rect 26424 9503 26476 9512
rect 26424 9469 26433 9503
rect 26433 9469 26467 9503
rect 26467 9469 26476 9503
rect 26424 9460 26476 9469
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 27620 9460 27672 9512
rect 27804 9503 27856 9512
rect 27804 9469 27813 9503
rect 27813 9469 27847 9503
rect 27847 9469 27856 9503
rect 27804 9460 27856 9469
rect 28448 9460 28500 9512
rect 29736 9503 29788 9512
rect 15384 9324 15436 9376
rect 15936 9324 15988 9376
rect 16948 9324 17000 9376
rect 18052 9324 18104 9376
rect 18604 9324 18656 9376
rect 21180 9324 21232 9376
rect 27344 9392 27396 9444
rect 24584 9324 24636 9376
rect 27712 9392 27764 9444
rect 29736 9469 29745 9503
rect 29745 9469 29779 9503
rect 29779 9469 29788 9503
rect 29736 9460 29788 9469
rect 27528 9324 27580 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 11336 9120 11388 9172
rect 12900 9120 12952 9172
rect 15200 9120 15252 9172
rect 15292 9120 15344 9172
rect 1860 9095 1912 9104
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 13452 9052 13504 9104
rect 13728 9052 13780 9104
rect 16396 9120 16448 9172
rect 19708 9120 19760 9172
rect 23388 9163 23440 9172
rect 10416 8984 10468 9036
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 8576 8891 8628 8900
rect 8576 8857 8585 8891
rect 8585 8857 8619 8891
rect 8619 8857 8628 8891
rect 12348 8916 12400 8968
rect 14004 8984 14056 9036
rect 18144 9052 18196 9104
rect 20076 9052 20128 9104
rect 22284 9052 22336 9104
rect 23112 9052 23164 9104
rect 23388 9129 23397 9163
rect 23397 9129 23431 9163
rect 23431 9129 23440 9163
rect 23388 9120 23440 9129
rect 23940 9163 23992 9172
rect 23940 9129 23949 9163
rect 23949 9129 23983 9163
rect 23983 9129 23992 9163
rect 23940 9120 23992 9129
rect 26148 9120 26200 9172
rect 26240 9120 26292 9172
rect 27436 9120 27488 9172
rect 27528 9120 27580 9172
rect 19432 8984 19484 9036
rect 8576 8848 8628 8857
rect 13268 8848 13320 8900
rect 16304 8916 16356 8968
rect 16764 8916 16816 8968
rect 20536 8916 20588 8968
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 23664 8916 23716 8968
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 26148 8916 26200 8968
rect 26700 8959 26752 8968
rect 26700 8925 26709 8959
rect 26709 8925 26743 8959
rect 26743 8925 26752 8959
rect 26700 8916 26752 8925
rect 26884 8959 26936 8968
rect 26884 8925 26893 8959
rect 26893 8925 26927 8959
rect 26927 8925 26936 8959
rect 26884 8916 26936 8925
rect 27896 9120 27948 9172
rect 27712 8984 27764 9036
rect 29736 9052 29788 9104
rect 30932 9120 30984 9172
rect 37372 9120 37424 9172
rect 28172 8984 28224 9036
rect 29828 9027 29880 9036
rect 28908 8959 28960 8968
rect 28908 8925 28917 8959
rect 28917 8925 28951 8959
rect 28951 8925 28960 8959
rect 28908 8916 28960 8925
rect 29828 8993 29837 9027
rect 29837 8993 29871 9027
rect 29871 8993 29880 9027
rect 29828 8984 29880 8993
rect 30472 9027 30524 9036
rect 30472 8993 30481 9027
rect 30481 8993 30515 9027
rect 30515 8993 30524 9027
rect 30472 8984 30524 8993
rect 29276 8916 29328 8968
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 9680 8780 9732 8832
rect 10508 8780 10560 8832
rect 12808 8780 12860 8832
rect 12992 8780 13044 8832
rect 14372 8780 14424 8832
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 16488 8848 16540 8900
rect 16672 8848 16724 8900
rect 19616 8891 19668 8900
rect 15936 8780 15988 8832
rect 17316 8780 17368 8832
rect 17960 8780 18012 8832
rect 19616 8857 19625 8891
rect 19625 8857 19659 8891
rect 19659 8857 19668 8891
rect 19616 8848 19668 8857
rect 19708 8891 19760 8900
rect 19708 8857 19717 8891
rect 19717 8857 19751 8891
rect 19751 8857 19760 8891
rect 19708 8848 19760 8857
rect 20812 8848 20864 8900
rect 24492 8848 24544 8900
rect 24584 8891 24636 8900
rect 24584 8857 24593 8891
rect 24593 8857 24627 8891
rect 24627 8857 24636 8891
rect 24584 8848 24636 8857
rect 20720 8780 20772 8832
rect 22192 8780 22244 8832
rect 25504 8848 25556 8900
rect 26424 8848 26476 8900
rect 29644 8848 29696 8900
rect 29920 8891 29972 8900
rect 29920 8857 29929 8891
rect 29929 8857 29963 8891
rect 29963 8857 29972 8891
rect 29920 8848 29972 8857
rect 27068 8780 27120 8832
rect 30932 8823 30984 8832
rect 30932 8789 30941 8823
rect 30941 8789 30975 8823
rect 30975 8789 30984 8823
rect 30932 8780 30984 8789
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 11152 8576 11204 8628
rect 12992 8576 13044 8628
rect 13084 8576 13136 8628
rect 15660 8576 15712 8628
rect 8300 8508 8352 8560
rect 13636 8508 13688 8560
rect 18604 8576 18656 8628
rect 19156 8576 19208 8628
rect 20996 8576 21048 8628
rect 16764 8508 16816 8560
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 16304 8483 16356 8492
rect 16304 8449 16306 8483
rect 16306 8449 16340 8483
rect 16340 8449 16356 8483
rect 17868 8508 17920 8560
rect 19432 8508 19484 8560
rect 20628 8508 20680 8560
rect 21272 8508 21324 8560
rect 25780 8576 25832 8628
rect 26240 8619 26292 8628
rect 26240 8585 26249 8619
rect 26249 8585 26283 8619
rect 26283 8585 26292 8619
rect 26240 8576 26292 8585
rect 26424 8576 26476 8628
rect 23756 8551 23808 8560
rect 23756 8517 23765 8551
rect 23765 8517 23799 8551
rect 23799 8517 23808 8551
rect 23756 8508 23808 8517
rect 23848 8508 23900 8560
rect 16304 8440 16356 8449
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 24124 8508 24176 8560
rect 24768 8551 24820 8560
rect 24768 8517 24777 8551
rect 24777 8517 24811 8551
rect 24811 8517 24820 8551
rect 24768 8508 24820 8517
rect 29460 8576 29512 8628
rect 30380 8619 30432 8628
rect 30380 8585 30389 8619
rect 30389 8585 30423 8619
rect 30423 8585 30432 8619
rect 30380 8576 30432 8585
rect 28264 8551 28316 8560
rect 28264 8517 28273 8551
rect 28273 8517 28307 8551
rect 28307 8517 28316 8551
rect 28264 8508 28316 8517
rect 29184 8551 29236 8560
rect 29184 8517 29193 8551
rect 29193 8517 29227 8551
rect 29227 8517 29236 8551
rect 29184 8508 29236 8517
rect 30840 8508 30892 8560
rect 21456 8440 21508 8449
rect 26240 8440 26292 8492
rect 26792 8440 26844 8492
rect 27528 8440 27580 8492
rect 29092 8440 29144 8492
rect 30748 8440 30800 8492
rect 15476 8372 15528 8424
rect 15660 8372 15712 8424
rect 17960 8372 18012 8424
rect 20168 8304 20220 8356
rect 21916 8304 21968 8356
rect 9680 8236 9732 8288
rect 14464 8236 14516 8288
rect 17592 8236 17644 8288
rect 17684 8236 17736 8288
rect 18972 8236 19024 8288
rect 19156 8236 19208 8288
rect 22284 8236 22336 8288
rect 24492 8304 24544 8356
rect 26148 8372 26200 8424
rect 27620 8372 27672 8424
rect 29368 8372 29420 8424
rect 30288 8304 30340 8356
rect 29552 8236 29604 8288
rect 29736 8279 29788 8288
rect 29736 8245 29745 8279
rect 29745 8245 29779 8279
rect 29779 8245 29788 8279
rect 29736 8236 29788 8245
rect 31024 8279 31076 8288
rect 31024 8245 31033 8279
rect 31033 8245 31067 8279
rect 31067 8245 31076 8279
rect 31576 8279 31628 8288
rect 31024 8236 31076 8245
rect 31576 8245 31585 8279
rect 31585 8245 31619 8279
rect 31619 8245 31628 8279
rect 31576 8236 31628 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 12164 8032 12216 8084
rect 13268 8032 13320 8084
rect 13728 8032 13780 8084
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 17040 8032 17092 8084
rect 17316 8032 17368 8084
rect 20536 8032 20588 8084
rect 23664 8032 23716 8084
rect 24032 8032 24084 8084
rect 24860 8032 24912 8084
rect 25596 8032 25648 8084
rect 29644 8032 29696 8084
rect 30472 8075 30524 8084
rect 30472 8041 30481 8075
rect 30481 8041 30515 8075
rect 30515 8041 30524 8075
rect 30472 8032 30524 8041
rect 31760 8075 31812 8084
rect 31760 8041 31769 8075
rect 31769 8041 31803 8075
rect 31803 8041 31812 8075
rect 31760 8032 31812 8041
rect 37740 8032 37792 8084
rect 14096 7964 14148 8016
rect 15016 7964 15068 8016
rect 13176 7896 13228 7948
rect 16304 7896 16356 7948
rect 16396 7896 16448 7948
rect 18972 7964 19024 8016
rect 17868 7896 17920 7948
rect 19432 7896 19484 7948
rect 19800 7896 19852 7948
rect 20720 7896 20772 7948
rect 22836 7896 22888 7948
rect 15200 7871 15252 7880
rect 12164 7803 12216 7812
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 12164 7769 12173 7803
rect 12173 7769 12207 7803
rect 12207 7769 12216 7803
rect 12164 7760 12216 7769
rect 13452 7760 13504 7812
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 22008 7871 22060 7880
rect 21456 7828 21508 7837
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 23940 7896 23992 7948
rect 25688 7896 25740 7948
rect 26792 7939 26844 7948
rect 26792 7905 26801 7939
rect 26801 7905 26835 7939
rect 26835 7905 26844 7939
rect 26792 7896 26844 7905
rect 27068 7939 27120 7948
rect 27068 7905 27077 7939
rect 27077 7905 27111 7939
rect 27111 7905 27120 7939
rect 27068 7896 27120 7905
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27620 7896 27672 7905
rect 29000 7896 29052 7948
rect 12532 7692 12584 7744
rect 15844 7760 15896 7812
rect 16028 7760 16080 7812
rect 16212 7760 16264 7812
rect 17592 7760 17644 7812
rect 18604 7760 18656 7812
rect 19800 7692 19852 7744
rect 20352 7692 20404 7744
rect 22192 7692 22244 7744
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 25412 7871 25464 7880
rect 24768 7828 24820 7837
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 28724 7828 28776 7880
rect 25964 7760 26016 7812
rect 27068 7760 27120 7812
rect 23664 7692 23716 7744
rect 26332 7692 26384 7744
rect 28540 7760 28592 7812
rect 29736 7760 29788 7812
rect 30748 7828 30800 7880
rect 31300 7828 31352 7880
rect 28356 7692 28408 7744
rect 28448 7692 28500 7744
rect 31392 7760 31444 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 2044 7420 2096 7472
rect 13452 7488 13504 7540
rect 15200 7488 15252 7540
rect 13360 7463 13412 7472
rect 13360 7429 13369 7463
rect 13369 7429 13403 7463
rect 13403 7429 13412 7463
rect 13360 7420 13412 7429
rect 13728 7420 13780 7472
rect 16488 7420 16540 7472
rect 1584 7352 1636 7404
rect 11796 7352 11848 7404
rect 12256 7352 12308 7404
rect 16304 7352 16356 7404
rect 17684 7420 17736 7472
rect 19064 7488 19116 7540
rect 18880 7420 18932 7472
rect 18972 7463 19024 7472
rect 18972 7429 18981 7463
rect 18981 7429 19015 7463
rect 19015 7429 19024 7463
rect 20904 7488 20956 7540
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 22376 7488 22428 7540
rect 18972 7420 19024 7429
rect 21916 7420 21968 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 23664 7488 23716 7540
rect 24216 7488 24268 7540
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 25412 7420 25464 7472
rect 25872 7420 25924 7472
rect 27160 7463 27212 7472
rect 27160 7429 27169 7463
rect 27169 7429 27203 7463
rect 27203 7429 27212 7463
rect 27160 7420 27212 7429
rect 27712 7463 27764 7472
rect 27712 7429 27721 7463
rect 27721 7429 27755 7463
rect 27755 7429 27764 7463
rect 27712 7420 27764 7429
rect 28356 7488 28408 7540
rect 28908 7488 28960 7540
rect 30564 7488 30616 7540
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 14924 7284 14976 7336
rect 17316 7284 17368 7336
rect 18512 7352 18564 7404
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 20536 7352 20588 7404
rect 21364 7352 21416 7404
rect 23388 7352 23440 7404
rect 24860 7352 24912 7404
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 28172 7352 28224 7404
rect 29184 7352 29236 7404
rect 18420 7284 18472 7336
rect 22008 7327 22060 7336
rect 12072 7216 12124 7268
rect 15568 7216 15620 7268
rect 22008 7293 22017 7327
rect 22017 7293 22051 7327
rect 22051 7293 22060 7327
rect 22008 7284 22060 7293
rect 26148 7327 26200 7336
rect 26148 7293 26157 7327
rect 26157 7293 26191 7327
rect 26191 7293 26200 7327
rect 26148 7284 26200 7293
rect 28908 7284 28960 7336
rect 21548 7216 21600 7268
rect 23480 7216 23532 7268
rect 23848 7216 23900 7268
rect 24768 7216 24820 7268
rect 27344 7216 27396 7268
rect 31116 7395 31168 7404
rect 31116 7361 31125 7395
rect 31125 7361 31159 7395
rect 31159 7361 31168 7395
rect 31116 7352 31168 7361
rect 35900 7352 35952 7404
rect 38292 7327 38344 7336
rect 38292 7293 38301 7327
rect 38301 7293 38335 7327
rect 38335 7293 38344 7327
rect 38292 7284 38344 7293
rect 31024 7259 31076 7268
rect 31024 7225 31033 7259
rect 31033 7225 31067 7259
rect 31067 7225 31076 7259
rect 31024 7216 31076 7225
rect 31576 7216 31628 7268
rect 32588 7216 32640 7268
rect 10232 7148 10284 7200
rect 12164 7148 12216 7200
rect 18604 7148 18656 7200
rect 18696 7148 18748 7200
rect 19432 7148 19484 7200
rect 19524 7148 19576 7200
rect 21088 7148 21140 7200
rect 22376 7148 22428 7200
rect 23388 7148 23440 7200
rect 27896 7148 27948 7200
rect 28080 7148 28132 7200
rect 28540 7148 28592 7200
rect 32220 7148 32272 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 14648 6944 14700 6996
rect 16396 6944 16448 6996
rect 17408 6987 17460 6996
rect 17408 6953 17438 6987
rect 17438 6953 17460 6987
rect 17408 6944 17460 6953
rect 18512 6944 18564 6996
rect 19524 6944 19576 6996
rect 20260 6944 20312 6996
rect 21272 6944 21324 6996
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 13636 6851 13688 6860
rect 12440 6740 12492 6792
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 14096 6808 14148 6860
rect 14556 6808 14608 6860
rect 15016 6808 15068 6860
rect 16304 6876 16356 6928
rect 24676 6944 24728 6996
rect 27068 6944 27120 6996
rect 27160 6944 27212 6996
rect 15844 6808 15896 6860
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 19432 6851 19484 6860
rect 19432 6817 19441 6851
rect 19441 6817 19475 6851
rect 19475 6817 19484 6851
rect 19432 6808 19484 6817
rect 9128 6715 9180 6724
rect 9128 6681 9137 6715
rect 9137 6681 9171 6715
rect 9171 6681 9180 6715
rect 9128 6672 9180 6681
rect 10784 6672 10836 6724
rect 14004 6672 14056 6724
rect 16396 6740 16448 6792
rect 23296 6808 23348 6860
rect 23756 6808 23808 6860
rect 24216 6808 24268 6860
rect 27252 6876 27304 6928
rect 27804 6944 27856 6996
rect 28724 6944 28776 6996
rect 29184 6944 29236 6996
rect 38292 6919 38344 6928
rect 23664 6740 23716 6792
rect 24768 6808 24820 6860
rect 38292 6885 38301 6919
rect 38301 6885 38335 6919
rect 38335 6885 38344 6919
rect 38292 6876 38344 6885
rect 31576 6808 31628 6860
rect 25320 6783 25372 6792
rect 14464 6672 14516 6724
rect 14832 6672 14884 6724
rect 17316 6672 17368 6724
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 12532 6604 12584 6656
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13084 6604 13136 6613
rect 14372 6604 14424 6656
rect 18972 6604 19024 6656
rect 22836 6672 22888 6724
rect 23204 6672 23256 6724
rect 24400 6672 24452 6724
rect 25320 6749 25329 6783
rect 25329 6749 25363 6783
rect 25363 6749 25372 6783
rect 25320 6740 25372 6749
rect 26700 6740 26752 6792
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 27712 6740 27764 6792
rect 28080 6740 28132 6792
rect 26148 6672 26200 6724
rect 26424 6715 26476 6724
rect 26424 6681 26433 6715
rect 26433 6681 26467 6715
rect 26467 6681 26476 6715
rect 26424 6672 26476 6681
rect 26516 6715 26568 6724
rect 26516 6681 26525 6715
rect 26525 6681 26559 6715
rect 26559 6681 26568 6715
rect 28356 6715 28408 6724
rect 26516 6672 26568 6681
rect 28356 6681 28365 6715
rect 28365 6681 28399 6715
rect 28399 6681 28408 6715
rect 28356 6672 28408 6681
rect 28448 6715 28500 6724
rect 28448 6681 28457 6715
rect 28457 6681 28491 6715
rect 28491 6681 28500 6715
rect 28448 6672 28500 6681
rect 28816 6672 28868 6724
rect 29184 6740 29236 6792
rect 29368 6740 29420 6792
rect 31116 6740 31168 6792
rect 31300 6740 31352 6792
rect 32496 6740 32548 6792
rect 20720 6604 20772 6656
rect 21180 6647 21232 6656
rect 21180 6613 21189 6647
rect 21189 6613 21223 6647
rect 21223 6613 21232 6647
rect 21180 6604 21232 6613
rect 22284 6604 22336 6656
rect 29184 6604 29236 6656
rect 30472 6647 30524 6656
rect 30472 6613 30481 6647
rect 30481 6613 30515 6647
rect 30515 6613 30524 6647
rect 30472 6604 30524 6613
rect 31116 6647 31168 6656
rect 31116 6613 31125 6647
rect 31125 6613 31159 6647
rect 31159 6613 31168 6647
rect 31116 6604 31168 6613
rect 31208 6604 31260 6656
rect 31852 6604 31904 6656
rect 32588 6604 32640 6656
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 33324 6604 33376 6656
rect 33968 6647 34020 6656
rect 33968 6613 33977 6647
rect 33977 6613 34011 6647
rect 34011 6613 34020 6647
rect 33968 6604 34020 6613
rect 37648 6647 37700 6656
rect 37648 6613 37657 6647
rect 37657 6613 37691 6647
rect 37691 6613 37700 6647
rect 37648 6604 37700 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 8300 6400 8352 6452
rect 10876 6400 10928 6452
rect 11704 6400 11756 6452
rect 13452 6400 13504 6452
rect 14004 6400 14056 6452
rect 4620 6332 4672 6384
rect 13728 6332 13780 6384
rect 15752 6400 15804 6452
rect 16488 6400 16540 6452
rect 24032 6400 24084 6452
rect 17868 6332 17920 6384
rect 4068 6264 4120 6316
rect 8024 6264 8076 6316
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9220 6264 9272 6316
rect 16028 6264 16080 6316
rect 16212 6264 16264 6316
rect 19432 6332 19484 6384
rect 19800 6332 19852 6384
rect 22284 6332 22336 6384
rect 27712 6400 27764 6452
rect 27896 6443 27948 6452
rect 27896 6409 27905 6443
rect 27905 6409 27939 6443
rect 27939 6409 27948 6443
rect 27896 6400 27948 6409
rect 28632 6443 28684 6452
rect 28632 6409 28641 6443
rect 28641 6409 28675 6443
rect 28675 6409 28684 6443
rect 28632 6400 28684 6409
rect 28724 6400 28776 6452
rect 26884 6332 26936 6384
rect 27068 6332 27120 6384
rect 30748 6400 30800 6452
rect 32404 6443 32456 6452
rect 30564 6375 30616 6384
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 13636 6196 13688 6248
rect 9772 6060 9824 6112
rect 10232 6060 10284 6112
rect 11980 6128 12032 6180
rect 13084 6128 13136 6180
rect 14556 6196 14608 6248
rect 14648 6196 14700 6248
rect 15752 6196 15804 6248
rect 18972 6196 19024 6248
rect 21364 6196 21416 6248
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22376 6196 22428 6248
rect 26240 6264 26292 6316
rect 26700 6264 26752 6316
rect 28724 6307 28776 6316
rect 28724 6273 28733 6307
rect 28733 6273 28767 6307
rect 28767 6273 28776 6307
rect 28724 6264 28776 6273
rect 29368 6307 29420 6316
rect 29368 6273 29377 6307
rect 29377 6273 29411 6307
rect 29411 6273 29420 6307
rect 29368 6264 29420 6273
rect 30564 6341 30573 6375
rect 30573 6341 30607 6375
rect 30607 6341 30616 6375
rect 30564 6332 30616 6341
rect 30104 6264 30156 6316
rect 31208 6264 31260 6316
rect 32404 6409 32413 6443
rect 32413 6409 32447 6443
rect 32447 6409 32456 6443
rect 32404 6400 32456 6409
rect 31392 6264 31444 6316
rect 32496 6307 32548 6316
rect 32496 6273 32505 6307
rect 32505 6273 32539 6307
rect 32539 6273 32548 6307
rect 32496 6264 32548 6273
rect 27436 6196 27488 6248
rect 27712 6196 27764 6248
rect 31760 6196 31812 6248
rect 15936 6128 15988 6180
rect 16488 6128 16540 6180
rect 17408 6128 17460 6180
rect 13452 6060 13504 6112
rect 17316 6060 17368 6112
rect 21732 6060 21784 6112
rect 23480 6128 23532 6180
rect 22376 6060 22428 6112
rect 23664 6060 23716 6112
rect 24032 6060 24084 6112
rect 32588 6128 32640 6180
rect 33692 6128 33744 6180
rect 25964 6103 26016 6112
rect 25964 6069 25973 6103
rect 25973 6069 26007 6103
rect 26007 6069 26016 6103
rect 25964 6060 26016 6069
rect 26056 6060 26108 6112
rect 26516 6060 26568 6112
rect 26792 6060 26844 6112
rect 29644 6060 29696 6112
rect 33324 6060 33376 6112
rect 36452 6060 36504 6112
rect 38292 6103 38344 6112
rect 38292 6069 38301 6103
rect 38301 6069 38335 6103
rect 38335 6069 38344 6103
rect 38292 6060 38344 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4620 5856 4672 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 10324 5856 10376 5908
rect 14648 5856 14700 5908
rect 16304 5899 16356 5908
rect 16304 5865 16313 5899
rect 16313 5865 16347 5899
rect 16347 5865 16356 5899
rect 16304 5856 16356 5865
rect 17408 5856 17460 5908
rect 9220 5788 9272 5840
rect 13820 5788 13872 5840
rect 18880 5831 18932 5840
rect 18880 5797 18889 5831
rect 18889 5797 18923 5831
rect 18923 5797 18932 5831
rect 18880 5788 18932 5797
rect 19340 5856 19392 5908
rect 26332 5899 26384 5908
rect 11704 5720 11756 5772
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 13912 5720 13964 5772
rect 14832 5763 14884 5772
rect 14832 5729 14841 5763
rect 14841 5729 14875 5763
rect 14875 5729 14884 5763
rect 14832 5720 14884 5729
rect 16396 5720 16448 5772
rect 17132 5763 17184 5772
rect 17132 5729 17141 5763
rect 17141 5729 17175 5763
rect 17175 5729 17184 5763
rect 17132 5720 17184 5729
rect 19524 5720 19576 5772
rect 3608 5652 3660 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 14556 5695 14608 5704
rect 9496 5627 9548 5636
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 10784 5584 10836 5636
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 19064 5652 19116 5704
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 12440 5516 12492 5568
rect 13636 5584 13688 5636
rect 14372 5516 14424 5568
rect 15752 5516 15804 5568
rect 16488 5584 16540 5636
rect 19340 5584 19392 5636
rect 26332 5865 26341 5899
rect 26341 5865 26375 5899
rect 26375 5865 26384 5899
rect 26332 5856 26384 5865
rect 26424 5856 26476 5908
rect 28264 5856 28316 5908
rect 29552 5856 29604 5908
rect 30288 5856 30340 5908
rect 31024 5856 31076 5908
rect 31760 5899 31812 5908
rect 31760 5865 31769 5899
rect 31769 5865 31803 5899
rect 31803 5865 31812 5899
rect 35440 5899 35492 5908
rect 31760 5856 31812 5865
rect 35440 5865 35449 5899
rect 35449 5865 35483 5899
rect 35483 5865 35492 5899
rect 35440 5856 35492 5865
rect 26608 5788 26660 5840
rect 26976 5788 27028 5840
rect 28080 5788 28132 5840
rect 22560 5720 22612 5772
rect 22652 5720 22704 5772
rect 30380 5788 30432 5840
rect 37464 5788 37516 5840
rect 22008 5652 22060 5704
rect 24216 5652 24268 5704
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 26240 5652 26292 5704
rect 27804 5652 27856 5704
rect 28080 5695 28132 5704
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 20260 5584 20312 5636
rect 21732 5584 21784 5636
rect 21916 5516 21968 5568
rect 24492 5584 24544 5636
rect 24860 5627 24912 5636
rect 24860 5593 24869 5627
rect 24869 5593 24903 5627
rect 24903 5593 24912 5627
rect 24860 5584 24912 5593
rect 26148 5584 26200 5636
rect 31116 5720 31168 5772
rect 30104 5652 30156 5704
rect 30472 5652 30524 5704
rect 32496 5695 32548 5704
rect 32496 5661 32505 5695
rect 32505 5661 32539 5695
rect 32539 5661 32548 5695
rect 32496 5652 32548 5661
rect 32864 5652 32916 5704
rect 33324 5652 33376 5704
rect 35256 5652 35308 5704
rect 30380 5584 30432 5636
rect 38200 5627 38252 5636
rect 38200 5593 38209 5627
rect 38209 5593 38243 5627
rect 38243 5593 38252 5627
rect 38200 5584 38252 5593
rect 27436 5516 27488 5568
rect 29736 5516 29788 5568
rect 33048 5559 33100 5568
rect 33048 5525 33057 5559
rect 33057 5525 33091 5559
rect 33091 5525 33100 5559
rect 33048 5516 33100 5525
rect 33600 5559 33652 5568
rect 33600 5525 33609 5559
rect 33609 5525 33643 5559
rect 33643 5525 33652 5559
rect 33600 5516 33652 5525
rect 36084 5559 36136 5568
rect 36084 5525 36093 5559
rect 36093 5525 36127 5559
rect 36127 5525 36136 5559
rect 36084 5516 36136 5525
rect 36452 5516 36504 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 10416 5312 10468 5364
rect 12348 5312 12400 5364
rect 11888 5244 11940 5296
rect 12440 5244 12492 5296
rect 16028 5312 16080 5364
rect 16304 5312 16356 5364
rect 17316 5312 17368 5364
rect 1952 5176 2004 5228
rect 10140 5176 10192 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 15016 5244 15068 5296
rect 15476 5287 15528 5296
rect 15476 5253 15485 5287
rect 15485 5253 15519 5287
rect 15519 5253 15528 5287
rect 19892 5312 19944 5364
rect 23848 5355 23900 5364
rect 23848 5321 23857 5355
rect 23857 5321 23891 5355
rect 23891 5321 23900 5355
rect 23848 5312 23900 5321
rect 23940 5312 23992 5364
rect 25688 5355 25740 5364
rect 25688 5321 25697 5355
rect 25697 5321 25731 5355
rect 25731 5321 25740 5355
rect 25688 5312 25740 5321
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 27712 5312 27764 5364
rect 28448 5312 28500 5364
rect 29920 5355 29972 5364
rect 29920 5321 29929 5355
rect 29929 5321 29963 5355
rect 29963 5321 29972 5355
rect 29920 5312 29972 5321
rect 30564 5355 30616 5364
rect 30564 5321 30573 5355
rect 30573 5321 30607 5355
rect 30607 5321 30616 5355
rect 30564 5312 30616 5321
rect 34152 5355 34204 5364
rect 34152 5321 34161 5355
rect 34161 5321 34195 5355
rect 34195 5321 34204 5355
rect 34152 5312 34204 5321
rect 35256 5355 35308 5364
rect 35256 5321 35265 5355
rect 35265 5321 35299 5355
rect 35299 5321 35308 5355
rect 35256 5312 35308 5321
rect 19248 5287 19300 5296
rect 15476 5244 15528 5253
rect 19248 5253 19257 5287
rect 19257 5253 19291 5287
rect 19291 5253 19300 5287
rect 19248 5244 19300 5253
rect 22652 5244 22704 5296
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 17132 5176 17184 5228
rect 19800 5176 19852 5228
rect 24676 5219 24728 5228
rect 8024 4972 8076 5024
rect 8484 4972 8536 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 14188 5108 14240 5160
rect 15108 5108 15160 5160
rect 15384 5108 15436 5160
rect 13268 5040 13320 5092
rect 14280 5040 14332 5092
rect 15476 4972 15528 5024
rect 19248 5040 19300 5092
rect 19984 5040 20036 5092
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23020 5108 23072 5160
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 30380 5244 30432 5296
rect 25872 5219 25924 5228
rect 25872 5185 25881 5219
rect 25881 5185 25915 5219
rect 25915 5185 25924 5219
rect 25872 5176 25924 5185
rect 21824 5040 21876 5092
rect 20076 4972 20128 5024
rect 22468 4972 22520 5024
rect 23572 4972 23624 5024
rect 24584 4972 24636 5024
rect 25320 4972 25372 5024
rect 27988 5176 28040 5228
rect 28632 5176 28684 5228
rect 28724 5219 28776 5228
rect 28724 5185 28733 5219
rect 28733 5185 28767 5219
rect 28767 5185 28776 5219
rect 28724 5176 28776 5185
rect 29184 5176 29236 5228
rect 29828 5219 29880 5228
rect 29828 5185 29837 5219
rect 29837 5185 29871 5219
rect 29871 5185 29880 5219
rect 29828 5176 29880 5185
rect 30472 5176 30524 5228
rect 27620 5108 27672 5160
rect 31208 5176 31260 5228
rect 31392 5176 31444 5228
rect 32588 5176 32640 5228
rect 33232 5176 33284 5228
rect 32312 5108 32364 5160
rect 26792 5040 26844 5092
rect 29736 5040 29788 5092
rect 32404 5083 32456 5092
rect 32404 5049 32413 5083
rect 32413 5049 32447 5083
rect 32447 5049 32456 5083
rect 32404 5040 32456 5049
rect 27896 4972 27948 5024
rect 28448 4972 28500 5024
rect 28816 4972 28868 5024
rect 29184 4972 29236 5024
rect 30288 4972 30340 5024
rect 31668 4972 31720 5024
rect 33600 5015 33652 5024
rect 33600 4981 33609 5015
rect 33609 4981 33643 5015
rect 33643 4981 33652 5015
rect 33600 4972 33652 4981
rect 36452 4972 36504 5024
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 10048 4768 10100 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 11612 4768 11664 4820
rect 13544 4811 13596 4820
rect 9588 4700 9640 4752
rect 13268 4700 13320 4752
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14648 4768 14700 4820
rect 14832 4768 14884 4820
rect 18328 4768 18380 4820
rect 14556 4700 14608 4752
rect 8944 4632 8996 4684
rect 14280 4632 14332 4684
rect 17040 4675 17092 4684
rect 17040 4641 17049 4675
rect 17049 4641 17083 4675
rect 17083 4641 17092 4675
rect 17040 4632 17092 4641
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 8116 4564 8168 4616
rect 29460 4768 29512 4820
rect 30196 4768 30248 4820
rect 31208 4768 31260 4820
rect 31668 4768 31720 4820
rect 31760 4811 31812 4820
rect 31760 4777 31769 4811
rect 31769 4777 31803 4811
rect 31803 4777 31812 4811
rect 31760 4768 31812 4777
rect 18512 4700 18564 4752
rect 19340 4700 19392 4752
rect 21180 4743 21232 4752
rect 21180 4709 21189 4743
rect 21189 4709 21223 4743
rect 21223 4709 21232 4743
rect 21180 4700 21232 4709
rect 21456 4700 21508 4752
rect 24492 4700 24544 4752
rect 27712 4700 27764 4752
rect 28264 4700 28316 4752
rect 30012 4700 30064 4752
rect 31484 4700 31536 4752
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 19800 4632 19852 4684
rect 13636 4539 13688 4548
rect 13636 4505 13645 4539
rect 13645 4505 13679 4539
rect 13679 4505 13688 4539
rect 13636 4496 13688 4505
rect 13728 4496 13780 4548
rect 23572 4564 23624 4616
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 26056 4564 26108 4616
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 14096 4428 14148 4480
rect 14556 4428 14608 4480
rect 22192 4496 22244 4548
rect 22284 4539 22336 4548
rect 22284 4505 22293 4539
rect 22293 4505 22327 4539
rect 22327 4505 22336 4539
rect 22284 4496 22336 4505
rect 22560 4496 22612 4548
rect 26424 4539 26476 4548
rect 26424 4505 26433 4539
rect 26433 4505 26467 4539
rect 26467 4505 26476 4539
rect 26424 4496 26476 4505
rect 27896 4564 27948 4616
rect 30196 4632 30248 4684
rect 28908 4564 28960 4616
rect 29552 4564 29604 4616
rect 30472 4564 30524 4616
rect 30656 4564 30708 4616
rect 31300 4564 31352 4616
rect 31852 4607 31904 4616
rect 31852 4573 31861 4607
rect 31861 4573 31895 4607
rect 31895 4573 31904 4607
rect 31852 4564 31904 4573
rect 33232 4632 33284 4684
rect 33692 4675 33744 4684
rect 33692 4641 33701 4675
rect 33701 4641 33735 4675
rect 33735 4641 33744 4675
rect 33692 4632 33744 4641
rect 34336 4632 34388 4684
rect 26792 4496 26844 4548
rect 27344 4539 27396 4548
rect 27344 4505 27353 4539
rect 27353 4505 27387 4539
rect 27387 4505 27396 4539
rect 27344 4496 27396 4505
rect 23664 4428 23716 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24308 4428 24360 4480
rect 24492 4428 24544 4480
rect 25044 4428 25096 4480
rect 27712 4496 27764 4548
rect 27620 4428 27672 4480
rect 29644 4428 29696 4480
rect 31484 4496 31536 4548
rect 32404 4539 32456 4548
rect 30012 4428 30064 4480
rect 32404 4505 32413 4539
rect 32413 4505 32447 4539
rect 32447 4505 32456 4539
rect 32404 4496 32456 4505
rect 34796 4496 34848 4548
rect 38016 4564 38068 4616
rect 36452 4496 36504 4548
rect 33600 4428 33652 4480
rect 35716 4428 35768 4480
rect 38108 4471 38160 4480
rect 38108 4437 38117 4471
rect 38117 4437 38151 4471
rect 38151 4437 38160 4471
rect 38108 4428 38160 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 11980 4224 12032 4276
rect 14372 4224 14424 4276
rect 19248 4224 19300 4276
rect 13360 4156 13412 4208
rect 14740 4156 14792 4208
rect 12532 4088 12584 4140
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 8024 3952 8076 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 4068 3884 4120 3936
rect 6920 3884 6972 3936
rect 7012 3884 7064 3936
rect 8668 3884 8720 3936
rect 10324 4020 10376 4072
rect 12716 3952 12768 4004
rect 11060 3884 11112 3936
rect 11244 3884 11296 3936
rect 14188 4020 14240 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 17040 4088 17092 4140
rect 18972 4088 19024 4140
rect 17868 4063 17920 4072
rect 17868 4029 17877 4063
rect 17877 4029 17911 4063
rect 17911 4029 17920 4063
rect 21180 4156 21232 4208
rect 19248 4088 19300 4140
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 17868 4020 17920 4029
rect 22284 4224 22336 4276
rect 24860 4224 24912 4276
rect 25504 4224 25556 4276
rect 29828 4224 29880 4276
rect 22192 4156 22244 4208
rect 24124 4156 24176 4208
rect 24584 4156 24636 4208
rect 27436 4156 27488 4208
rect 36452 4267 36504 4276
rect 36452 4233 36461 4267
rect 36461 4233 36495 4267
rect 36495 4233 36504 4267
rect 36452 4224 36504 4233
rect 21364 4020 21416 4072
rect 22376 4020 22428 4072
rect 19156 3952 19208 4004
rect 20720 3952 20772 4004
rect 22008 3952 22060 4004
rect 16764 3884 16816 3936
rect 19984 3927 20036 3936
rect 19984 3893 19993 3927
rect 19993 3893 20027 3927
rect 20027 3893 20036 3927
rect 19984 3884 20036 3893
rect 21732 3884 21784 3936
rect 23020 3884 23072 3936
rect 24124 4020 24176 4072
rect 26240 4088 26292 4140
rect 26700 4088 26752 4140
rect 28816 4088 28868 4140
rect 29000 4088 29052 4140
rect 26148 4020 26200 4072
rect 27528 4063 27580 4072
rect 26424 3952 26476 4004
rect 26608 3952 26660 4004
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 27804 4063 27856 4072
rect 27804 4029 27813 4063
rect 27813 4029 27847 4063
rect 27847 4029 27856 4063
rect 27804 4020 27856 4029
rect 28540 4020 28592 4072
rect 25964 3884 26016 3936
rect 26148 3884 26200 3936
rect 26976 3884 27028 3936
rect 28080 3884 28132 3936
rect 30196 4131 30248 4140
rect 29276 4020 29328 4072
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 30288 4088 30340 4140
rect 31484 4131 31536 4140
rect 30104 4020 30156 4072
rect 31484 4097 31493 4131
rect 31493 4097 31527 4131
rect 31527 4097 31536 4131
rect 31484 4088 31536 4097
rect 32128 4088 32180 4140
rect 33324 4156 33376 4208
rect 32588 4088 32640 4140
rect 38292 4156 38344 4208
rect 35716 4088 35768 4140
rect 37924 4088 37976 4140
rect 30196 3884 30248 3936
rect 30748 3927 30800 3936
rect 30748 3893 30757 3927
rect 30757 3893 30791 3927
rect 30791 3893 30800 3927
rect 30748 3884 30800 3893
rect 36268 4020 36320 4072
rect 31576 3952 31628 4004
rect 32128 3884 32180 3936
rect 32404 3927 32456 3936
rect 32404 3893 32413 3927
rect 32413 3893 32447 3927
rect 32447 3893 32456 3927
rect 32404 3884 32456 3893
rect 32680 3884 32732 3936
rect 33692 3927 33744 3936
rect 33692 3893 33701 3927
rect 33701 3893 33735 3927
rect 33735 3893 33744 3927
rect 33692 3884 33744 3893
rect 33784 3884 33836 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 5448 3612 5500 3664
rect 9772 3680 9824 3732
rect 10048 3680 10100 3732
rect 10324 3723 10376 3732
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 12440 3680 12492 3732
rect 12624 3680 12676 3732
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 4068 3476 4120 3528
rect 8116 3544 8168 3596
rect 10968 3544 11020 3596
rect 8208 3476 8260 3528
rect 10048 3476 10100 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 13268 3612 13320 3664
rect 11336 3544 11388 3596
rect 11888 3544 11940 3596
rect 12716 3544 12768 3596
rect 13636 3612 13688 3664
rect 14280 3612 14332 3664
rect 13728 3587 13780 3596
rect 10140 3476 10192 3485
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 16120 3544 16172 3596
rect 14096 3476 14148 3528
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 3240 3340 3292 3392
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 7012 3340 7064 3392
rect 8392 3340 8444 3392
rect 8944 3340 8996 3392
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11152 3340 11204 3349
rect 11520 3408 11572 3460
rect 12256 3451 12308 3460
rect 12256 3417 12265 3451
rect 12265 3417 12299 3451
rect 12299 3417 12308 3451
rect 12256 3408 12308 3417
rect 12532 3408 12584 3460
rect 13544 3408 13596 3460
rect 16212 3408 16264 3460
rect 16580 3340 16632 3392
rect 17224 3680 17276 3732
rect 21732 3680 21784 3732
rect 21824 3680 21876 3732
rect 18144 3612 18196 3664
rect 22192 3544 22244 3596
rect 16856 3408 16908 3460
rect 19984 3408 20036 3460
rect 20076 3408 20128 3460
rect 20536 3451 20588 3460
rect 20536 3417 20545 3451
rect 20545 3417 20579 3451
rect 20579 3417 20588 3451
rect 20536 3408 20588 3417
rect 21824 3408 21876 3460
rect 22376 3408 22428 3460
rect 24952 3544 25004 3596
rect 25228 3544 25280 3596
rect 26608 3544 26660 3596
rect 27344 3680 27396 3732
rect 32588 3680 32640 3732
rect 33784 3680 33836 3732
rect 34336 3723 34388 3732
rect 34336 3689 34345 3723
rect 34345 3689 34379 3723
rect 34379 3689 34388 3723
rect 34336 3680 34388 3689
rect 35716 3680 35768 3732
rect 27436 3612 27488 3664
rect 30932 3612 30984 3664
rect 31852 3612 31904 3664
rect 24584 3519 24636 3528
rect 17040 3340 17092 3392
rect 18420 3340 18472 3392
rect 19432 3340 19484 3392
rect 20720 3340 20772 3392
rect 21272 3340 21324 3392
rect 23204 3340 23256 3392
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 25964 3476 26016 3528
rect 27528 3519 27580 3528
rect 27528 3485 27537 3519
rect 27537 3485 27571 3519
rect 27571 3485 27580 3519
rect 27528 3476 27580 3485
rect 27988 3476 28040 3528
rect 28172 3519 28224 3528
rect 28172 3485 28181 3519
rect 28181 3485 28215 3519
rect 28215 3485 28224 3519
rect 28172 3476 28224 3485
rect 28356 3476 28408 3528
rect 28908 3476 28960 3528
rect 24216 3408 24268 3460
rect 25136 3408 25188 3460
rect 25688 3340 25740 3392
rect 26516 3408 26568 3460
rect 26424 3340 26476 3392
rect 26976 3451 27028 3460
rect 26976 3417 26985 3451
rect 26985 3417 27019 3451
rect 27019 3417 27028 3451
rect 26976 3408 27028 3417
rect 27712 3408 27764 3460
rect 30288 3476 30340 3528
rect 31024 3476 31076 3528
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 33876 3612 33928 3664
rect 34796 3612 34848 3664
rect 33324 3544 33376 3596
rect 32864 3476 32916 3528
rect 29368 3340 29420 3392
rect 31668 3408 31720 3460
rect 33232 3476 33284 3528
rect 34428 3476 34480 3528
rect 36452 3476 36504 3528
rect 30472 3383 30524 3392
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 31760 3340 31812 3392
rect 33232 3340 33284 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 3424 3136 3476 3188
rect 8024 3136 8076 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 11796 3136 11848 3188
rect 13544 3136 13596 3188
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 4068 3000 4120 3052
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 7932 2932 7984 2984
rect 10508 3068 10560 3120
rect 10692 3068 10744 3120
rect 10968 3068 11020 3120
rect 13728 3068 13780 3120
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 10048 3000 10100 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11612 3000 11664 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12440 3000 12492 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 16580 3136 16632 3188
rect 16672 3136 16724 3188
rect 19432 3136 19484 3188
rect 16120 3068 16172 3120
rect 14096 3000 14148 3009
rect 4712 2864 4764 2916
rect 5908 2864 5960 2916
rect 6736 2864 6788 2916
rect 8208 2864 8260 2916
rect 12532 2932 12584 2984
rect 13820 2932 13872 2984
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 6000 2796 6052 2805
rect 6920 2796 6972 2848
rect 8392 2796 8444 2848
rect 9588 2796 9640 2848
rect 11888 2796 11940 2848
rect 17224 3068 17276 3120
rect 19156 3068 19208 3120
rect 16580 3000 16632 3052
rect 19432 3000 19484 3052
rect 20076 3068 20128 3120
rect 22928 3136 22980 3188
rect 24216 3136 24268 3188
rect 24676 3136 24728 3188
rect 26148 3136 26200 3188
rect 22192 3068 22244 3120
rect 22284 3111 22336 3120
rect 22284 3077 22293 3111
rect 22293 3077 22327 3111
rect 22327 3077 22336 3111
rect 22284 3068 22336 3077
rect 24400 3068 24452 3120
rect 38108 3136 38160 3188
rect 18880 2932 18932 2984
rect 19064 2864 19116 2916
rect 26148 3000 26200 3052
rect 26608 3043 26660 3052
rect 26608 3009 26617 3043
rect 26617 3009 26651 3043
rect 26651 3009 26660 3043
rect 26608 3000 26660 3009
rect 22284 2932 22336 2984
rect 22376 2932 22428 2984
rect 25320 2932 25372 2984
rect 25596 2932 25648 2984
rect 26056 2932 26108 2984
rect 27712 3000 27764 3052
rect 28816 3000 28868 3052
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 31852 3068 31904 3120
rect 33692 3111 33744 3120
rect 30932 3043 30984 3052
rect 30932 3009 30941 3043
rect 30941 3009 30975 3043
rect 30975 3009 30984 3043
rect 30932 3000 30984 3009
rect 31024 3043 31076 3052
rect 31024 3009 31033 3043
rect 31033 3009 31067 3043
rect 31067 3009 31076 3043
rect 31024 3000 31076 3009
rect 33692 3077 33701 3111
rect 33701 3077 33735 3111
rect 33735 3077 33744 3111
rect 33692 3068 33744 3077
rect 36268 3111 36320 3120
rect 36268 3077 36277 3111
rect 36277 3077 36311 3111
rect 36311 3077 36320 3111
rect 36268 3068 36320 3077
rect 33876 3000 33928 3052
rect 34428 3043 34480 3052
rect 34428 3009 34437 3043
rect 34437 3009 34471 3043
rect 34471 3009 34480 3043
rect 34428 3000 34480 3009
rect 21916 2796 21968 2848
rect 24124 2864 24176 2916
rect 23664 2796 23716 2848
rect 24492 2796 24544 2848
rect 25044 2796 25096 2848
rect 27804 2975 27856 2984
rect 27804 2941 27813 2975
rect 27813 2941 27847 2975
rect 27847 2941 27856 2975
rect 27804 2932 27856 2941
rect 30564 2932 30616 2984
rect 36452 3000 36504 3052
rect 36912 3000 36964 3052
rect 32404 2907 32456 2916
rect 32404 2873 32413 2907
rect 32413 2873 32447 2907
rect 32447 2873 32456 2907
rect 32404 2864 32456 2873
rect 32496 2864 32548 2916
rect 26516 2839 26568 2848
rect 26516 2805 26525 2839
rect 26525 2805 26559 2839
rect 26559 2805 26568 2839
rect 26516 2796 26568 2805
rect 26608 2796 26660 2848
rect 28080 2796 28132 2848
rect 28816 2796 28868 2848
rect 29000 2839 29052 2848
rect 29000 2805 29009 2839
rect 29009 2805 29043 2839
rect 29043 2805 29052 2839
rect 29000 2796 29052 2805
rect 31208 2796 31260 2848
rect 32312 2796 32364 2848
rect 33048 2839 33100 2848
rect 33048 2805 33057 2839
rect 33057 2805 33091 2839
rect 33091 2805 33100 2839
rect 33048 2796 33100 2805
rect 34520 2796 34572 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 6920 2592 6972 2644
rect 20 2524 72 2576
rect 2412 2388 2464 2440
rect 5448 2456 5500 2508
rect 5908 2524 5960 2576
rect 6736 2456 6788 2508
rect 3240 2388 3292 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 8208 2320 8260 2372
rect 9680 2388 9732 2440
rect 31484 2592 31536 2644
rect 34336 2592 34388 2644
rect 35808 2635 35860 2644
rect 35808 2601 35817 2635
rect 35817 2601 35851 2635
rect 35851 2601 35860 2635
rect 35808 2592 35860 2601
rect 11336 2524 11388 2576
rect 12256 2524 12308 2576
rect 16856 2524 16908 2576
rect 21180 2524 21232 2576
rect 14096 2456 14148 2508
rect 15844 2456 15896 2508
rect 17316 2456 17368 2508
rect 19432 2456 19484 2508
rect 19892 2456 19944 2508
rect 22100 2499 22152 2508
rect 22100 2465 22109 2499
rect 22109 2465 22143 2499
rect 22143 2465 22152 2499
rect 22100 2456 22152 2465
rect 23388 2456 23440 2508
rect 30472 2524 30524 2576
rect 32312 2567 32364 2576
rect 32312 2533 32321 2567
rect 32321 2533 32355 2567
rect 32355 2533 32364 2567
rect 32312 2524 32364 2533
rect 33508 2524 33560 2576
rect 24492 2456 24544 2508
rect 25044 2499 25096 2508
rect 25044 2465 25053 2499
rect 25053 2465 25087 2499
rect 25087 2465 25096 2499
rect 25044 2456 25096 2465
rect 26516 2456 26568 2508
rect 26332 2388 26384 2440
rect 28264 2456 28316 2508
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 28356 2388 28408 2440
rect 30564 2456 30616 2508
rect 28908 2388 28960 2440
rect 31392 2456 31444 2508
rect 32220 2456 32272 2508
rect 33876 2456 33928 2508
rect 37648 2456 37700 2508
rect 31576 2388 31628 2440
rect 32588 2388 32640 2440
rect 33508 2388 33560 2440
rect 33968 2388 34020 2440
rect 35440 2388 35492 2440
rect 36084 2388 36136 2440
rect 36728 2388 36780 2440
rect 36912 2431 36964 2440
rect 36912 2397 36921 2431
rect 36921 2397 36955 2431
rect 36955 2397 36964 2431
rect 36912 2388 36964 2397
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 1308 2252 1360 2304
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 6460 2252 6512 2304
rect 11152 2320 11204 2372
rect 13452 2363 13504 2372
rect 13452 2329 13461 2363
rect 13461 2329 13495 2363
rect 13495 2329 13504 2363
rect 13452 2320 13504 2329
rect 15292 2320 15344 2372
rect 17868 2320 17920 2372
rect 19064 2320 19116 2372
rect 19340 2320 19392 2372
rect 11244 2252 11296 2304
rect 16672 2252 16724 2304
rect 22284 2320 22336 2372
rect 26148 2320 26200 2372
rect 20628 2252 20680 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 28448 2252 28500 2304
rect 29644 2252 29696 2304
rect 30564 2295 30616 2304
rect 30564 2261 30573 2295
rect 30573 2261 30607 2295
rect 30607 2261 30616 2295
rect 30564 2252 30616 2261
rect 31208 2295 31260 2304
rect 31208 2261 31217 2295
rect 31217 2261 31251 2295
rect 31251 2261 31260 2295
rect 31208 2252 31260 2261
rect 34796 2252 34848 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3424 2048 3476 2100
rect 9680 2048 9732 2100
rect 24584 2048 24636 2100
rect 27160 2048 27212 2100
rect 28172 2048 28224 2100
rect 8208 1980 8260 2032
rect 10600 1980 10652 2032
rect 24952 1980 25004 2032
rect 30564 1980 30616 2032
rect 5448 1912 5500 1964
rect 15292 1912 15344 1964
rect 25780 1912 25832 1964
rect 31208 1912 31260 1964
rect 37740 1912 37792 1964
rect 22284 1844 22336 1896
rect 33048 1844 33100 1896
rect 20536 1776 20588 1828
rect 24308 1776 24360 1828
rect 32220 1776 32272 1828
<< metal2 >>
rect 18 39200 74 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18694 39200 18750 39800
rect 20626 39200 20682 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 32 36378 60 39200
rect 1964 37262 1992 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2884 37262 2912 38791
rect 2964 37664 3016 37670
rect 2964 37606 3016 37612
rect 2976 37466 3004 37606
rect 2964 37460 3016 37466
rect 2964 37402 3016 37408
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 2872 37256 2924 37262
rect 2872 37198 2924 37204
rect 1674 36816 1730 36825
rect 1674 36751 1676 36760
rect 1728 36751 1730 36760
rect 1676 36722 1728 36728
rect 1768 36576 1820 36582
rect 1768 36518 1820 36524
rect 1780 36378 1808 36518
rect 20 36372 72 36378
rect 20 36314 72 36320
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1964 36310 1992 37198
rect 2884 36922 2912 37198
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5184 37126 5212 39200
rect 7116 37330 7144 39200
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 5264 37256 5316 37262
rect 5264 37198 5316 37204
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 5172 37120 5224 37126
rect 5172 37062 5224 37068
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 1952 36304 2004 36310
rect 1952 36246 2004 36252
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1688 33425 1716 33458
rect 1674 33416 1730 33425
rect 1674 33351 1730 33360
rect 1688 33114 1716 33351
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 5276 33114 5304 37198
rect 8404 37126 8432 39200
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 5448 36168 5500 36174
rect 5448 36110 5500 36116
rect 1676 33108 1728 33114
rect 1676 33050 1728 33056
rect 5264 33108 5316 33114
rect 5264 33050 5316 33056
rect 5460 32842 5488 36110
rect 5448 32836 5500 32842
rect 5448 32778 5500 32784
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31414 1624 31758
rect 1584 31408 1636 31414
rect 1582 31376 1584 31385
rect 1636 31376 1638 31385
rect 1582 31311 1638 31320
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 1584 30184 1636 30190
rect 1584 30126 1636 30132
rect 2504 30184 2556 30190
rect 2504 30126 2556 30132
rect 1596 30025 1624 30126
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 29850 1624 29951
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1676 24608 1728 24614
rect 1674 24576 1676 24585
rect 1728 24576 1730 24585
rect 1674 24511 1730 24520
rect 1872 23322 1900 28018
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1674 22536 1730 22545
rect 1674 22471 1676 22480
rect 1728 22471 1730 22480
rect 1676 22442 1728 22448
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1596 21185 1624 21490
rect 1582 21176 1638 21185
rect 1582 21111 1584 21120
rect 1636 21111 1638 21120
rect 1584 21082 1636 21088
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 19145 1624 19246
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1596 18970 1624 19071
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17785 1716 18022
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1780 15162 1808 22578
rect 1860 21412 1912 21418
rect 1860 21354 1912 21360
rect 1872 20466 1900 21354
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1872 14890 1900 18226
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 13938 1716 14214
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1688 13705 1716 13874
rect 1674 13696 1730 13705
rect 1674 13631 1730 13640
rect 1964 13462 1992 19314
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1674 8936 1730 8945
rect 1674 8871 1676 8880
rect 1728 8871 1730 8880
rect 1676 8842 1728 8848
rect 1688 8634 1716 8842
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1780 6914 1808 13126
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 9110 1900 10950
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 2056 7478 2084 16730
rect 2424 15502 2452 22918
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 12986 2176 14962
rect 2516 13190 2544 30126
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6840 21894 6868 26930
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2148 6914 2176 12922
rect 2516 12918 2544 13126
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 1582 6896 1638 6905
rect 1780 6886 1900 6914
rect 1582 6831 1638 6840
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4865 1624 5102
rect 1582 4856 1638 4865
rect 1582 4791 1584 4800
rect 1636 4791 1638 4800
rect 1584 4762 1636 4768
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3534 1716 3878
rect 1676 3528 1728 3534
rect 1674 3496 1676 3505
rect 1728 3496 1730 3505
rect 1674 3431 1730 3440
rect 1872 3058 1900 6886
rect 1964 6886 2176 6914
rect 1964 5234 1992 6886
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2424 2446 2452 3130
rect 3252 2446 3280 3334
rect 3436 3194 3464 17274
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15162 4108 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 7392 15026 7420 37062
rect 9312 33380 9364 33386
rect 9312 33322 9364 33328
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 7760 12918 7788 13738
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5552 12442 5580 12786
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 8404 11150 8432 11698
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 8312 6458 8340 8502
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 5710 4108 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 6326
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8036 5914 8064 6258
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3620 5370 3648 5646
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 8036 5114 8064 5850
rect 7944 5086 8064 5114
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 4080 3534 4108 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4080 3058 4108 3470
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2446 4752 2858
rect 5460 2514 5488 3606
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5920 2582 5948 2858
rect 6012 2854 6040 3334
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6012 2650 6040 2790
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 6748 2514 6776 2858
rect 6932 2854 6960 3878
rect 7024 3398 7052 3878
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7944 2990 7972 5086
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8036 4486 8064 4966
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4010 8064 4422
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8128 3641 8156 4558
rect 8114 3632 8170 3641
rect 8114 3567 8116 3576
rect 8168 3567 8170 3576
rect 8116 3538 8168 3544
rect 8128 3507 8156 3538
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 3058 8064 3130
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2650 6960 2790
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 8036 2446 8064 2994
rect 8220 2922 8248 3470
rect 8404 3398 8432 11086
rect 8588 8906 8616 12038
rect 9232 11762 9260 32710
rect 9324 13258 9352 33322
rect 9416 26586 9444 37198
rect 9496 37188 9548 37194
rect 9496 37130 9548 37136
rect 9508 32026 9536 37130
rect 10336 37126 10364 39200
rect 10692 37256 10744 37262
rect 10692 37198 10744 37204
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10704 36922 10732 37198
rect 12268 37108 12296 39200
rect 13556 37466 13584 39200
rect 13544 37460 13596 37466
rect 13544 37402 13596 37408
rect 13556 37330 13584 37402
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 12440 37120 12492 37126
rect 12268 37080 12440 37108
rect 12440 37062 12492 37068
rect 14292 36922 14320 37198
rect 15488 37126 15516 39200
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 14280 36916 14332 36922
rect 14280 36858 14332 36864
rect 13820 36372 13872 36378
rect 13820 36314 13872 36320
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 10508 31816 10560 31822
rect 10506 31784 10508 31793
rect 10560 31784 10562 31793
rect 10506 31719 10562 31728
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 13462 9904 21830
rect 12084 16574 12112 29106
rect 12084 16546 12204 16574
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10704 15706 10732 15982
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10244 12238 10272 13194
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9784 11801 9812 12106
rect 9770 11792 9826 11801
rect 9220 11756 9272 11762
rect 9770 11727 9826 11736
rect 9220 11698 9272 11704
rect 9876 11218 9904 12106
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9968 11354 9996 11766
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 9586 8708 10406
rect 9416 10266 9444 10610
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9600 10198 9628 10950
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 10152 10130 10180 12174
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9864 9648 9916 9654
rect 9862 9616 9864 9625
rect 9916 9616 9918 9625
rect 8668 9580 8720 9586
rect 9862 9551 9918 9560
rect 8668 9522 8720 9528
rect 8680 9382 8708 9522
rect 9310 9480 9366 9489
rect 9310 9415 9312 9424
rect 9364 9415 9366 9424
rect 9312 9386 9364 9392
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5030 8524 5510
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8680 3942 8708 9318
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8294 9720 8774
rect 9680 8288 9732 8294
rect 10244 8242 10272 12174
rect 10336 10674 10364 13262
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10428 11898 10456 12854
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10520 11762 10548 13670
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9680 8230 9732 8236
rect 9692 7750 9720 8230
rect 10152 8214 10272 8242
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 6322 9168 6666
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9232 5846 9260 6258
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9494 5672 9550 5681
rect 9494 5607 9496 5616
rect 9548 5607 9550 5616
rect 9496 5578 9548 5584
rect 9784 5409 9812 6054
rect 9770 5400 9826 5409
rect 9770 5335 9826 5344
rect 10152 5234 10180 8214
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 6662 10272 7142
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10244 6118 10272 6598
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10336 5914 10364 10610
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 5370 10456 8978
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 8956 4690 8984 4966
rect 10060 4826 10088 4966
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3058 8984 3334
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 9600 2854 9628 4694
rect 10060 4282 10088 4762
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10060 3738 10088 4218
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9784 3194 9812 3674
rect 10152 3534 10180 5170
rect 10428 4865 10456 5306
rect 10414 4856 10470 4865
rect 10414 4791 10470 4800
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10336 3738 10364 4014
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 10060 3058 10088 3470
rect 10520 3126 10548 8774
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2382
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2106 3464 2246
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 4724 1850 4752 2382
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5460 1970 5488 2246
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 4540 1822 4752 1850
rect 4540 800 4568 1822
rect 6472 800 6500 2246
rect 8220 2038 8248 2314
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8404 800 8432 2790
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 2106 9720 2382
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9692 800 9720 2042
rect 10612 2038 10640 15438
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 3126 10732 13194
rect 10796 11694 10824 14894
rect 10888 14074 10916 16390
rect 12176 15366 12204 16546
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13648 15706 13676 16458
rect 13832 16250 13860 36314
rect 15856 32230 15884 37198
rect 16776 37126 16804 39200
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 17144 26897 17172 37198
rect 18432 34202 18460 37198
rect 18708 35834 18736 39200
rect 20536 37392 20588 37398
rect 20536 37334 20588 37340
rect 19340 37188 19392 37194
rect 19340 37130 19392 37136
rect 19352 36786 19380 37130
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 18788 36712 18840 36718
rect 18788 36654 18840 36660
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 17684 33856 17736 33862
rect 17684 33798 17736 33804
rect 17130 26888 17186 26897
rect 17130 26823 17186 26832
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13832 16130 13860 16186
rect 13832 16102 13952 16130
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13832 15502 13860 15982
rect 13924 15570 13952 16102
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14346 11284 14758
rect 11716 14550 11744 14962
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10888 13954 10916 14010
rect 11060 14000 11112 14006
rect 10888 13926 11008 13954
rect 11060 13942 11112 13948
rect 10980 13326 11008 13926
rect 11072 13530 11100 13942
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11716 12238 11744 14486
rect 12176 14414 12204 15302
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 13938 12204 14350
rect 12268 13938 12296 14486
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12544 13870 12572 14282
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 13870 13400 14214
rect 13556 14006 13584 14758
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13544 14000 13596 14006
rect 13648 13977 13676 14214
rect 13544 13942 13596 13948
rect 13634 13968 13690 13977
rect 13634 13903 13690 13912
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12434 11836 13126
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 11808 12406 12020 12434
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11898 11008 12038
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 11060 11280 11112 11286
rect 11058 11248 11060 11257
rect 11112 11248 11114 11257
rect 11058 11183 11114 11192
rect 11164 11150 11192 11698
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10606 10916 10746
rect 11164 10742 11192 10950
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10600 10928 10606
rect 10980 10577 11008 10610
rect 10876 10542 10928 10548
rect 10966 10568 11022 10577
rect 10966 10503 10968 10512
rect 11020 10503 11022 10512
rect 10968 10474 11020 10480
rect 10980 10443 11008 10474
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 7546 11100 9930
rect 11256 9654 11284 10678
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11348 9178 11376 9590
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10874 6896 10930 6905
rect 10874 6831 10876 6840
rect 10928 6831 10930 6840
rect 10876 6802 10928 6808
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 5642 10824 6666
rect 10888 6458 10916 6802
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 4826 10824 5578
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 3126 11008 3538
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 11072 3058 11100 3878
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11164 2378 11192 3334
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11256 2310 11284 3878
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 2582 11376 3538
rect 11532 3466 11560 11018
rect 11624 4826 11652 11086
rect 11716 6458 11744 12174
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5234 11744 5714
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11808 3194 11836 7346
rect 11900 5302 11928 9522
rect 11992 7154 12020 12406
rect 12268 12322 12296 12718
rect 12544 12714 12572 13806
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 13266 13696 13322 13705
rect 12912 13326 12940 13670
rect 13266 13631 13322 13640
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 13161 12940 13262
rect 12898 13152 12954 13161
rect 12898 13087 12954 13096
rect 13174 12744 13230 12753
rect 12532 12708 12584 12714
rect 13174 12679 13230 12688
rect 12532 12650 12584 12656
rect 12176 12294 12296 12322
rect 12176 12186 12204 12294
rect 12084 12170 12204 12186
rect 12072 12164 12204 12170
rect 12124 12158 12204 12164
rect 12072 12106 12124 12112
rect 12176 11558 12204 12158
rect 12394 12164 12446 12170
rect 12394 12106 12446 12112
rect 12256 11756 12308 11762
rect 12406 11744 12434 12106
rect 12256 11698 12308 11704
rect 12360 11716 12434 11744
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10606 12204 11154
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 7274 12112 9522
rect 12176 8090 12204 9930
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12268 7970 12296 11698
rect 12360 11354 12388 11716
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 9518 12388 10950
rect 12544 10130 12572 12650
rect 13188 12646 13216 12679
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12636 11762 12664 12242
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12636 9994 12664 11086
rect 12728 10742 12756 12242
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10266 12848 11154
rect 12992 11144 13044 11150
rect 13044 11104 13216 11132
rect 12992 11086 13044 11092
rect 13188 11014 13216 11104
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12176 7942 12296 7970
rect 12176 7818 12204 7942
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12176 7206 12204 7754
rect 12254 7440 12310 7449
rect 12254 7375 12256 7384
rect 12308 7375 12310 7384
rect 12256 7346 12308 7352
rect 12164 7200 12216 7206
rect 11992 7126 12112 7154
rect 12164 7142 12216 7148
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11992 5778 12020 6122
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11888 5296 11940 5302
rect 11940 5256 12020 5284
rect 11888 5238 11940 5244
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4282 11928 4422
rect 11992 4282 12020 5256
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11900 3602 11928 4218
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12084 3233 12112 7126
rect 12360 5370 12388 8910
rect 12820 8838 12848 9454
rect 12912 9178 12940 10678
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9722 13124 9998
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8634 13032 8774
rect 13096 8634 13124 9386
rect 13280 8906 13308 13631
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13556 12850 13584 13398
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13464 12238 13492 12310
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13280 8090 13308 8842
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12440 6792 12492 6798
rect 12438 6760 12440 6769
rect 12492 6760 12494 6769
rect 12438 6695 12494 6704
rect 12544 6662 12572 7686
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 6186 13124 6598
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5302 12480 5510
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12532 4140 12584 4146
rect 12452 3738 12480 4111
rect 12532 4082 12584 4088
rect 12544 3890 12572 4082
rect 12714 4040 12770 4049
rect 12714 3975 12716 3984
rect 12768 3975 12770 3984
rect 12716 3946 12768 3952
rect 12544 3862 12756 3890
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12070 3224 12126 3233
rect 11796 3188 11848 3194
rect 12070 3159 12126 3168
rect 11796 3130 11848 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 10600 2032 10652 2038
rect 10600 1974 10652 1980
rect 11624 800 11652 2994
rect 11900 2854 11928 2994
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 12268 2582 12296 3402
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 12452 762 12480 2994
rect 12544 2990 12572 3402
rect 12636 3233 12664 3674
rect 12728 3602 12756 3862
rect 13188 3754 13216 7890
rect 13372 7478 13400 9998
rect 13464 9110 13492 10678
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7546 13492 7754
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13464 6118 13492 6394
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13280 4758 13308 5034
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13372 3913 13400 4150
rect 13358 3904 13414 3913
rect 13358 3839 13414 3848
rect 13188 3726 13308 3754
rect 13280 3670 13308 3726
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12622 3224 12678 3233
rect 12622 3159 12678 3168
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 13464 2378 13492 6054
rect 13556 4826 13584 12786
rect 13648 9518 13676 13806
rect 13740 13705 13768 14962
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13820 13728 13872 13734
rect 13726 13696 13782 13705
rect 13820 13670 13872 13676
rect 13726 13631 13782 13640
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13740 13462 13768 13495
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13832 13326 13860 13670
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13924 12782 13952 13874
rect 14016 12918 14044 14758
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14200 12866 14228 14554
rect 14292 13326 14320 16730
rect 14844 16658 14872 17070
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 14660 15706 14688 16118
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14752 15502 14780 15642
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14384 14550 14412 15030
rect 14568 15026 14596 15302
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 13410 14412 14486
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14476 14074 14504 14282
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14384 13382 14504 13410
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12986 14412 13126
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14200 12838 14412 12866
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 10554 13768 11562
rect 13818 11384 13874 11393
rect 13818 11319 13874 11328
rect 13832 11082 13860 11319
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 10656 13860 11018
rect 13912 10668 13964 10674
rect 13832 10628 13912 10656
rect 13912 10610 13964 10616
rect 13740 10538 13952 10554
rect 13740 10532 13964 10538
rect 13740 10526 13912 10532
rect 13912 10474 13964 10480
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9110 13768 9454
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13648 6866 13676 8502
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13740 7478 13768 8026
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13648 5817 13676 6190
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13648 5642 13676 5743
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13740 4554 13768 6326
rect 13832 5846 13860 9862
rect 13924 9382 13952 9930
rect 14016 9674 14044 12174
rect 14108 11830 14136 12650
rect 14200 12306 14228 12718
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14200 11626 14228 12242
rect 14292 12238 14320 12718
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14278 11248 14334 11257
rect 14278 11183 14334 11192
rect 14292 11150 14320 11183
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14186 10840 14242 10849
rect 14186 10775 14242 10784
rect 14016 9646 14136 9674
rect 14200 9654 14228 10775
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13648 3670 13676 4490
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 3194 13584 3402
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13740 3126 13768 3538
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13832 2990 13860 5782
rect 13924 5778 13952 9318
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14016 8498 14044 8978
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14108 8022 14136 9646
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 6866 14136 7278
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6458 14044 6666
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14188 5160 14240 5166
rect 14292 5137 14320 11086
rect 14384 9994 14412 12838
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14370 8936 14426 8945
rect 14476 8922 14504 13382
rect 14568 13138 14596 14962
rect 14660 13274 14688 15438
rect 14752 14618 14780 15438
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 15028 14482 15056 15574
rect 15120 15570 15148 15914
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15396 15094 15424 16934
rect 15488 15162 15516 17070
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13530 14964 14214
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14660 13246 14964 13274
rect 14568 13110 14872 13138
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14568 11132 14596 12174
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11286 14688 12038
rect 14752 11830 14780 12650
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14568 11104 14688 11132
rect 14554 9072 14610 9081
rect 14554 9007 14610 9016
rect 14568 8922 14596 9007
rect 14476 8906 14596 8922
rect 14476 8900 14608 8906
rect 14476 8894 14556 8900
rect 14370 8871 14426 8880
rect 14384 8838 14412 8871
rect 14556 8842 14608 8848
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 8090 14504 8230
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14660 7002 14688 11104
rect 14844 10713 14872 13110
rect 14830 10704 14886 10713
rect 14830 10639 14886 10648
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14752 9489 14780 9590
rect 14738 9480 14794 9489
rect 14738 9415 14794 9424
rect 14752 7313 14780 9415
rect 14738 7304 14794 7313
rect 14738 7239 14794 7248
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14738 6896 14794 6905
rect 14556 6860 14608 6866
rect 14844 6848 14872 10639
rect 14936 7342 14964 13246
rect 15028 10849 15056 14418
rect 15120 13258 15148 14758
rect 15212 14006 15240 14826
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15304 13818 15332 14962
rect 15580 14226 15608 16594
rect 15672 16046 15700 26726
rect 17696 22094 17724 33798
rect 18800 27130 18828 36654
rect 19352 30258 19380 36722
rect 19444 35834 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20548 36922 20576 37334
rect 20640 37330 20668 39200
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 20628 37324 20680 37330
rect 20628 37266 20680 37272
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 21284 36922 21312 37198
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 21272 36916 21324 36922
rect 21272 36858 21324 36864
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 17604 22066 17724 22094
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15672 15570 15700 15982
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15764 15162 15792 16118
rect 16040 15434 16068 16934
rect 16224 16658 16252 17138
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16132 16250 16160 16458
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 15936 15360 15988 15366
rect 16224 15348 16252 16594
rect 16592 16522 16620 16934
rect 17328 16590 17356 17138
rect 17604 16794 17632 22066
rect 18156 17542 18184 26250
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17066 18184 17478
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15936 15302 15988 15308
rect 16132 15320 16252 15348
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15212 13790 15332 13818
rect 15488 14198 15608 14226
rect 15488 13802 15516 14198
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15476 13796 15528 13802
rect 15212 13734 15240 13790
rect 15476 13738 15528 13744
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13394 15332 13670
rect 15488 13530 15516 13738
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15200 13184 15252 13190
rect 15198 13152 15200 13161
rect 15252 13152 15254 13161
rect 15198 13087 15254 13096
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15200 11144 15252 11150
rect 15304 11132 15332 12718
rect 15396 11354 15424 12854
rect 15488 12306 15516 13466
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15580 11898 15608 14010
rect 15672 13870 15700 14554
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15764 14362 15792 14486
rect 15948 14482 15976 15302
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15764 14334 15976 14362
rect 15948 14278 15976 14334
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15672 12782 15700 13194
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15764 12442 15792 13942
rect 16040 13326 16068 14962
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16132 13138 16160 15320
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16224 14657 16252 14962
rect 16316 14822 16344 15846
rect 16408 14890 16436 15982
rect 16592 15706 16620 16050
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16776 15638 16804 16458
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16868 15366 16896 15982
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16210 14648 16266 14657
rect 16210 14583 16266 14592
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 15948 13110 16160 13138
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15252 11104 15332 11132
rect 15200 11086 15252 11092
rect 15014 10840 15070 10849
rect 15014 10775 15070 10784
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 15028 10441 15056 10474
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15106 10024 15162 10033
rect 15106 9959 15108 9968
rect 15160 9959 15162 9968
rect 15108 9930 15160 9936
rect 15120 9625 15148 9930
rect 15200 9648 15252 9654
rect 15106 9616 15162 9625
rect 15200 9590 15252 9596
rect 15106 9551 15162 9560
rect 15212 9178 15240 9590
rect 15382 9480 15438 9489
rect 15382 9415 15438 9424
rect 15396 9382 15424 9415
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15106 9072 15162 9081
rect 15304 9058 15332 9114
rect 15162 9030 15332 9058
rect 15106 9007 15162 9016
rect 15106 8800 15162 8809
rect 15106 8735 15162 8744
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14794 6840 14872 6848
rect 14738 6831 14872 6840
rect 14556 6802 14608 6808
rect 14752 6820 14872 6831
rect 14462 6760 14518 6769
rect 14462 6695 14464 6704
rect 14516 6695 14518 6704
rect 14464 6666 14516 6672
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 5574 14412 6598
rect 14568 6254 14596 6802
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14568 5710 14596 6190
rect 14660 5914 14688 6190
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14188 5102 14240 5108
rect 14278 5128 14334 5137
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14108 4146 14136 4422
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3534 14136 4082
rect 14200 4078 14228 5102
rect 14278 5063 14280 5072
rect 14332 5063 14334 5072
rect 14280 5034 14332 5040
rect 14292 5003 14320 5034
rect 14278 4720 14334 4729
rect 14278 4655 14280 4664
rect 14332 4655 14334 4664
rect 14280 4626 14332 4632
rect 14384 4282 14412 5510
rect 14660 4826 14688 5850
rect 14752 5760 14780 6820
rect 14936 6746 14964 7278
rect 15028 6866 15056 7958
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14844 6730 14964 6746
rect 14832 6724 14964 6730
rect 14884 6718 14964 6724
rect 14832 6666 14884 6672
rect 14832 5772 14884 5778
rect 14752 5732 14832 5760
rect 14832 5714 14884 5720
rect 15014 5672 15070 5681
rect 15014 5607 15070 5616
rect 14738 5400 14794 5409
rect 14738 5335 14794 5344
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14568 4486 14596 4694
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14568 4078 14596 4422
rect 14752 4214 14780 5335
rect 15028 5302 15056 5607
rect 15016 5296 15068 5302
rect 15014 5264 15016 5273
rect 15068 5264 15070 5273
rect 15014 5199 15070 5208
rect 15120 5166 15148 8735
rect 15488 8430 15516 11698
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 10577 15608 11290
rect 15566 10568 15622 10577
rect 15566 10503 15622 10512
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7546 15240 7822
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15580 7274 15608 10503
rect 15672 9489 15700 12106
rect 15856 11914 15884 12378
rect 15764 11886 15884 11914
rect 15764 11354 15792 11886
rect 15844 11824 15896 11830
rect 15842 11792 15844 11801
rect 15896 11792 15898 11801
rect 15948 11762 15976 13110
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15842 11727 15898 11736
rect 15936 11756 15988 11762
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15856 11200 15884 11727
rect 15936 11698 15988 11704
rect 16040 11558 16068 12854
rect 16118 11792 16174 11801
rect 16118 11727 16174 11736
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15856 11172 15976 11200
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15672 8430 15700 8570
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15108 5160 15160 5166
rect 15384 5160 15436 5166
rect 15108 5102 15160 5108
rect 15382 5128 15384 5137
rect 15436 5128 15438 5137
rect 15382 5063 15438 5072
rect 15488 5030 15516 5238
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14844 4729 14872 4762
rect 14830 4720 14886 4729
rect 14830 4655 14886 4664
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 3058 14136 3470
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 14108 2514 14136 2994
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 14292 898 14320 3606
rect 15580 2774 15608 7210
rect 15764 6458 15792 11018
rect 15856 10538 15884 11018
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15856 7818 15884 9930
rect 15948 9674 15976 11172
rect 16040 11150 16068 11290
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 11014 16068 11086
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16132 10198 16160 11727
rect 16224 11354 16252 14418
rect 16316 13870 16344 14758
rect 16500 14634 16528 15098
rect 16408 14606 16528 14634
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 10192 16172 10198
rect 16316 10146 16344 13262
rect 16408 11762 16436 14606
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16500 14006 16528 14486
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16592 13569 16620 14282
rect 16578 13560 16634 13569
rect 16578 13495 16634 13504
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16486 12200 16542 12209
rect 16486 12135 16488 12144
rect 16540 12135 16542 12144
rect 16488 12106 16540 12112
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16500 11354 16528 12106
rect 16684 11694 16712 13330
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16120 10134 16172 10140
rect 16224 10118 16344 10146
rect 15948 9646 16068 9674
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 8945 15976 9318
rect 15934 8936 15990 8945
rect 15934 8871 15990 8880
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15856 6866 15884 7754
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5574 15792 6190
rect 15948 6186 15976 8774
rect 16040 7818 16068 9646
rect 16224 9586 16252 10118
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16316 9518 16344 9998
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16316 8974 16344 9454
rect 16408 9178 16436 11154
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16486 8936 16542 8945
rect 16316 8498 16344 8910
rect 16486 8871 16488 8880
rect 16540 8871 16542 8880
rect 16488 8842 16540 8848
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16316 7954 16344 8434
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16224 6322 16252 7754
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6934 16344 7346
rect 16408 7002 16436 7890
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15764 5234 15792 5510
rect 16040 5370 16068 6258
rect 16224 5681 16252 6258
rect 16316 5914 16344 6870
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16210 5672 16266 5681
rect 16210 5607 16266 5616
rect 16316 5370 16344 5850
rect 16408 5778 16436 6734
rect 16500 6458 16528 7414
rect 16592 6866 16620 10678
rect 16684 10198 16712 10950
rect 16776 10674 16804 12718
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 10441 16804 10610
rect 16762 10432 16818 10441
rect 16762 10367 16818 10376
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 8906 16712 9522
rect 16776 9518 16804 10367
rect 16868 9874 16896 15302
rect 17236 15094 17264 16390
rect 17328 15502 17356 16526
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 16960 14906 16988 15030
rect 17040 14952 17092 14958
rect 16960 14900 17040 14906
rect 16960 14894 17092 14900
rect 16960 14878 17080 14894
rect 17222 13968 17278 13977
rect 17222 13903 17278 13912
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13394 17080 13806
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17236 13258 17264 13903
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17040 12776 17092 12782
rect 17038 12744 17040 12753
rect 17092 12744 17094 12753
rect 17038 12679 17094 12688
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 10606 16988 11154
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16868 9846 16988 9874
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16776 8566 16804 8910
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 16040 4078 16068 5306
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16132 3126 16160 3538
rect 16408 3534 16436 5714
rect 16500 5642 16528 6122
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16396 3528 16448 3534
rect 16210 3496 16266 3505
rect 16396 3470 16448 3476
rect 16210 3431 16212 3440
rect 16264 3431 16266 3440
rect 16212 3402 16264 3408
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3194 16620 3334
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16120 3120 16172 3126
rect 16118 3088 16120 3097
rect 16172 3088 16174 3097
rect 16592 3058 16620 3130
rect 16118 3023 16174 3032
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 15580 2746 15884 2774
rect 15856 2514 15884 2746
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15290 2408 15346 2417
rect 15290 2343 15292 2352
rect 15344 2343 15346 2352
rect 15292 2314 15344 2320
rect 15304 1970 15332 2314
rect 16684 2310 16712 3130
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 12820 870 12940 898
rect 14292 870 14504 898
rect 12820 762 12848 870
rect 12912 800 12940 870
rect 12452 734 12848 762
rect 12898 200 12954 800
rect 14476 762 14504 870
rect 14752 870 14872 898
rect 14752 762 14780 870
rect 14844 800 14872 870
rect 16776 800 16804 3878
rect 16868 3466 16896 9658
rect 16960 9382 16988 9846
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17052 8090 17080 11766
rect 17144 9450 17172 11766
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17328 8838 17356 15438
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17512 14550 17540 14826
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17696 14482 17724 15574
rect 18248 15094 18276 15846
rect 18340 15586 18368 26726
rect 19352 18290 19380 29990
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20548 26926 20576 36858
rect 21836 36786 21864 37606
rect 21928 37210 21956 39200
rect 23020 37460 23072 37466
rect 23020 37402 23072 37408
rect 21928 37182 22140 37210
rect 22112 37126 22140 37182
rect 22100 37120 22152 37126
rect 22100 37062 22152 37068
rect 23032 36854 23060 37402
rect 23860 37126 23888 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 23020 36848 23072 36854
rect 23020 36790 23072 36796
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 22020 26586 22048 36722
rect 23032 27606 23060 36790
rect 24596 29306 24624 37198
rect 25148 37126 25176 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 22008 26580 22060 26586
rect 22008 26522 22060 26528
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17882 19288 18022
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19260 17270 19288 17818
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18432 16114 18460 16458
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18340 15570 18460 15586
rect 18328 15564 18460 15570
rect 18380 15558 18460 15564
rect 18328 15506 18380 15512
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18340 14618 18368 15370
rect 18432 14958 18460 15558
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18524 14618 18552 14826
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17696 14006 17724 14418
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12306 17724 12854
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17788 11914 17816 13126
rect 17696 11898 17816 11914
rect 17684 11892 17816 11898
rect 17736 11886 17816 11892
rect 17684 11834 17736 11840
rect 17880 11830 17908 14554
rect 18616 14074 18644 17206
rect 19260 16998 19288 17206
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19352 15162 19380 18090
rect 19444 17746 19472 18294
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19524 17672 19576 17678
rect 19444 17620 19524 17626
rect 19444 17614 19576 17620
rect 19444 17598 19564 17614
rect 19444 16794 19472 17598
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20088 16182 20116 26250
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19444 16046 19472 16118
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19444 15638 19472 15982
rect 19536 15706 19564 15982
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17868 11688 17920 11694
rect 17866 11656 17868 11665
rect 17920 11656 17922 11665
rect 17866 11591 17922 11600
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17420 10470 17448 10678
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 8832 17368 8838
rect 17368 8792 17448 8820
rect 17316 8774 17368 8780
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17328 7342 17356 8026
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17420 7002 17448 8792
rect 17604 8294 17632 11018
rect 17880 9518 17908 11591
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 18064 9382 18092 13874
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18432 12238 18460 13194
rect 18800 12918 18828 14214
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18248 11393 18276 12106
rect 18234 11384 18290 11393
rect 18234 11319 18290 11328
rect 18326 10840 18382 10849
rect 18326 10775 18382 10784
rect 18340 10606 18368 10775
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18432 9674 18460 12174
rect 18616 12102 18644 12854
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11286 18644 12038
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 19076 11218 19104 14758
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18892 10198 18920 10406
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18340 9646 18460 9674
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 17960 8832 18012 8838
rect 18156 8809 18184 9046
rect 17960 8774 18012 8780
rect 18142 8800 18198 8809
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17316 6724 17368 6730
rect 17316 6666 17368 6672
rect 17328 6118 17356 6666
rect 17604 6361 17632 7754
rect 17696 7478 17724 8230
rect 17880 7954 17908 8502
rect 17972 8430 18000 8774
rect 18142 8735 18198 8744
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17868 6384 17920 6390
rect 17590 6352 17646 6361
rect 17868 6326 17920 6332
rect 17590 6287 17646 6296
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17420 5914 17448 6122
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5234 17172 5714
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17132 5228 17184 5234
rect 17052 5188 17132 5216
rect 17052 4690 17080 5188
rect 17132 5170 17184 5176
rect 17328 4865 17356 5306
rect 17314 4856 17370 4865
rect 17314 4791 17370 4800
rect 17328 4690 17356 4791
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17052 4146 17080 4626
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 2582 16896 3402
rect 17052 3398 17080 4082
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17236 3126 17264 3674
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17420 2774 17448 5850
rect 17880 5137 17908 6326
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 18340 4826 18368 9646
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 8634 18644 9318
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18892 7886 18920 9862
rect 18984 8294 19012 9998
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18432 4842 18460 7278
rect 18524 7002 18552 7346
rect 18616 7206 18644 7754
rect 18984 7478 19012 7958
rect 19076 7546 19104 10678
rect 19168 8634 19196 14962
rect 19444 14498 19472 15574
rect 19628 15434 19656 15846
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19352 14470 19472 14498
rect 19904 14482 19932 14962
rect 19892 14476 19944 14482
rect 19352 14090 19380 14470
rect 19892 14418 19944 14424
rect 19996 14346 20024 16050
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19260 14062 19380 14090
rect 19260 13394 19288 14062
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19352 12442 19380 13942
rect 19444 13870 19472 14282
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19798 13696 19854 13705
rect 19798 13631 19854 13640
rect 19812 13326 19840 13631
rect 20180 13394 20208 18022
rect 20272 16114 20300 20198
rect 21652 17882 21680 24754
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21652 17202 21680 17818
rect 22112 17746 22140 27270
rect 25240 24410 25268 37130
rect 25332 36718 25360 37198
rect 27080 37126 27108 39200
rect 29012 37126 29040 39200
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 30300 37210 30328 39200
rect 30748 37256 30800 37262
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 25320 36712 25372 36718
rect 25320 36654 25372 36660
rect 25228 24404 25280 24410
rect 25228 24346 25280 24352
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 22112 17134 22140 17682
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23124 17338 23152 17478
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20272 14482 20300 16050
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20732 15162 20760 15982
rect 20824 15706 20852 17070
rect 21732 17060 21784 17066
rect 21732 17002 21784 17008
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 21284 15434 21312 16458
rect 21468 15502 21496 16934
rect 21744 16522 21772 17002
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21928 15722 21956 16458
rect 22112 16114 22140 16594
rect 22192 16448 22244 16454
rect 22296 16402 22324 17206
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16658 22416 16934
rect 23124 16658 23152 17002
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 22244 16396 22324 16402
rect 22192 16390 22324 16396
rect 22204 16374 22324 16390
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 21836 15706 21956 15722
rect 22020 15706 22048 15846
rect 21824 15700 21956 15706
rect 21876 15694 21956 15700
rect 22008 15700 22060 15706
rect 21824 15642 21876 15648
rect 22008 15642 22060 15648
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 13938 20300 14418
rect 20824 14414 20852 15030
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20640 13530 20668 13806
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20180 12918 20208 13330
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 20088 12209 20116 12854
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20074 12200 20130 12209
rect 20074 12135 20130 12144
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20088 11354 20116 11630
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10792 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20088 10810 20116 11154
rect 20076 10804 20128 10810
rect 19444 10764 19932 10792
rect 19430 10568 19486 10577
rect 19430 10503 19486 10512
rect 19338 10296 19394 10305
rect 19444 10266 19472 10503
rect 19338 10231 19394 10240
rect 19432 10260 19484 10266
rect 19246 10160 19302 10169
rect 19352 10146 19380 10231
rect 19432 10202 19484 10208
rect 19352 10118 19472 10146
rect 19246 10095 19302 10104
rect 19260 9994 19288 10095
rect 19444 10062 19472 10118
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19340 9988 19392 9994
rect 19628 9982 19748 10010
rect 19904 9994 19932 10764
rect 20076 10746 20128 10752
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19628 9976 19656 9982
rect 19340 9930 19392 9936
rect 19536 9948 19656 9976
rect 19352 9897 19380 9930
rect 19432 9920 19484 9926
rect 19338 9888 19394 9897
rect 19536 9908 19564 9948
rect 19720 9926 19748 9982
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19484 9880 19564 9908
rect 19708 9920 19760 9926
rect 19432 9862 19484 9868
rect 19708 9862 19760 9868
rect 19338 9823 19394 9832
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19338 9752 19394 9761
rect 19574 9755 19882 9764
rect 19338 9687 19394 9696
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 8294 19196 8570
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18708 7206 18736 7346
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18892 5846 18920 7414
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 6254 19012 6598
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19352 5914 19380 9687
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8566 19472 8978
rect 19628 8906 19656 9454
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19720 8906 19748 9114
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19444 7206 19472 7890
rect 19812 7750 19840 7890
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19444 6866 19472 7142
rect 19536 7002 19564 7142
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6390 19472 6802
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6384 19484 6390
rect 19800 6384 19852 6390
rect 19484 6344 19564 6372
rect 19432 6326 19484 6332
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18328 4820 18380 4826
rect 18432 4814 18552 4842
rect 18328 4762 18380 4768
rect 17868 4072 17920 4078
rect 17866 4040 17868 4049
rect 17920 4040 17922 4049
rect 17866 3975 17922 3984
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 17328 2746 17448 2774
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17328 2514 17356 2746
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 17880 1873 17908 2314
rect 17866 1864 17922 1873
rect 18156 1850 18184 3606
rect 18340 3380 18368 4762
rect 18524 4758 18552 4814
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18420 3392 18472 3398
rect 18340 3352 18420 3380
rect 18420 3334 18472 3340
rect 18892 2990 18920 5782
rect 19536 5778 19564 6344
rect 19996 6372 20024 9998
rect 20088 9722 20116 10542
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20088 9110 20116 9658
rect 20180 9518 20208 12718
rect 20732 12442 20760 13194
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21008 12374 21036 12718
rect 21192 12714 21220 13670
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20180 6633 20208 8298
rect 20272 7002 20300 10406
rect 20364 7750 20392 12174
rect 20824 12073 20852 12174
rect 20810 12064 20866 12073
rect 20810 11999 20866 12008
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20456 10062 20484 10474
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20548 9674 20576 10542
rect 20640 9761 20668 11018
rect 20626 9752 20682 9761
rect 20626 9687 20682 9696
rect 20456 9646 20576 9674
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20166 6624 20222 6633
rect 20166 6559 20222 6568
rect 19852 6344 20024 6372
rect 19800 6326 19852 6332
rect 19524 5772 19576 5778
rect 19444 5732 19524 5760
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18880 2984 18932 2990
rect 18984 2961 19012 4082
rect 18880 2926 18932 2932
rect 18970 2952 19026 2961
rect 19076 2922 19104 5646
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19260 5098 19288 5238
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19352 5001 19380 5578
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19260 4146 19288 4218
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19168 3913 19196 3946
rect 19154 3904 19210 3913
rect 19154 3839 19210 3848
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 18970 2887 19026 2896
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19076 2378 19104 2858
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 19168 2009 19196 3062
rect 19352 2378 19380 4694
rect 19444 4690 19472 5732
rect 19524 5714 19576 5720
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19892 5364 19944 5370
rect 19996 5352 20024 6344
rect 19944 5324 20024 5352
rect 19892 5306 19944 5312
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19812 4690 19840 5170
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19996 4729 20024 5034
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19982 4720 20038 4729
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19800 4684 19852 4690
rect 19982 4655 20038 4664
rect 19800 4626 19852 4632
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19996 3466 20024 3878
rect 20088 3466 20116 4966
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3194 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 20076 3120 20128 3126
rect 20180 3108 20208 6559
rect 20258 5672 20314 5681
rect 20258 5607 20260 5616
rect 20312 5607 20314 5616
rect 20260 5578 20312 5584
rect 20456 4185 20484 9646
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 8974 20576 9454
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20824 8906 20852 11999
rect 20916 11150 20944 12242
rect 21192 11898 21220 12650
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20994 10704 21050 10713
rect 20994 10639 20996 10648
rect 21048 10639 21050 10648
rect 20996 10610 21048 10616
rect 21100 9518 21128 11766
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21192 9382 21220 11290
rect 21284 11218 21312 15370
rect 21468 14006 21496 15438
rect 22020 15162 22048 15642
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21560 14890 21588 15098
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21546 14648 21602 14657
rect 21546 14583 21602 14592
rect 21560 14550 21588 14583
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21270 10568 21326 10577
rect 21270 10503 21326 10512
rect 21284 9994 21312 10503
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8673 20760 8774
rect 20718 8664 20774 8673
rect 21008 8634 21036 8910
rect 20718 8599 20774 8608
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20548 7585 20576 8026
rect 20534 7576 20590 7585
rect 20534 7511 20590 7520
rect 20548 7410 20576 7511
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20640 6905 20668 8502
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 7041 20760 7890
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20916 7177 20944 7482
rect 21088 7200 21140 7206
rect 20902 7168 20958 7177
rect 21088 7142 21140 7148
rect 20902 7103 20958 7112
rect 20718 7032 20774 7041
rect 20718 6967 20774 6976
rect 20626 6896 20682 6905
rect 20626 6831 20682 6840
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 5953 20760 6598
rect 20718 5944 20774 5953
rect 20718 5879 20774 5888
rect 20442 4176 20498 4185
rect 20442 4111 20498 4120
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 4010 20760 4082
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20128 3080 20208 3108
rect 20076 3062 20128 3068
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 2514 19472 2994
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19892 2508 19944 2514
rect 19944 2468 20024 2496
rect 19892 2450 19944 2456
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19154 2000 19210 2009
rect 19154 1935 19210 1944
rect 17866 1799 17922 1808
rect 18064 1822 18184 1850
rect 18064 800 18092 1822
rect 19996 800 20024 2468
rect 20548 1834 20576 3402
rect 20732 3398 20760 3946
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20626 2816 20682 2825
rect 20626 2751 20682 2760
rect 21100 2774 21128 7142
rect 21192 6662 21220 9318
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21284 7002 21312 8502
rect 21376 7546 21404 13194
rect 21468 12850 21496 13942
rect 21560 13802 21588 14282
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21732 13456 21784 13462
rect 21732 13398 21784 13404
rect 21744 13326 21772 13398
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21560 10810 21588 12106
rect 21652 11558 21680 12106
rect 21744 11830 21772 13126
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21836 12170 21864 12718
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21744 11218 21772 11766
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21824 11008 21876 11014
rect 21824 10950 21876 10956
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21836 10538 21864 10950
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21928 10538 21956 10610
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 22112 10266 22140 16050
rect 23216 16046 23244 17614
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23676 17134 23704 17546
rect 23952 17270 23980 17750
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23676 16726 23704 17070
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23308 16250 23336 16526
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23204 16040 23256 16046
rect 23952 15994 23980 17206
rect 24596 16998 24624 17614
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24780 16250 24808 17614
rect 24872 16250 24900 18158
rect 24964 17338 24992 24142
rect 25332 22094 25360 36654
rect 29748 36582 29776 37198
rect 30300 37182 30420 37210
rect 30748 37198 30800 37204
rect 30392 37126 30420 37182
rect 30656 37188 30708 37194
rect 30656 37130 30708 37136
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 29736 36576 29788 36582
rect 29736 36518 29788 36524
rect 27896 35488 27948 35494
rect 27896 35430 27948 35436
rect 26148 33312 26200 33318
rect 26148 33254 26200 33260
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25516 24886 25544 32710
rect 25504 24880 25556 24886
rect 25504 24822 25556 24828
rect 25056 22066 25360 22094
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24964 16794 24992 17274
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 16289 24992 16458
rect 24950 16280 25006 16289
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24860 16244 24912 16250
rect 24950 16215 25006 16224
rect 24860 16186 24912 16192
rect 25056 16130 25084 22066
rect 26160 18970 26188 33254
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26160 18766 26188 18906
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25148 17542 25176 18022
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25148 16658 25176 17478
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25148 16504 25176 16594
rect 25228 16516 25280 16522
rect 25148 16476 25228 16504
rect 25228 16458 25280 16464
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24872 16102 25084 16130
rect 23204 15982 23256 15988
rect 23860 15966 23980 15994
rect 23860 15706 23888 15966
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23952 15638 23980 15846
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23940 15632 23992 15638
rect 23940 15574 23992 15580
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22204 13734 22232 13942
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22296 13258 22324 15030
rect 22756 14958 22784 15438
rect 23492 15162 23520 15574
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 23020 14340 23072 14346
rect 23020 14282 23072 14288
rect 22388 14006 22416 14282
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 23032 13530 23060 14282
rect 23124 14006 23152 14894
rect 23216 14482 23244 14894
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23216 13394 23244 14418
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22296 12434 22324 12854
rect 22296 12406 22416 12434
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22204 11064 22232 11222
rect 22388 11200 22416 12406
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22468 11688 22520 11694
rect 22466 11656 22468 11665
rect 22520 11656 22522 11665
rect 22466 11591 22522 11600
rect 22468 11212 22520 11218
rect 22388 11172 22468 11200
rect 22468 11154 22520 11160
rect 22468 11076 22520 11082
rect 22204 11036 22468 11064
rect 22468 11018 22520 11024
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 7886 21496 8434
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21454 7712 21510 7721
rect 21454 7647 21510 7656
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21376 6254 21404 7346
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21192 4214 21220 4694
rect 21180 4208 21232 4214
rect 21180 4150 21232 4156
rect 21376 4078 21404 6190
rect 21468 4758 21496 7647
rect 21560 7274 21588 9658
rect 22112 9518 22140 10202
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22204 9722 22232 9930
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22204 8838 22232 9522
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22296 8650 22324 9046
rect 22112 8622 22324 8650
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21928 7478 21956 8298
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 22020 7342 22048 7822
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 22020 6254 22048 7278
rect 22008 6248 22060 6254
rect 21822 6216 21878 6225
rect 22008 6190 22060 6196
rect 21822 6151 21878 6160
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21744 5642 21772 6054
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21836 5098 21864 6151
rect 22020 5710 22048 6190
rect 22112 5930 22140 8622
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 6089 22232 7686
rect 22296 7478 22324 8230
rect 22374 7576 22430 7585
rect 22374 7511 22376 7520
rect 22428 7511 22430 7520
rect 22376 7482 22428 7488
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22282 6896 22338 6905
rect 22282 6831 22338 6840
rect 22296 6662 22324 6831
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22282 6488 22338 6497
rect 22282 6423 22338 6432
rect 22296 6390 22324 6423
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22388 6254 22416 7142
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 22190 6080 22246 6089
rect 22190 6015 22246 6024
rect 22296 5930 22324 6190
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22112 5902 22324 5930
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21744 3738 21772 3878
rect 21928 3777 21956 5510
rect 22020 5148 22048 5646
rect 22388 5166 22416 6054
rect 22100 5160 22152 5166
rect 22020 5120 22100 5148
rect 22376 5160 22428 5166
rect 22152 5120 22232 5148
rect 22100 5102 22152 5108
rect 22204 4554 22232 5120
rect 22376 5102 22428 5108
rect 22480 5030 22508 11018
rect 22572 5778 22600 11766
rect 22664 10742 22692 12242
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22652 10736 22704 10742
rect 22652 10678 22704 10684
rect 22664 10130 22692 10678
rect 22756 10606 22784 11562
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22756 10198 22784 10542
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 23124 9110 23152 11154
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 22848 6730 22876 7890
rect 23216 7154 23244 10610
rect 23400 9178 23428 14214
rect 23492 9654 23520 15098
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 12442 23796 12718
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23754 12200 23810 12209
rect 23754 12135 23810 12144
rect 23768 11218 23796 12135
rect 23860 11762 23888 13398
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23952 11898 23980 12718
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 12073 24072 12174
rect 24030 12064 24086 12073
rect 24030 11999 24086 12008
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23848 11756 23900 11762
rect 23900 11716 24072 11744
rect 23848 11698 23900 11704
rect 23848 11620 23900 11626
rect 23848 11562 23900 11568
rect 23860 11354 23888 11562
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 24044 11234 24072 11716
rect 24136 11354 24164 15030
rect 24504 14822 24532 16050
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24688 14482 24716 15370
rect 24780 15162 24808 16050
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 23756 11212 23808 11218
rect 24044 11206 24164 11234
rect 23756 11154 23808 11160
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10810 23612 11086
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23492 7562 23520 9590
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23676 8090 23704 8910
rect 23754 8800 23810 8809
rect 23754 8735 23810 8744
rect 23768 8566 23796 8735
rect 23860 8566 23888 9454
rect 23952 9178 23980 10474
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23860 8412 23888 8502
rect 23768 8384 23888 8412
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23676 7750 23704 8026
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23492 7546 23704 7562
rect 23492 7540 23716 7546
rect 23492 7534 23664 7540
rect 23664 7482 23716 7488
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23400 7206 23428 7346
rect 23480 7268 23532 7274
rect 23480 7210 23532 7216
rect 22940 7126 23244 7154
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 22836 6724 22888 6730
rect 22836 6666 22888 6672
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22664 5658 22692 5714
rect 22572 5630 22692 5658
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22572 4554 22600 5630
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22664 4593 22692 5238
rect 22650 4584 22706 4593
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 22284 4548 22336 4554
rect 22284 4490 22336 4496
rect 22560 4548 22612 4554
rect 22650 4519 22706 4528
rect 22560 4490 22612 4496
rect 22204 4214 22232 4490
rect 22296 4282 22324 4490
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22374 4176 22430 4185
rect 22006 4040 22062 4049
rect 22006 3975 22008 3984
rect 22060 3975 22062 3984
rect 22008 3946 22060 3952
rect 21914 3768 21970 3777
rect 21732 3732 21784 3738
rect 21732 3674 21784 3680
rect 21824 3732 21876 3738
rect 21914 3703 21970 3712
rect 21824 3674 21876 3680
rect 21836 3466 21864 3674
rect 22204 3602 22232 4150
rect 22374 4111 22430 4120
rect 22388 4078 22416 4111
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 20640 2310 20668 2751
rect 21100 2746 21220 2774
rect 21192 2582 21220 2746
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20536 1828 20588 1834
rect 20536 1770 20588 1776
rect 21284 800 21312 3334
rect 22098 3224 22154 3233
rect 22098 3159 22154 3168
rect 22112 2938 22140 3159
rect 22204 3126 22232 3538
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 21928 2910 22140 2938
rect 21928 2854 21956 2910
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 22100 2508 22152 2514
rect 22204 2496 22232 3062
rect 22296 2990 22324 3062
rect 22388 2990 22416 3402
rect 22940 3194 22968 7126
rect 23492 6984 23520 7210
rect 23216 6956 23520 6984
rect 23216 6730 23244 6956
rect 23294 6896 23350 6905
rect 23768 6866 23796 8384
rect 24044 8090 24072 10542
rect 24136 8566 24164 11206
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23294 6831 23296 6840
rect 23348 6831 23350 6840
rect 23756 6860 23808 6866
rect 23296 6802 23348 6808
rect 23756 6802 23808 6808
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23204 6724 23256 6730
rect 23204 6666 23256 6672
rect 23478 6216 23534 6225
rect 23478 6151 23480 6160
rect 23532 6151 23534 6160
rect 23480 6122 23532 6128
rect 23676 6118 23704 6734
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23860 5370 23888 7210
rect 23952 5370 23980 7890
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24044 6118 24072 6394
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24136 5930 24164 8502
rect 24228 7546 24256 13670
rect 24320 12374 24348 13738
rect 24412 13462 24440 13806
rect 24400 13456 24452 13462
rect 24400 13398 24452 13404
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24504 13190 24532 13262
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24308 12368 24360 12374
rect 24308 12310 24360 12316
rect 24320 12170 24348 12310
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24228 6322 24256 6802
rect 24412 6730 24440 13126
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24504 11218 24532 11290
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24504 10674 24532 11154
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24596 10266 24624 13194
rect 24688 12986 24716 13806
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 11354 24716 12582
rect 24872 12434 24900 16102
rect 25608 15570 25636 18566
rect 25700 17882 25728 18702
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25596 15564 25648 15570
rect 25596 15506 25648 15512
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25056 15162 25084 15438
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 24780 12406 24900 12434
rect 24780 11830 24808 12406
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24596 9722 24624 10202
rect 24780 10130 24808 10746
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24596 8906 24624 9318
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24504 8362 24532 8842
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24044 5902 24164 5930
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 23032 3942 23060 5102
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4622 23612 4966
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23020 3936 23072 3942
rect 23676 3913 23704 4422
rect 23020 3878 23072 3884
rect 23662 3904 23718 3913
rect 23662 3839 23718 3848
rect 23768 3754 23796 4422
rect 23584 3726 23796 3754
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22152 2468 22232 2496
rect 22100 2450 22152 2456
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22296 1902 22324 2314
rect 22284 1896 22336 1902
rect 22284 1838 22336 1844
rect 23216 800 23244 3334
rect 23584 2774 23612 3726
rect 24044 3233 24072 5902
rect 24228 5710 24256 6258
rect 24596 6236 24624 8842
rect 24688 7002 24716 9590
rect 24766 9208 24822 9217
rect 24766 9143 24822 9152
rect 24780 8566 24808 9143
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24766 8120 24822 8129
rect 24872 8090 24900 10678
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24964 9518 24992 9590
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24766 8055 24822 8064
rect 24860 8084 24912 8090
rect 24780 7886 24808 8055
rect 24860 8026 24912 8032
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24780 7274 24808 7822
rect 25056 7546 25084 13942
rect 25148 13394 25176 15438
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25240 14482 25268 14894
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25148 12986 25176 13194
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25332 12374 25360 15506
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25700 12442 25728 12718
rect 25688 12436 25740 12442
rect 25688 12378 25740 12384
rect 25320 12368 25372 12374
rect 25320 12310 25372 12316
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25332 11529 25360 11630
rect 25318 11520 25374 11529
rect 25318 11455 25374 11464
rect 25424 11354 25452 12038
rect 25516 11762 25544 12038
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25884 11694 25912 17070
rect 26332 14408 26384 14414
rect 26332 14350 26384 14356
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 25976 12850 26004 14214
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 26068 12714 26096 13194
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 26068 12442 26096 12650
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26068 11898 26096 12378
rect 26160 12322 26188 13330
rect 26160 12294 26280 12322
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 26252 11558 26280 12294
rect 26344 12209 26372 14350
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26436 12374 26464 13466
rect 26620 12918 26648 14214
rect 26608 12912 26660 12918
rect 26608 12854 26660 12860
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26608 12232 26660 12238
rect 26330 12200 26386 12209
rect 26608 12174 26660 12180
rect 26330 12135 26386 12144
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25148 10742 25176 10950
rect 25240 10810 25268 10950
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 25516 10674 25544 10950
rect 25792 10674 25820 11086
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24768 7268 24820 7274
rect 24768 7210 24820 7216
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24768 6860 24820 6866
rect 24412 6208 24624 6236
rect 24688 6820 24768 6848
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24306 4856 24362 4865
rect 24306 4791 24362 4800
rect 24320 4486 24348 4791
rect 24308 4480 24360 4486
rect 24122 4448 24178 4457
rect 24308 4422 24360 4428
rect 24122 4383 24178 4392
rect 24136 4214 24164 4383
rect 24412 4298 24440 6208
rect 24584 5704 24636 5710
rect 24688 5692 24716 6820
rect 24768 6802 24820 6808
rect 24636 5664 24716 5692
rect 24584 5646 24636 5652
rect 24492 5636 24544 5642
rect 24492 5578 24544 5584
rect 24504 4758 24532 5578
rect 24596 5030 24624 5646
rect 24872 5642 24900 7346
rect 24964 6225 24992 7346
rect 25332 6798 25360 10542
rect 25884 10305 25912 11086
rect 26344 10470 26372 11698
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 25870 10296 25926 10305
rect 26436 10266 26464 10542
rect 25870 10231 25926 10240
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26240 10192 26292 10198
rect 26240 10134 26292 10140
rect 26252 10062 26280 10134
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25410 7984 25466 7993
rect 25410 7919 25466 7928
rect 25424 7886 25452 7919
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 24950 6216 25006 6225
rect 24950 6151 25006 6160
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24492 4752 24544 4758
rect 24492 4694 24544 4700
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24320 4270 24440 4298
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24030 3224 24086 3233
rect 24030 3159 24086 3168
rect 24136 2922 24164 4014
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 3194 24256 3402
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24124 2916 24176 2922
rect 24124 2858 24176 2864
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23492 2746 23612 2774
rect 23388 2508 23440 2514
rect 23492 2496 23520 2746
rect 23440 2468 23520 2496
rect 23388 2450 23440 2456
rect 23676 2281 23704 2790
rect 23662 2272 23718 2281
rect 23662 2207 23718 2216
rect 24320 1834 24348 4270
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24412 2553 24440 3062
rect 24504 2938 24532 4422
rect 24596 4214 24624 4966
rect 24688 4321 24716 5170
rect 24674 4312 24730 4321
rect 24872 4282 24900 5578
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24674 4247 24730 4256
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24584 4208 24636 4214
rect 24584 4150 24636 4156
rect 24596 3534 24624 4150
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24584 3528 24636 3534
rect 24636 3488 24716 3516
rect 24584 3470 24636 3476
rect 24688 3194 24716 3488
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24504 2910 24624 2938
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 24398 2544 24454 2553
rect 24504 2514 24532 2790
rect 24398 2479 24454 2488
rect 24492 2508 24544 2514
rect 24492 2450 24544 2456
rect 24596 2106 24624 2910
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 24964 2038 24992 3538
rect 25056 2854 25084 4422
rect 25228 3596 25280 3602
rect 25228 3538 25280 3544
rect 25240 3482 25268 3538
rect 25148 3466 25268 3482
rect 25136 3460 25268 3466
rect 25188 3454 25268 3460
rect 25136 3402 25188 3408
rect 25332 2990 25360 4966
rect 25424 3233 25452 7414
rect 25516 6769 25544 8842
rect 25608 8090 25636 8910
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25700 7954 25728 9930
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25688 7948 25740 7954
rect 25688 7890 25740 7896
rect 25502 6760 25558 6769
rect 25502 6695 25558 6704
rect 25792 5817 25820 8570
rect 25884 7478 25912 9522
rect 26160 9178 26188 9930
rect 26240 9512 26292 9518
rect 26424 9512 26476 9518
rect 26292 9472 26372 9500
rect 26240 9454 26292 9460
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26146 9072 26202 9081
rect 26146 9007 26202 9016
rect 26160 8974 26188 9007
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26252 8634 26280 9114
rect 26240 8628 26292 8634
rect 26344 8616 26372 9472
rect 26424 9454 26476 9460
rect 26436 8906 26464 9454
rect 26528 9353 26556 11086
rect 26620 10606 26648 12174
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26712 9674 26740 24822
rect 27908 20058 27936 35430
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 27896 20052 27948 20058
rect 27896 19994 27948 20000
rect 27250 16280 27306 16289
rect 27250 16215 27306 16224
rect 27160 14884 27212 14890
rect 27160 14826 27212 14832
rect 27172 13938 27200 14826
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27172 12850 27200 13874
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 26804 12374 26832 12786
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26792 12368 26844 12374
rect 26792 12310 26844 12316
rect 27080 12238 27108 12718
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 26804 10130 26832 10406
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26712 9646 26832 9674
rect 26608 9512 26660 9518
rect 26606 9480 26608 9489
rect 26660 9480 26662 9489
rect 26606 9415 26662 9424
rect 26514 9344 26570 9353
rect 26514 9279 26570 9288
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26424 8628 26476 8634
rect 26344 8588 26424 8616
rect 26240 8570 26292 8576
rect 26424 8570 26476 8576
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26148 8424 26200 8430
rect 26148 8366 26200 8372
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 25976 6118 26004 7754
rect 26160 7342 26188 8366
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26160 6730 26188 7278
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 26252 6322 26280 8434
rect 26606 8256 26662 8265
rect 26606 8191 26662 8200
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 25778 5808 25834 5817
rect 25778 5743 25834 5752
rect 25870 5400 25926 5409
rect 25688 5364 25740 5370
rect 25870 5335 25926 5344
rect 25688 5306 25740 5312
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 25410 3224 25466 3233
rect 25410 3159 25466 3168
rect 25516 3108 25544 4218
rect 25700 3398 25728 5306
rect 25884 5234 25912 5335
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25516 3080 25636 3108
rect 25608 2990 25636 3080
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25056 2514 25084 2790
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24952 2032 25004 2038
rect 24952 1974 25004 1980
rect 24308 1828 24360 1834
rect 24308 1770 24360 1776
rect 25148 800 25176 2246
rect 25792 1970 25820 4558
rect 25976 3942 26004 6054
rect 26068 4622 26096 6054
rect 26344 5914 26372 7686
rect 26424 6724 26476 6730
rect 26424 6666 26476 6672
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26436 5914 26464 6666
rect 26528 6118 26556 6666
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26424 5908 26476 5914
rect 26424 5850 26476 5856
rect 26620 5846 26648 8191
rect 26712 6798 26740 8910
rect 26804 8498 26832 9646
rect 26896 9586 26924 12174
rect 27264 11898 27292 16215
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27344 13252 27396 13258
rect 27344 13194 27396 13200
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27252 11620 27304 11626
rect 27252 11562 27304 11568
rect 27264 11529 27292 11562
rect 27250 11520 27306 11529
rect 27250 11455 27306 11464
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26790 8256 26846 8265
rect 26790 8191 26846 8200
rect 26804 7954 26832 8191
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26790 6896 26846 6905
rect 26790 6831 26846 6840
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26712 6225 26740 6258
rect 26698 6216 26754 6225
rect 26698 6151 26754 6160
rect 26804 6118 26832 6831
rect 26896 6390 26924 8910
rect 26884 6384 26936 6390
rect 26884 6326 26936 6332
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 26988 5846 27016 11018
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 27080 9994 27108 10474
rect 27264 10470 27292 11455
rect 27356 10470 27384 13194
rect 27540 12986 27568 13942
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 28000 12850 28028 13670
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27540 12442 27568 12650
rect 27528 12436 27580 12442
rect 28000 12434 28028 12786
rect 27528 12378 27580 12384
rect 27908 12406 28028 12434
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 27448 11898 27476 12242
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27540 12073 27568 12174
rect 27526 12064 27582 12073
rect 27526 11999 27582 12008
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27448 11558 27476 11630
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27068 9988 27120 9994
rect 27068 9930 27120 9936
rect 27068 8832 27120 8838
rect 27068 8774 27120 8780
rect 27080 7954 27108 8774
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27066 7848 27122 7857
rect 27066 7783 27068 7792
rect 27120 7783 27122 7792
rect 27068 7754 27120 7760
rect 27172 7478 27200 10066
rect 27252 9716 27304 9722
rect 27540 9674 27568 11999
rect 27252 9658 27304 9664
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 27172 7002 27200 7414
rect 27264 7392 27292 9658
rect 27448 9646 27568 9674
rect 27632 9982 27844 10010
rect 27632 9654 27660 9982
rect 27712 9920 27764 9926
rect 27712 9862 27764 9868
rect 27620 9648 27672 9654
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27356 9058 27384 9386
rect 27448 9178 27476 9646
rect 27620 9590 27672 9596
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27540 9178 27568 9318
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27356 9030 27476 9058
rect 27448 8242 27476 9030
rect 27526 8528 27582 8537
rect 27526 8463 27528 8472
rect 27580 8463 27582 8472
rect 27528 8434 27580 8440
rect 27632 8430 27660 9454
rect 27724 9450 27752 9862
rect 27816 9518 27844 9982
rect 27908 9738 27936 12406
rect 28172 12368 28224 12374
rect 28172 12310 28224 12316
rect 28080 12232 28132 12238
rect 28078 12200 28080 12209
rect 28132 12200 28134 12209
rect 28078 12135 28134 12144
rect 27988 11620 28040 11626
rect 27988 11562 28040 11568
rect 28000 11150 28028 11562
rect 28080 11280 28132 11286
rect 28080 11222 28132 11228
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27988 11008 28040 11014
rect 27986 10976 27988 10985
rect 28040 10976 28042 10985
rect 27986 10911 28042 10920
rect 28092 10674 28120 11222
rect 28184 10674 28212 12310
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10810 28304 11018
rect 28264 10804 28316 10810
rect 28264 10746 28316 10752
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 27908 9710 28120 9738
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27724 9042 27752 9386
rect 27802 9344 27858 9353
rect 27802 9279 27858 9288
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27448 8214 27660 8242
rect 27632 7954 27660 8214
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27712 7472 27764 7478
rect 27712 7414 27764 7420
rect 27264 7364 27568 7392
rect 27344 7268 27396 7274
rect 27344 7210 27396 7216
rect 27068 6996 27120 7002
rect 27068 6938 27120 6944
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27080 6390 27108 6938
rect 27252 6928 27304 6934
rect 27356 6916 27384 7210
rect 27304 6888 27384 6916
rect 27252 6870 27304 6876
rect 27264 6798 27292 6870
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27068 6384 27120 6390
rect 27068 6326 27120 6332
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 26160 4078 26188 5578
rect 26252 4146 26280 5646
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26436 4010 26464 4490
rect 26620 4128 26648 5782
rect 27448 5574 27476 6190
rect 27436 5568 27488 5574
rect 27250 5536 27306 5545
rect 27436 5510 27488 5516
rect 27250 5471 27306 5480
rect 27264 5370 27292 5471
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 26792 5092 26844 5098
rect 26792 5034 26844 5040
rect 26804 4554 26832 5034
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 27344 4548 27396 4554
rect 27344 4490 27396 4496
rect 26528 4100 26648 4128
rect 26700 4140 26752 4146
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 25964 3528 26016 3534
rect 26160 3516 26188 3878
rect 25964 3470 26016 3476
rect 26068 3488 26188 3516
rect 25976 2689 26004 3470
rect 26068 2990 26096 3488
rect 26528 3466 26556 4100
rect 26700 4082 26752 4088
rect 26608 4004 26660 4010
rect 26608 3946 26660 3952
rect 26620 3602 26648 3946
rect 26608 3596 26660 3602
rect 26608 3538 26660 3544
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 26160 3058 26188 3130
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 25962 2680 26018 2689
rect 25962 2615 26018 2624
rect 26160 2378 26188 2994
rect 26436 2774 26464 3334
rect 26712 3233 26740 4082
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26988 3466 27016 3878
rect 27356 3738 27384 4490
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27448 3670 27476 4150
rect 27540 4078 27568 7364
rect 27724 6798 27752 7414
rect 27816 7002 27844 9279
rect 27894 9208 27950 9217
rect 27894 9143 27896 9152
rect 27948 9143 27950 9152
rect 27896 9114 27948 9120
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27816 6633 27844 6938
rect 27802 6624 27858 6633
rect 27802 6559 27858 6568
rect 27618 6488 27674 6497
rect 27618 6423 27674 6432
rect 27712 6452 27764 6458
rect 27632 5166 27660 6423
rect 27712 6394 27764 6400
rect 27724 6254 27752 6394
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27710 5808 27766 5817
rect 27710 5743 27766 5752
rect 27724 5370 27752 5743
rect 27816 5710 27844 6559
rect 27908 6458 27936 7142
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27804 5704 27856 5710
rect 27804 5646 27856 5652
rect 28000 5386 28028 9522
rect 28092 7206 28120 9710
rect 28368 9654 28396 12038
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28460 9518 28488 12922
rect 28644 11762 28672 32166
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 30116 30734 30144 31758
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 29276 19780 29328 19786
rect 29276 19722 29328 19728
rect 28816 13864 28868 13870
rect 28816 13806 28868 13812
rect 28828 12986 28856 13806
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28540 11008 28592 11014
rect 28540 10950 28592 10956
rect 28630 10976 28686 10985
rect 28552 10130 28580 10950
rect 28630 10911 28686 10920
rect 28644 10810 28672 10911
rect 28632 10804 28684 10810
rect 28632 10746 28684 10752
rect 28540 10124 28592 10130
rect 28540 10066 28592 10072
rect 28448 9512 28500 9518
rect 28170 9480 28226 9489
rect 28448 9454 28500 9460
rect 28170 9415 28226 9424
rect 28184 9042 28212 9415
rect 28814 9072 28870 9081
rect 28172 9036 28224 9042
rect 28814 9007 28870 9016
rect 28172 8978 28224 8984
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 28080 7200 28132 7206
rect 28078 7168 28080 7177
rect 28132 7168 28134 7177
rect 28078 7103 28134 7112
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28092 5846 28120 6734
rect 28080 5840 28132 5846
rect 28080 5782 28132 5788
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 27712 5364 27764 5370
rect 27712 5306 27764 5312
rect 27908 5358 28028 5386
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27908 5030 27936 5358
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27724 4554 27752 4694
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27620 4480 27672 4486
rect 27618 4448 27620 4457
rect 27672 4448 27674 4457
rect 27618 4383 27674 4392
rect 27908 4321 27936 4558
rect 27894 4312 27950 4321
rect 27894 4247 27950 4256
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27804 4072 27856 4078
rect 27804 4014 27856 4020
rect 27436 3664 27488 3670
rect 27436 3606 27488 3612
rect 27540 3534 27568 4014
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 26698 3224 26754 3233
rect 26698 3159 26754 3168
rect 27724 3058 27752 3402
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 26620 2854 26648 2994
rect 27816 2990 27844 4014
rect 28000 3534 28028 5170
rect 28092 3942 28120 5646
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 28184 3618 28212 7346
rect 28276 5914 28304 8502
rect 28724 7880 28776 7886
rect 28538 7848 28594 7857
rect 28724 7822 28776 7828
rect 28538 7783 28540 7792
rect 28592 7783 28594 7792
rect 28540 7754 28592 7760
rect 28356 7744 28408 7750
rect 28448 7744 28500 7750
rect 28356 7686 28408 7692
rect 28446 7712 28448 7721
rect 28500 7712 28502 7721
rect 28368 7546 28396 7686
rect 28446 7647 28502 7656
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28448 6724 28500 6730
rect 28448 6666 28500 6672
rect 28264 5908 28316 5914
rect 28264 5850 28316 5856
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28092 3590 28212 3618
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 28092 2854 28120 3590
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 26516 2848 26568 2854
rect 26608 2848 26660 2854
rect 26516 2790 26568 2796
rect 26606 2816 26608 2825
rect 28080 2848 28132 2854
rect 26660 2816 26662 2825
rect 26344 2746 26464 2774
rect 26344 2446 26372 2746
rect 26528 2514 26556 2790
rect 28080 2790 28132 2796
rect 26606 2751 26662 2760
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 25780 1964 25832 1970
rect 25780 1906 25832 1912
rect 26436 800 26464 2246
rect 27172 2106 27200 2382
rect 28184 2106 28212 3470
rect 28276 2514 28304 4694
rect 28368 3534 28396 6666
rect 28460 5370 28488 6666
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 27160 2100 27212 2106
rect 27160 2042 27212 2048
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28368 800 28396 2382
rect 28460 2310 28488 4966
rect 28552 4078 28580 7142
rect 28736 7002 28764 7822
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 28828 6730 28856 9007
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 28920 7546 28948 8910
rect 29012 8129 29040 12174
rect 29288 12102 29316 19722
rect 30116 18154 30144 30670
rect 30668 28218 30696 37130
rect 30760 29306 30788 37198
rect 32232 37126 32260 39200
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37466 35480 39200
rect 36726 38856 36782 38865
rect 36726 38791 36782 38800
rect 36740 37466 36768 38791
rect 35440 37460 35492 37466
rect 35440 37402 35492 37408
rect 36728 37460 36780 37466
rect 36728 37402 36780 37408
rect 35452 37262 35480 37402
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 36912 37256 36964 37262
rect 36912 37198 36964 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30656 28212 30708 28218
rect 30656 28154 30708 28160
rect 30104 18148 30156 18154
rect 30104 18090 30156 18096
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 29288 11801 29316 12038
rect 29274 11792 29330 11801
rect 29274 11727 29276 11736
rect 29328 11727 29330 11736
rect 29276 11698 29328 11704
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 29748 11354 29776 11494
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29840 11286 29868 15438
rect 30104 12640 30156 12646
rect 30104 12582 30156 12588
rect 30116 12374 30144 12582
rect 30944 12434 30972 29106
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 31220 27878 31248 28018
rect 31208 27872 31260 27878
rect 31208 27814 31260 27820
rect 31220 13462 31248 27814
rect 33612 26042 33640 37198
rect 35532 37188 35584 37194
rect 35532 37130 35584 37136
rect 35544 36718 35572 37130
rect 35532 36712 35584 36718
rect 35532 36654 35584 36660
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 34164 24410 34192 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 36924 26586 36952 37198
rect 37384 37126 37412 39200
rect 38198 37496 38254 37505
rect 38198 37431 38254 37440
rect 37464 37256 37516 37262
rect 37464 37198 37516 37204
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 37476 36718 37504 37198
rect 37464 36712 37516 36718
rect 37464 36654 37516 36660
rect 37924 36644 37976 36650
rect 37924 36586 37976 36592
rect 37740 36168 37792 36174
rect 37740 36110 37792 36116
rect 37372 26920 37424 26926
rect 37372 26862 37424 26868
rect 36912 26580 36964 26586
rect 36912 26522 36964 26528
rect 34244 25900 34296 25906
rect 34244 25842 34296 25848
rect 34256 25702 34284 25842
rect 34244 25696 34296 25702
rect 34244 25638 34296 25644
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 33416 24064 33468 24070
rect 33416 24006 33468 24012
rect 33428 20262 33456 24006
rect 33416 20256 33468 20262
rect 33416 20198 33468 20204
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 33060 18222 33088 18566
rect 33048 18216 33100 18222
rect 33048 18158 33100 18164
rect 32956 17128 33008 17134
rect 32956 17070 33008 17076
rect 32968 16250 32996 17070
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 31300 14544 31352 14550
rect 31300 14486 31352 14492
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 30852 12406 30972 12434
rect 30104 12368 30156 12374
rect 30104 12310 30156 12316
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30392 11626 30420 11834
rect 30380 11620 30432 11626
rect 30380 11562 30432 11568
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 29828 11280 29880 11286
rect 29828 11222 29880 11228
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 29656 11014 29684 11222
rect 29840 11150 29868 11222
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29748 9110 29776 9454
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 29840 9042 29868 9998
rect 29828 9036 29880 9042
rect 29828 8978 29880 8984
rect 29276 8968 29328 8974
rect 29276 8910 29328 8916
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 29104 8401 29132 8434
rect 29090 8392 29146 8401
rect 29090 8327 29146 8336
rect 29196 8265 29224 8502
rect 29182 8256 29238 8265
rect 29182 8191 29238 8200
rect 28998 8120 29054 8129
rect 29054 8064 29224 8072
rect 28998 8055 29224 8064
rect 29012 8044 29224 8055
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 28908 7336 28960 7342
rect 29012 7290 29040 7890
rect 29090 7440 29146 7449
rect 29196 7410 29224 8044
rect 29090 7375 29146 7384
rect 29184 7404 29236 7410
rect 28960 7284 29040 7290
rect 28908 7278 29040 7284
rect 28920 7262 29040 7278
rect 28816 6724 28868 6730
rect 28816 6666 28868 6672
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 28644 5953 28672 6394
rect 28736 6322 28764 6394
rect 28724 6316 28776 6322
rect 28724 6258 28776 6264
rect 28630 5944 28686 5953
rect 28630 5879 28686 5888
rect 28736 5352 28764 6258
rect 28814 6216 28870 6225
rect 28814 6151 28870 6160
rect 28644 5324 28764 5352
rect 28644 5234 28672 5324
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28644 4128 28672 5170
rect 28736 4865 28764 5170
rect 28828 5030 28856 6151
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28722 4856 28778 4865
rect 28722 4791 28778 4800
rect 28908 4616 28960 4622
rect 28908 4558 28960 4564
rect 28816 4140 28868 4146
rect 28644 4100 28816 4128
rect 28816 4082 28868 4088
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28828 3058 28856 4082
rect 28920 3534 28948 4558
rect 29012 4146 29040 7262
rect 29104 5386 29132 7375
rect 29184 7346 29236 7352
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29196 6798 29224 6938
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29184 6656 29236 6662
rect 29182 6624 29184 6633
rect 29236 6624 29238 6633
rect 29182 6559 29238 6568
rect 29288 6202 29316 8910
rect 29644 8900 29696 8906
rect 29644 8842 29696 8848
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 29366 8528 29422 8537
rect 29366 8463 29422 8472
rect 29380 8430 29408 8463
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 29368 6792 29420 6798
rect 29368 6734 29420 6740
rect 29380 6322 29408 6734
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29288 6174 29408 6202
rect 29104 5358 29316 5386
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29196 5030 29224 5170
rect 29184 5024 29236 5030
rect 29090 4992 29146 5001
rect 29184 4966 29236 4972
rect 29090 4927 29146 4936
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29104 2938 29132 4927
rect 29196 4049 29224 4966
rect 29288 4078 29316 5358
rect 29276 4072 29328 4078
rect 29182 4040 29238 4049
rect 29276 4014 29328 4020
rect 29182 3975 29238 3984
rect 29380 3398 29408 6174
rect 29472 4826 29500 8570
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 5914 29592 8230
rect 29656 8090 29684 8842
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29748 7818 29776 8230
rect 29736 7812 29788 7818
rect 29736 7754 29788 7760
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29564 4457 29592 4558
rect 29656 4486 29684 6054
rect 29736 5568 29788 5574
rect 29736 5510 29788 5516
rect 29748 5098 29776 5510
rect 29932 5370 29960 8842
rect 29920 5364 29972 5370
rect 29920 5306 29972 5312
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29736 5092 29788 5098
rect 29736 5034 29788 5040
rect 29734 4720 29790 4729
rect 29734 4655 29790 4664
rect 29644 4480 29696 4486
rect 29550 4448 29606 4457
rect 29644 4422 29696 4428
rect 29550 4383 29606 4392
rect 29368 3392 29420 3398
rect 29748 3369 29776 4655
rect 29840 4282 29868 5170
rect 30024 4865 30052 11086
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 10198 30144 10406
rect 30104 10192 30156 10198
rect 30104 10134 30156 10140
rect 30288 10056 30340 10062
rect 30340 10004 30420 10010
rect 30288 9998 30420 10004
rect 30300 9982 30420 9998
rect 30392 9586 30420 9982
rect 30484 9654 30512 11222
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 30562 10160 30618 10169
rect 30562 10095 30618 10104
rect 30472 9648 30524 9654
rect 30472 9590 30524 9596
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30392 9058 30420 9522
rect 30300 9030 30420 9058
rect 30484 9042 30512 9590
rect 30472 9036 30524 9042
rect 30300 8514 30328 9030
rect 30472 8978 30524 8984
rect 30378 8936 30434 8945
rect 30378 8871 30434 8880
rect 30392 8634 30420 8871
rect 30470 8664 30526 8673
rect 30380 8628 30432 8634
rect 30470 8599 30526 8608
rect 30380 8570 30432 8576
rect 30300 8486 30420 8514
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30116 5710 30144 6258
rect 30300 5914 30328 8298
rect 30288 5908 30340 5914
rect 30288 5850 30340 5856
rect 30392 5846 30420 8486
rect 30484 8090 30512 8599
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30576 7546 30604 10095
rect 30564 7540 30616 7546
rect 30564 7482 30616 7488
rect 30470 6760 30526 6769
rect 30470 6695 30526 6704
rect 30484 6662 30512 6695
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30564 6384 30616 6390
rect 30562 6352 30564 6361
rect 30616 6352 30618 6361
rect 30562 6287 30618 6296
rect 30562 6080 30618 6089
rect 30562 6015 30618 6024
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30010 4856 30066 4865
rect 30010 4791 30066 4800
rect 30012 4752 30064 4758
rect 30012 4694 30064 4700
rect 30024 4486 30052 4694
rect 30012 4480 30064 4486
rect 30012 4422 30064 4428
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 30116 4078 30144 5646
rect 30380 5636 30432 5642
rect 30380 5578 30432 5584
rect 30392 5302 30420 5578
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 30484 5234 30512 5646
rect 30576 5370 30604 6015
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30208 4690 30236 4762
rect 30196 4684 30248 4690
rect 30196 4626 30248 4632
rect 30300 4146 30328 4966
rect 30484 4622 30512 5170
rect 30668 4622 30696 11086
rect 30852 8566 30880 12406
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 30944 11558 30972 11766
rect 30932 11552 30984 11558
rect 30932 11494 30984 11500
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 30932 9172 30984 9178
rect 30932 9114 30984 9120
rect 30944 8838 30972 9114
rect 30932 8832 30984 8838
rect 30930 8800 30932 8809
rect 30984 8800 30986 8809
rect 30930 8735 30986 8744
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30760 7886 30788 8434
rect 31036 8294 31064 11154
rect 31312 11014 31340 14486
rect 34256 14278 34284 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 37292 21894 37320 22578
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35440 15632 35492 15638
rect 35440 15574 35492 15580
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 34256 13870 34284 14214
rect 34244 13864 34296 13870
rect 34244 13806 34296 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34152 12776 34204 12782
rect 34152 12718 34204 12724
rect 34164 11898 34192 12718
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 31482 11656 31538 11665
rect 31482 11591 31538 11600
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31300 11008 31352 11014
rect 31300 10950 31352 10956
rect 31404 10674 31432 11018
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31404 10470 31432 10610
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 31024 8288 31076 8294
rect 31024 8230 31076 8236
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 31300 7880 31352 7886
rect 31300 7822 31352 7828
rect 30760 6458 30788 7822
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 31022 7304 31078 7313
rect 31022 7239 31024 7248
rect 31076 7239 31078 7248
rect 31024 7210 31076 7216
rect 31022 7032 31078 7041
rect 31022 6967 31078 6976
rect 30748 6452 30800 6458
rect 30748 6394 30800 6400
rect 31036 5914 31064 6967
rect 31128 6798 31156 7346
rect 31312 6798 31340 7822
rect 31404 7818 31432 10406
rect 31392 7812 31444 7818
rect 31392 7754 31444 7760
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31116 6656 31168 6662
rect 31208 6656 31260 6662
rect 31116 6598 31168 6604
rect 31206 6624 31208 6633
rect 31260 6624 31262 6633
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 31128 5778 31156 6598
rect 31206 6559 31262 6568
rect 31208 6316 31260 6322
rect 31312 6304 31340 6734
rect 31260 6276 31340 6304
rect 31208 6258 31260 6264
rect 31116 5772 31168 5778
rect 31116 5714 31168 5720
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31220 4826 31248 5170
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31312 4622 31340 6276
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 31404 5234 31432 6258
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31496 4758 31524 11591
rect 32402 10024 32458 10033
rect 32402 9959 32458 9968
rect 31576 8288 31628 8294
rect 31576 8230 31628 8236
rect 31588 7274 31616 8230
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 31772 7993 31800 8026
rect 31758 7984 31814 7993
rect 31758 7919 31814 7928
rect 31576 7268 31628 7274
rect 31576 7210 31628 7216
rect 31588 6866 31616 7210
rect 32220 7200 32272 7206
rect 32220 7142 32272 7148
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 31852 6656 31904 6662
rect 31852 6598 31904 6604
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 31772 5914 31800 6190
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31758 5672 31814 5681
rect 31758 5607 31814 5616
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31680 4826 31708 4966
rect 31772 4826 31800 5607
rect 31668 4820 31720 4826
rect 31668 4762 31720 4768
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31484 4752 31536 4758
rect 31404 4700 31484 4706
rect 31404 4694 31536 4700
rect 31404 4678 31524 4694
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 30668 4457 30696 4558
rect 30654 4448 30710 4457
rect 30654 4383 30710 4392
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 30208 3942 30236 4082
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30300 3534 30328 4082
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30760 3777 30788 3878
rect 30746 3768 30802 3777
rect 30746 3703 30802 3712
rect 30932 3664 30984 3670
rect 30932 3606 30984 3612
rect 31206 3632 31262 3641
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30472 3392 30524 3398
rect 29368 3334 29420 3340
rect 29734 3360 29790 3369
rect 30472 3334 30524 3340
rect 29734 3295 29790 3304
rect 29748 3058 29776 3295
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 29012 2910 29132 2938
rect 29012 2854 29040 2910
rect 28816 2848 28868 2854
rect 29000 2848 29052 2854
rect 28868 2808 28948 2836
rect 28816 2790 28868 2796
rect 28920 2446 28948 2808
rect 29000 2790 29052 2796
rect 30484 2582 30512 3334
rect 30944 3058 30972 3606
rect 31206 3567 31262 3576
rect 31220 3534 31248 3567
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31036 3058 31064 3470
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 30564 2984 30616 2990
rect 30564 2926 30616 2932
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30576 2514 30604 2926
rect 31220 2854 31248 3470
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 31404 2514 31432 4678
rect 31484 4548 31536 4554
rect 31484 4490 31536 4496
rect 31496 4146 31524 4490
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31496 2650 31524 4082
rect 31576 4004 31628 4010
rect 31576 3946 31628 3952
rect 31588 3233 31616 3946
rect 31680 3584 31708 4762
rect 31864 4622 31892 6598
rect 31852 4616 31904 4622
rect 31852 4558 31904 4564
rect 31864 3670 31892 4558
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32140 3942 32168 4082
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 31680 3556 31800 3584
rect 31772 3516 31800 3556
rect 31852 3528 31904 3534
rect 31772 3488 31852 3516
rect 31852 3470 31904 3476
rect 31668 3460 31720 3466
rect 31668 3402 31720 3408
rect 31574 3224 31630 3233
rect 31574 3159 31630 3168
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 31392 2508 31444 2514
rect 31392 2450 31444 2456
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 28448 2304 28500 2310
rect 28448 2246 28500 2252
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 30564 2304 30616 2310
rect 30564 2246 30616 2252
rect 31208 2304 31260 2310
rect 31208 2246 31260 2252
rect 29656 800 29684 2246
rect 30576 2038 30604 2246
rect 30564 2032 30616 2038
rect 30564 1974 30616 1980
rect 31220 1970 31248 2246
rect 31208 1964 31260 1970
rect 31208 1906 31260 1912
rect 31588 800 31616 2382
rect 31680 2281 31708 3402
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 31666 2272 31722 2281
rect 31666 2207 31722 2216
rect 31772 1873 31800 3334
rect 31864 3126 31892 3470
rect 31852 3120 31904 3126
rect 31852 3062 31904 3068
rect 32232 2514 32260 7142
rect 32416 6458 32444 9959
rect 32588 7268 32640 7274
rect 32588 7210 32640 7216
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32404 6452 32456 6458
rect 32404 6394 32456 6400
rect 32508 6322 32536 6734
rect 32600 6662 32628 7210
rect 32588 6656 32640 6662
rect 32864 6656 32916 6662
rect 32588 6598 32640 6604
rect 32862 6624 32864 6633
rect 32916 6624 32918 6633
rect 32496 6316 32548 6322
rect 32496 6258 32548 6264
rect 32508 5710 32536 6258
rect 32600 6186 32628 6598
rect 32862 6559 32918 6568
rect 32588 6180 32640 6186
rect 32588 6122 32640 6128
rect 32496 5704 32548 5710
rect 32496 5646 32548 5652
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32402 5128 32458 5137
rect 32324 2854 32352 5102
rect 32402 5063 32404 5072
rect 32456 5063 32458 5072
rect 32404 5034 32456 5040
rect 32402 4584 32458 4593
rect 32402 4519 32404 4528
rect 32456 4519 32458 4528
rect 32404 4490 32456 4496
rect 32600 4146 32628 5170
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 32404 3936 32456 3942
rect 32402 3904 32404 3913
rect 32680 3936 32732 3942
rect 32456 3904 32458 3913
rect 32680 3878 32732 3884
rect 32402 3839 32458 3848
rect 32588 3732 32640 3738
rect 32588 3674 32640 3680
rect 32402 2952 32458 2961
rect 32402 2887 32404 2896
rect 32456 2887 32458 2896
rect 32496 2916 32548 2922
rect 32404 2858 32456 2864
rect 32496 2858 32548 2864
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 32324 2582 32352 2790
rect 32312 2576 32364 2582
rect 32508 2553 32536 2858
rect 32312 2518 32364 2524
rect 32494 2544 32550 2553
rect 32220 2508 32272 2514
rect 32494 2479 32550 2488
rect 32220 2450 32272 2456
rect 31758 1864 31814 1873
rect 32232 1834 32260 2450
rect 32600 2446 32628 3674
rect 32588 2440 32640 2446
rect 32692 2417 32720 3878
rect 32876 3534 32904 5646
rect 33048 5568 33100 5574
rect 33048 5510 33100 5516
rect 33060 5273 33088 5510
rect 33244 5409 33272 11834
rect 33508 11552 33560 11558
rect 33508 11494 33560 11500
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6118 33364 6598
rect 33324 6112 33376 6118
rect 33324 6054 33376 6060
rect 33336 5710 33364 6054
rect 33324 5704 33376 5710
rect 33324 5646 33376 5652
rect 33230 5400 33286 5409
rect 33230 5335 33286 5344
rect 33046 5264 33102 5273
rect 33046 5199 33102 5208
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 33244 4690 33272 5170
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 33244 3534 33272 4626
rect 33336 4214 33364 5646
rect 33324 4208 33376 4214
rect 33324 4150 33376 4156
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 33232 3392 33284 3398
rect 33336 3369 33364 3538
rect 33232 3334 33284 3340
rect 33322 3360 33378 3369
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 32588 2382 32640 2388
rect 32678 2408 32734 2417
rect 32678 2343 32734 2352
rect 33060 1902 33088 2790
rect 33244 2009 33272 3334
rect 33322 3295 33378 3304
rect 33520 2582 33548 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 33692 6180 33744 6186
rect 33692 6122 33744 6128
rect 33600 5568 33652 5574
rect 33600 5510 33652 5516
rect 33612 5030 33640 5510
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 4486 33640 4966
rect 33704 4690 33732 6122
rect 33692 4684 33744 4690
rect 33692 4626 33744 4632
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 33692 3936 33744 3942
rect 33692 3878 33744 3884
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33704 3505 33732 3878
rect 33796 3738 33824 3878
rect 33784 3732 33836 3738
rect 33784 3674 33836 3680
rect 33876 3664 33928 3670
rect 33876 3606 33928 3612
rect 33690 3496 33746 3505
rect 33690 3431 33746 3440
rect 33692 3120 33744 3126
rect 33690 3088 33692 3097
rect 33744 3088 33746 3097
rect 33888 3058 33916 3606
rect 33690 3023 33746 3032
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 33508 2576 33560 2582
rect 33508 2518 33560 2524
rect 33888 2514 33916 2994
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 33980 2446 34008 6598
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35452 5914 35480 15574
rect 37292 14074 37320 21830
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 35808 13864 35860 13870
rect 35808 13806 35860 13812
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 35256 5704 35308 5710
rect 35256 5646 35308 5652
rect 34150 5400 34206 5409
rect 35268 5370 35296 5646
rect 34150 5335 34152 5344
rect 34204 5335 34206 5344
rect 35256 5364 35308 5370
rect 34152 5306 34204 5312
rect 35256 5306 35308 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 34348 3738 34376 4626
rect 34796 4548 34848 4554
rect 34796 4490 34848 4496
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 34348 2650 34376 3674
rect 34808 3670 34836 4490
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3664 34848 3670
rect 34796 3606 34848 3612
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34440 3058 34468 3470
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34532 2689 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34518 2680 34574 2689
rect 34934 2683 35242 2692
rect 34336 2644 34388 2650
rect 34518 2615 34574 2624
rect 34336 2586 34388 2592
rect 35452 2446 35480 5850
rect 35716 4480 35768 4486
rect 35716 4422 35768 4428
rect 35728 4146 35756 4422
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35728 3738 35756 4082
rect 35716 3732 35768 3738
rect 35716 3674 35768 3680
rect 35820 2650 35848 13806
rect 35900 11688 35952 11694
rect 35900 11630 35952 11636
rect 35912 7410 35940 11630
rect 37384 9178 37412 26862
rect 37464 24948 37516 24954
rect 37464 24890 37516 24896
rect 37476 12374 37504 24890
rect 37464 12368 37516 12374
rect 37464 12310 37516 12316
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 36452 6112 36504 6118
rect 36452 6054 36504 6060
rect 36464 5574 36492 6054
rect 37476 5846 37504 12310
rect 37752 8090 37780 36110
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37844 16114 37872 25230
rect 37936 24818 37964 36586
rect 38212 36378 38240 37431
rect 38672 36854 38700 39200
rect 38660 36848 38712 36854
rect 38660 36790 38712 36796
rect 38200 36372 38252 36378
rect 38200 36314 38252 36320
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38200 33516 38252 33522
rect 38200 33458 38252 33464
rect 38212 33425 38240 33458
rect 38198 33416 38254 33425
rect 38198 33351 38254 33360
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 38016 30864 38068 30870
rect 38016 30806 38068 30812
rect 38028 30258 38056 30806
rect 38016 30252 38068 30258
rect 38016 30194 38068 30200
rect 38016 26376 38068 26382
rect 38016 26318 38068 26324
rect 38028 25702 38056 26318
rect 38120 26234 38148 32370
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38292 27328 38344 27334
rect 38292 27270 38344 27276
rect 38304 26926 38332 27270
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 38304 26625 38332 26862
rect 38290 26616 38346 26625
rect 38290 26551 38346 26560
rect 38120 26206 38240 26234
rect 38016 25696 38068 25702
rect 38016 25638 38068 25644
rect 38028 24954 38056 25638
rect 38212 25498 38240 26206
rect 38200 25492 38252 25498
rect 38200 25434 38252 25440
rect 38016 24948 38068 24954
rect 38016 24890 38068 24896
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 38108 24812 38160 24818
rect 38108 24754 38160 24760
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 38028 22778 38056 23666
rect 38016 22772 38068 22778
rect 38016 22714 38068 22720
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 38028 15706 38056 21490
rect 38120 21146 38148 24754
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38200 23520 38252 23526
rect 38200 23462 38252 23468
rect 38212 23225 38240 23462
rect 38198 23216 38254 23225
rect 38198 23151 38254 23160
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38108 21140 38160 21146
rect 38198 21111 38254 21120
rect 38108 21082 38160 21088
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38120 19718 38148 20878
rect 38292 19848 38344 19854
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 38290 19751 38346 19760
rect 38108 19712 38160 19718
rect 38108 19654 38160 19660
rect 38120 18766 38148 19654
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 38292 16040 38344 16046
rect 38292 15982 38344 15988
rect 38304 15745 38332 15982
rect 38290 15736 38346 15745
rect 38016 15700 38068 15706
rect 38290 15671 38292 15680
rect 38016 15642 38068 15648
rect 38344 15671 38346 15680
rect 38292 15642 38344 15648
rect 38016 14408 38068 14414
rect 38292 14408 38344 14414
rect 38016 14350 38068 14356
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38028 12918 38056 14350
rect 38290 14311 38346 14320
rect 38304 14074 38332 14311
rect 38292 14068 38344 14074
rect 38292 14010 38344 14016
rect 38016 12912 38068 12918
rect 38016 12854 38068 12860
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37464 5840 37516 5846
rect 37464 5782 37516 5788
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 36096 2446 36124 5510
rect 36464 5030 36492 5510
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36464 4554 36492 4966
rect 36452 4548 36504 4554
rect 36452 4490 36504 4496
rect 36464 4282 36492 4490
rect 36452 4276 36504 4282
rect 36452 4218 36504 4224
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36280 3126 36308 4014
rect 36464 3534 36492 4218
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 36268 3120 36320 3126
rect 36268 3062 36320 3068
rect 36464 3058 36492 3470
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 36924 2446 36952 2994
rect 37660 2514 37688 6598
rect 37936 4146 37964 10950
rect 38028 10674 38056 12854
rect 38292 12776 38344 12782
rect 38292 12718 38344 12724
rect 38304 12374 38332 12718
rect 38292 12368 38344 12374
rect 38290 12336 38292 12345
rect 38344 12336 38346 12345
rect 38290 12271 38346 12280
rect 38304 12245 38332 12271
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38304 11150 38332 11494
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 38028 8974 38056 10406
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 38304 6934 38332 7278
rect 38292 6928 38344 6934
rect 38290 6896 38292 6905
rect 38344 6896 38346 6905
rect 38290 6831 38346 6840
rect 38292 6112 38344 6118
rect 38292 6054 38344 6060
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 38212 5545 38240 5578
rect 38198 5536 38254 5545
rect 38198 5471 38254 5480
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 38028 4622 38056 4966
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 33230 2000 33286 2009
rect 33230 1935 33286 1944
rect 33048 1896 33100 1902
rect 33048 1838 33100 1844
rect 31758 1799 31814 1808
rect 32220 1828 32272 1834
rect 32220 1770 32272 1776
rect 33520 800 33548 2382
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 34808 800 34836 2246
rect 36740 800 36768 2382
rect 37660 2145 37688 2450
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37646 2136 37702 2145
rect 37646 2071 37702 2080
rect 37752 1970 37780 2382
rect 37740 1964 37792 1970
rect 37740 1906 37792 1912
rect 38028 800 38056 4558
rect 38108 4480 38160 4486
rect 38108 4422 38160 4428
rect 38120 3194 38148 4422
rect 38304 4214 38332 6054
rect 38292 4208 38344 4214
rect 38292 4150 38344 4156
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 38108 3188 38160 3194
rect 38108 3130 38160 3136
rect 14476 734 14780 762
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36726 200 36782 800
rect 38014 200 38070 800
rect 38304 105 38332 4150
rect 38290 96 38346 105
rect 38290 31 38346 40
<< via2 >>
rect 2870 38800 2926 38856
rect 1674 36780 1730 36816
rect 1674 36760 1676 36780
rect 1676 36760 1728 36780
rect 1728 36760 1730 36780
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1674 33360 1730 33416
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1582 31356 1584 31376
rect 1584 31356 1636 31376
rect 1636 31356 1638 31376
rect 1582 31320 1638 31356
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1582 29960 1638 30016
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 26560 1730 26616
rect 1674 24556 1676 24576
rect 1676 24556 1728 24576
rect 1728 24556 1730 24576
rect 1674 24520 1730 24556
rect 1674 22500 1730 22536
rect 1674 22480 1676 22500
rect 1676 22480 1728 22500
rect 1728 22480 1730 22500
rect 1582 21140 1638 21176
rect 1582 21120 1584 21140
rect 1584 21120 1636 21140
rect 1636 21120 1638 21140
rect 1582 19080 1638 19136
rect 1674 17720 1730 17776
rect 1674 15680 1730 15736
rect 1674 13640 1730 13696
rect 1674 12280 1730 12336
rect 1674 10240 1730 10296
rect 1674 8900 1730 8936
rect 1674 8880 1676 8900
rect 1676 8880 1728 8900
rect 1728 8880 1730 8900
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 6840 1638 6896
rect 1582 4820 1638 4856
rect 1582 4800 1584 4820
rect 1584 4800 1636 4820
rect 1636 4800 1638 4820
rect 1674 3476 1676 3496
rect 1676 3476 1728 3496
rect 1728 3476 1730 3496
rect 1674 3440 1730 3476
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8114 3596 8170 3632
rect 8114 3576 8116 3596
rect 8116 3576 8168 3596
rect 8168 3576 8170 3596
rect 10506 31764 10508 31784
rect 10508 31764 10560 31784
rect 10560 31764 10562 31784
rect 10506 31728 10562 31764
rect 9770 11736 9826 11792
rect 9862 9596 9864 9616
rect 9864 9596 9916 9616
rect 9916 9596 9918 9616
rect 9862 9560 9918 9596
rect 9310 9444 9366 9480
rect 9310 9424 9312 9444
rect 9312 9424 9364 9444
rect 9364 9424 9366 9444
rect 9494 5636 9550 5672
rect 9494 5616 9496 5636
rect 9496 5616 9548 5636
rect 9548 5616 9550 5636
rect 9770 5344 9826 5400
rect 10414 4800 10470 4856
rect 1674 1400 1730 1456
rect 17130 26832 17186 26888
rect 13634 13912 13690 13968
rect 11058 11228 11060 11248
rect 11060 11228 11112 11248
rect 11112 11228 11114 11248
rect 11058 11192 11114 11228
rect 10966 10532 11022 10568
rect 10966 10512 10968 10532
rect 10968 10512 11020 10532
rect 11020 10512 11022 10532
rect 10874 6860 10930 6896
rect 10874 6840 10876 6860
rect 10876 6840 10928 6860
rect 10928 6840 10930 6860
rect 13266 13640 13322 13696
rect 12898 13096 12954 13152
rect 13174 12688 13230 12744
rect 12254 7404 12310 7440
rect 12254 7384 12256 7404
rect 12256 7384 12308 7404
rect 12308 7384 12310 7404
rect 12438 6740 12440 6760
rect 12440 6740 12492 6760
rect 12492 6740 12494 6760
rect 12438 6704 12494 6740
rect 12438 4120 12494 4176
rect 12714 4004 12770 4040
rect 12714 3984 12716 4004
rect 12716 3984 12768 4004
rect 12768 3984 12770 4004
rect 12070 3168 12126 3224
rect 13358 3848 13414 3904
rect 12622 3168 12678 3224
rect 13726 13640 13782 13696
rect 13726 13504 13782 13560
rect 13818 11328 13874 11384
rect 13634 5752 13690 5808
rect 14278 11192 14334 11248
rect 14186 10784 14242 10840
rect 14370 8880 14426 8936
rect 14554 9016 14610 9072
rect 14830 10648 14886 10704
rect 14738 9424 14794 9480
rect 14738 7248 14794 7304
rect 14738 6840 14794 6896
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 15198 13132 15200 13152
rect 15200 13132 15252 13152
rect 15252 13132 15254 13152
rect 15198 13096 15254 13132
rect 16210 14592 16266 14648
rect 15014 10784 15070 10840
rect 15014 10376 15070 10432
rect 15106 9988 15162 10024
rect 15106 9968 15108 9988
rect 15108 9968 15160 9988
rect 15160 9968 15162 9988
rect 15106 9560 15162 9616
rect 15382 9424 15438 9480
rect 15106 9016 15162 9072
rect 15106 8744 15162 8800
rect 14462 6724 14518 6760
rect 14462 6704 14464 6724
rect 14464 6704 14516 6724
rect 14516 6704 14518 6724
rect 14278 5092 14334 5128
rect 14278 5072 14280 5092
rect 14280 5072 14332 5092
rect 14332 5072 14334 5092
rect 14278 4684 14334 4720
rect 14278 4664 14280 4684
rect 14280 4664 14332 4684
rect 14332 4664 14334 4684
rect 15014 5616 15070 5672
rect 14738 5344 14794 5400
rect 15014 5244 15016 5264
rect 15016 5244 15068 5264
rect 15068 5244 15070 5264
rect 15014 5208 15070 5244
rect 15566 10512 15622 10568
rect 15842 11772 15844 11792
rect 15844 11772 15896 11792
rect 15896 11772 15898 11792
rect 15842 11736 15898 11772
rect 16118 11736 16174 11792
rect 15658 9424 15714 9480
rect 15382 5108 15384 5128
rect 15384 5108 15436 5128
rect 15436 5108 15438 5128
rect 15382 5072 15438 5108
rect 14830 4664 14886 4720
rect 16578 13504 16634 13560
rect 16486 12164 16542 12200
rect 16486 12144 16488 12164
rect 16488 12144 16540 12164
rect 16540 12144 16542 12164
rect 15934 8880 15990 8936
rect 16486 8900 16542 8936
rect 16486 8880 16488 8900
rect 16488 8880 16540 8900
rect 16540 8880 16542 8900
rect 16210 5616 16266 5672
rect 16762 10376 16818 10432
rect 17222 13912 17278 13968
rect 17038 12724 17040 12744
rect 17040 12724 17092 12744
rect 17092 12724 17094 12744
rect 17038 12688 17094 12724
rect 16210 3460 16266 3496
rect 16210 3440 16212 3460
rect 16212 3440 16264 3460
rect 16264 3440 16266 3460
rect 16118 3068 16120 3088
rect 16120 3068 16172 3088
rect 16172 3068 16174 3088
rect 16118 3032 16174 3068
rect 15290 2372 15346 2408
rect 15290 2352 15292 2372
rect 15292 2352 15344 2372
rect 15344 2352 15346 2372
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 17866 11636 17868 11656
rect 17868 11636 17920 11656
rect 17920 11636 17922 11656
rect 17866 11600 17922 11636
rect 18234 11328 18290 11384
rect 18326 10784 18382 10840
rect 18142 8744 18198 8800
rect 17590 6296 17646 6352
rect 17314 4800 17370 4856
rect 17866 5072 17922 5128
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19798 13640 19854 13696
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20074 12144 20130 12200
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19430 10512 19486 10568
rect 19338 10240 19394 10296
rect 19246 10104 19302 10160
rect 19338 9832 19394 9888
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19338 9696 19394 9752
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 17866 4020 17868 4040
rect 17868 4020 17920 4040
rect 17920 4020 17922 4040
rect 17866 3984 17922 4020
rect 17866 1808 17922 1864
rect 20810 12008 20866 12064
rect 20626 9696 20682 9752
rect 20166 6568 20222 6624
rect 18970 2896 19026 2952
rect 19338 4936 19394 4992
rect 19154 3848 19210 3904
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19982 4664 20038 4720
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20258 5636 20314 5672
rect 20258 5616 20260 5636
rect 20260 5616 20312 5636
rect 20312 5616 20314 5636
rect 20994 10668 21050 10704
rect 20994 10648 20996 10668
rect 20996 10648 21048 10668
rect 21048 10648 21050 10668
rect 21546 14592 21602 14648
rect 21270 10512 21326 10568
rect 20718 8608 20774 8664
rect 20534 7520 20590 7576
rect 20902 7112 20958 7168
rect 20718 6976 20774 7032
rect 20626 6840 20682 6896
rect 20718 5888 20774 5944
rect 20442 4120 20498 4176
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 19154 1944 19210 2000
rect 20626 2760 20682 2816
rect 24950 16224 25006 16280
rect 22466 11636 22468 11656
rect 22468 11636 22520 11656
rect 22520 11636 22522 11656
rect 22466 11600 22522 11636
rect 21454 7656 21510 7712
rect 21822 6160 21878 6216
rect 22374 7540 22430 7576
rect 22374 7520 22376 7540
rect 22376 7520 22428 7540
rect 22428 7520 22430 7540
rect 22282 6840 22338 6896
rect 22282 6432 22338 6488
rect 22190 6024 22246 6080
rect 23754 12144 23810 12200
rect 24030 12008 24086 12064
rect 23754 8744 23810 8800
rect 22650 4528 22706 4584
rect 22006 4004 22062 4040
rect 22006 3984 22008 4004
rect 22008 3984 22060 4004
rect 22060 3984 22062 4004
rect 21914 3712 21970 3768
rect 22374 4120 22430 4176
rect 22098 3168 22154 3224
rect 23294 6860 23350 6896
rect 23294 6840 23296 6860
rect 23296 6840 23348 6860
rect 23348 6840 23350 6860
rect 23478 6180 23534 6216
rect 23478 6160 23480 6180
rect 23480 6160 23532 6180
rect 23532 6160 23534 6180
rect 23662 3848 23718 3904
rect 24766 9152 24822 9208
rect 24766 8064 24822 8120
rect 25318 11464 25374 11520
rect 26330 12144 26386 12200
rect 24306 4800 24362 4856
rect 24122 4392 24178 4448
rect 25870 10240 25926 10296
rect 25410 7928 25466 7984
rect 24950 6160 25006 6216
rect 24030 3168 24086 3224
rect 23662 2216 23718 2272
rect 24674 4256 24730 4312
rect 24398 2488 24454 2544
rect 25502 6704 25558 6760
rect 26146 9016 26202 9072
rect 27250 16224 27306 16280
rect 26606 9460 26608 9480
rect 26608 9460 26660 9480
rect 26660 9460 26662 9480
rect 26606 9424 26662 9460
rect 26514 9288 26570 9344
rect 26606 8200 26662 8256
rect 25778 5752 25834 5808
rect 25870 5344 25926 5400
rect 25410 3168 25466 3224
rect 27250 11464 27306 11520
rect 26790 8200 26846 8256
rect 26790 6840 26846 6896
rect 26698 6160 26754 6216
rect 27526 12008 27582 12064
rect 27066 7812 27122 7848
rect 27066 7792 27068 7812
rect 27068 7792 27120 7812
rect 27120 7792 27122 7812
rect 27526 8492 27582 8528
rect 27526 8472 27528 8492
rect 27528 8472 27580 8492
rect 27580 8472 27582 8492
rect 28078 12180 28080 12200
rect 28080 12180 28132 12200
rect 28132 12180 28134 12200
rect 28078 12144 28134 12180
rect 27986 10956 27988 10976
rect 27988 10956 28040 10976
rect 28040 10956 28042 10976
rect 27986 10920 28042 10956
rect 27802 9288 27858 9344
rect 27250 5480 27306 5536
rect 25962 2624 26018 2680
rect 27894 9172 27950 9208
rect 27894 9152 27896 9172
rect 27896 9152 27948 9172
rect 27948 9152 27950 9172
rect 27802 6568 27858 6624
rect 27618 6432 27674 6488
rect 27710 5752 27766 5808
rect 28630 10920 28686 10976
rect 28170 9424 28226 9480
rect 28814 9016 28870 9072
rect 28078 7148 28080 7168
rect 28080 7148 28132 7168
rect 28132 7148 28134 7168
rect 28078 7112 28134 7148
rect 27618 4428 27620 4448
rect 27620 4428 27672 4448
rect 27672 4428 27674 4448
rect 27618 4392 27674 4428
rect 27894 4256 27950 4312
rect 26698 3168 26754 3224
rect 28538 7812 28594 7848
rect 28538 7792 28540 7812
rect 28540 7792 28592 7812
rect 28592 7792 28594 7812
rect 28446 7692 28448 7712
rect 28448 7692 28500 7712
rect 28500 7692 28502 7712
rect 28446 7656 28502 7692
rect 26606 2796 26608 2816
rect 26608 2796 26660 2816
rect 26660 2796 26662 2816
rect 26606 2760 26662 2796
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36726 38800 36782 38856
rect 29274 11756 29330 11792
rect 29274 11736 29276 11756
rect 29276 11736 29328 11756
rect 29328 11736 29330 11756
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 38198 37440 38254 37496
rect 29090 8336 29146 8392
rect 29182 8200 29238 8256
rect 28998 8064 29054 8120
rect 29090 7384 29146 7440
rect 28630 5888 28686 5944
rect 28814 6160 28870 6216
rect 28722 4800 28778 4856
rect 29182 6604 29184 6624
rect 29184 6604 29236 6624
rect 29236 6604 29238 6624
rect 29182 6568 29238 6604
rect 29366 8472 29422 8528
rect 29090 4936 29146 4992
rect 29182 3984 29238 4040
rect 29734 4664 29790 4720
rect 29550 4392 29606 4448
rect 30562 10104 30618 10160
rect 30378 8880 30434 8936
rect 30470 8608 30526 8664
rect 30470 6704 30526 6760
rect 30562 6332 30564 6352
rect 30564 6332 30616 6352
rect 30616 6332 30618 6352
rect 30562 6296 30618 6332
rect 30562 6024 30618 6080
rect 30010 4800 30066 4856
rect 30930 8780 30932 8800
rect 30932 8780 30984 8800
rect 30984 8780 30986 8800
rect 30930 8744 30986 8780
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 31482 11600 31538 11656
rect 31022 7268 31078 7304
rect 31022 7248 31024 7268
rect 31024 7248 31076 7268
rect 31076 7248 31078 7268
rect 31022 6976 31078 7032
rect 31206 6604 31208 6624
rect 31208 6604 31260 6624
rect 31260 6604 31262 6624
rect 31206 6568 31262 6604
rect 32402 9968 32458 10024
rect 31758 7928 31814 7984
rect 31758 5616 31814 5672
rect 30654 4392 30710 4448
rect 30746 3712 30802 3768
rect 29734 3304 29790 3360
rect 31206 3576 31262 3632
rect 31574 3168 31630 3224
rect 31666 2216 31722 2272
rect 32862 6604 32864 6624
rect 32864 6604 32916 6624
rect 32916 6604 32918 6624
rect 32862 6568 32918 6604
rect 32402 5092 32458 5128
rect 32402 5072 32404 5092
rect 32404 5072 32456 5092
rect 32456 5072 32458 5092
rect 32402 4548 32458 4584
rect 32402 4528 32404 4548
rect 32404 4528 32456 4548
rect 32456 4528 32458 4548
rect 32402 3884 32404 3904
rect 32404 3884 32456 3904
rect 32456 3884 32458 3904
rect 32402 3848 32458 3884
rect 32402 2916 32458 2952
rect 32402 2896 32404 2916
rect 32404 2896 32456 2916
rect 32456 2896 32458 2916
rect 32494 2488 32550 2544
rect 31758 1808 31814 1864
rect 33230 5344 33286 5400
rect 33046 5208 33102 5264
rect 32678 2352 32734 2408
rect 33322 3304 33378 3360
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 33690 3440 33746 3496
rect 33690 3068 33692 3088
rect 33692 3068 33744 3088
rect 33744 3068 33746 3088
rect 33690 3032 33746 3068
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34150 5364 34206 5400
rect 34150 5344 34152 5364
rect 34152 5344 34204 5364
rect 34204 5344 34206 5364
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 34518 2624 34574 2680
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 33360 38254 33416
rect 38198 32000 38254 32056
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38198 28600 38254 28656
rect 38290 26560 38346 26616
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 23160 38254 23216
rect 38198 21120 38254 21176
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 38290 15700 38346 15736
rect 38290 15680 38292 15700
rect 38292 15680 38344 15700
rect 38344 15680 38346 15700
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38290 12316 38292 12336
rect 38292 12316 38344 12336
rect 38344 12316 38346 12336
rect 38290 12280 38346 12316
rect 38290 10920 38346 10976
rect 38198 8880 38254 8936
rect 38290 6876 38292 6896
rect 38292 6876 38344 6896
rect 38344 6876 38346 6896
rect 38290 6840 38346 6876
rect 38198 5480 38254 5536
rect 33230 1944 33286 2000
rect 37646 2080 37702 2136
rect 38198 3440 38254 3496
rect 38290 40 38346 96
<< metal3 >>
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 36721 38858 36787 38861
rect 39200 38858 39800 38888
rect 36721 38856 39800 38858
rect 36721 38800 36726 38856
rect 36782 38800 39800 38856
rect 36721 38798 39800 38800
rect 36721 38795 36787 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38193 37498 38259 37501
rect 39200 37498 39800 37528
rect 38193 37496 39800 37498
rect 38193 37440 38198 37496
rect 38254 37440 39800 37496
rect 38193 37438 39800 37440
rect 38193 37435 38259 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1669 36818 1735 36821
rect 200 36816 1735 36818
rect 200 36760 1674 36816
rect 1730 36760 1735 36816
rect 200 36758 1735 36760
rect 200 36728 800 36758
rect 1669 36755 1735 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1669 33418 1735 33421
rect 200 33416 1735 33418
rect 200 33360 1674 33416
rect 1730 33360 1735 33416
rect 200 33358 1735 33360
rect 200 33328 800 33358
rect 1669 33355 1735 33358
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 10501 31786 10567 31789
rect 16430 31786 16436 31788
rect 10501 31784 16436 31786
rect 10501 31728 10506 31784
rect 10562 31728 16436 31784
rect 10501 31726 16436 31728
rect 10501 31723 10567 31726
rect 16430 31724 16436 31726
rect 16500 31724 16506 31788
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1577 31378 1643 31381
rect 200 31376 1643 31378
rect 200 31320 1582 31376
rect 1638 31320 1643 31376
rect 200 31318 1643 31320
rect 200 31288 800 31318
rect 1577 31315 1643 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 200 30018 800 30048
rect 1577 30018 1643 30021
rect 200 30016 1643 30018
rect 200 29960 1582 30016
rect 1638 29960 1643 30016
rect 200 29958 1643 29960
rect 200 29928 800 29958
rect 1577 29955 1643 29958
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1669 27978 1735 27981
rect 200 27976 1735 27978
rect 200 27920 1674 27976
rect 1730 27920 1735 27976
rect 200 27918 1735 27920
rect 200 27888 800 27918
rect 1669 27915 1735 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 17125 26890 17191 26893
rect 27286 26890 27292 26892
rect 17125 26888 27292 26890
rect 17125 26832 17130 26888
rect 17186 26832 27292 26888
rect 17125 26830 27292 26832
rect 17125 26827 17191 26830
rect 27286 26828 27292 26830
rect 27356 26828 27362 26892
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1669 24578 1735 24581
rect 200 24576 1735 24578
rect 200 24520 1674 24576
rect 1730 24520 1735 24576
rect 200 24518 1735 24520
rect 200 24488 800 24518
rect 1669 24515 1735 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 38193 23218 38259 23221
rect 39200 23218 39800 23248
rect 38193 23216 39800 23218
rect 38193 23160 38198 23216
rect 38254 23160 39800 23216
rect 38193 23158 39800 23160
rect 38193 23155 38259 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1577 21178 1643 21181
rect 200 21176 1643 21178
rect 200 21120 1582 21176
rect 1638 21120 1643 21176
rect 200 21118 1643 21120
rect 200 21088 800 21118
rect 1577 21115 1643 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1577 19138 1643 19141
rect 200 19136 1643 19138
rect 200 19080 1582 19136
rect 1638 19080 1643 19136
rect 200 19078 1643 19080
rect 200 19048 800 19078
rect 1577 19075 1643 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1669 17778 1735 17781
rect 200 17776 1735 17778
rect 200 17720 1674 17776
rect 1730 17720 1735 17776
rect 200 17718 1735 17720
rect 200 17688 800 17718
rect 1669 17715 1735 17718
rect 39200 17688 39800 17808
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 24945 16282 25011 16285
rect 27245 16282 27311 16285
rect 24945 16280 27311 16282
rect 24945 16224 24950 16280
rect 25006 16224 27250 16280
rect 27306 16224 27311 16280
rect 24945 16222 27311 16224
rect 24945 16219 25011 16222
rect 27245 16219 27311 16222
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 16205 14650 16271 14653
rect 21541 14650 21607 14653
rect 16205 14648 21607 14650
rect 16205 14592 16210 14648
rect 16266 14592 21546 14648
rect 21602 14592 21607 14648
rect 16205 14590 21607 14592
rect 16205 14587 16271 14590
rect 21541 14587 21607 14590
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 13629 13970 13695 13973
rect 17217 13970 17283 13973
rect 13629 13968 17283 13970
rect 13629 13912 13634 13968
rect 13690 13912 17222 13968
rect 17278 13912 17283 13968
rect 13629 13910 17283 13912
rect 13629 13907 13695 13910
rect 17217 13907 17283 13910
rect 200 13698 800 13728
rect 1669 13698 1735 13701
rect 200 13696 1735 13698
rect 200 13640 1674 13696
rect 1730 13640 1735 13696
rect 200 13638 1735 13640
rect 200 13608 800 13638
rect 1669 13635 1735 13638
rect 13261 13698 13327 13701
rect 13721 13698 13787 13701
rect 19793 13698 19859 13701
rect 13261 13696 19859 13698
rect 13261 13640 13266 13696
rect 13322 13640 13726 13696
rect 13782 13640 19798 13696
rect 19854 13640 19859 13696
rect 13261 13638 19859 13640
rect 13261 13635 13327 13638
rect 13721 13635 13787 13638
rect 19793 13635 19859 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 13721 13562 13787 13565
rect 16573 13562 16639 13565
rect 13721 13560 16639 13562
rect 13721 13504 13726 13560
rect 13782 13504 16578 13560
rect 16634 13504 16639 13560
rect 13721 13502 16639 13504
rect 13721 13499 13787 13502
rect 16573 13499 16639 13502
rect 12893 13154 12959 13157
rect 15193 13154 15259 13157
rect 12893 13152 15259 13154
rect 12893 13096 12898 13152
rect 12954 13096 15198 13152
rect 15254 13096 15259 13152
rect 12893 13094 15259 13096
rect 12893 13091 12959 13094
rect 15193 13091 15259 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 13169 12746 13235 12749
rect 17033 12746 17099 12749
rect 13169 12744 17099 12746
rect 13169 12688 13174 12744
rect 13230 12688 17038 12744
rect 17094 12688 17099 12744
rect 13169 12686 17099 12688
rect 13169 12683 13235 12686
rect 17033 12683 17099 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 38285 12338 38351 12341
rect 39200 12338 39800 12368
rect 38285 12336 39800 12338
rect 38285 12280 38290 12336
rect 38346 12280 39800 12336
rect 38285 12278 39800 12280
rect 38285 12275 38351 12278
rect 39200 12248 39800 12278
rect 16481 12204 16547 12205
rect 16430 12202 16436 12204
rect 16390 12142 16436 12202
rect 16500 12200 16547 12204
rect 16542 12144 16547 12200
rect 16430 12140 16436 12142
rect 16500 12140 16547 12144
rect 19374 12140 19380 12204
rect 19444 12202 19450 12204
rect 20069 12202 20135 12205
rect 19444 12200 20135 12202
rect 19444 12144 20074 12200
rect 20130 12144 20135 12200
rect 19444 12142 20135 12144
rect 19444 12140 19450 12142
rect 16481 12139 16547 12140
rect 20069 12139 20135 12142
rect 23749 12202 23815 12205
rect 26325 12202 26391 12205
rect 28073 12202 28139 12205
rect 23749 12200 28139 12202
rect 23749 12144 23754 12200
rect 23810 12144 26330 12200
rect 26386 12144 28078 12200
rect 28134 12144 28139 12200
rect 23749 12142 28139 12144
rect 23749 12139 23815 12142
rect 26325 12139 26391 12142
rect 28073 12139 28139 12142
rect 20805 12066 20871 12069
rect 24025 12066 24091 12069
rect 27521 12066 27587 12069
rect 20805 12064 27587 12066
rect 20805 12008 20810 12064
rect 20866 12008 24030 12064
rect 24086 12008 27526 12064
rect 27582 12008 27587 12064
rect 20805 12006 27587 12008
rect 20805 12003 20871 12006
rect 24025 12003 24091 12006
rect 27521 12003 27587 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 9765 11794 9831 11797
rect 15837 11794 15903 11797
rect 9765 11792 15903 11794
rect 9765 11736 9770 11792
rect 9826 11736 15842 11792
rect 15898 11736 15903 11792
rect 9765 11734 15903 11736
rect 9765 11731 9831 11734
rect 15837 11731 15903 11734
rect 16113 11794 16179 11797
rect 29269 11794 29335 11797
rect 16113 11792 29335 11794
rect 16113 11736 16118 11792
rect 16174 11736 29274 11792
rect 29330 11736 29335 11792
rect 16113 11734 29335 11736
rect 16113 11731 16179 11734
rect 29269 11731 29335 11734
rect 17861 11658 17927 11661
rect 22461 11658 22527 11661
rect 31477 11658 31543 11661
rect 17861 11656 31543 11658
rect 17861 11600 17866 11656
rect 17922 11600 22466 11656
rect 22522 11600 31482 11656
rect 31538 11600 31543 11656
rect 17861 11598 31543 11600
rect 17861 11595 17927 11598
rect 22461 11595 22527 11598
rect 31477 11595 31543 11598
rect 25313 11522 25379 11525
rect 27245 11522 27311 11525
rect 25313 11520 27311 11522
rect 25313 11464 25318 11520
rect 25374 11464 27250 11520
rect 27306 11464 27311 11520
rect 25313 11462 27311 11464
rect 25313 11459 25379 11462
rect 27245 11459 27311 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 13813 11386 13879 11389
rect 18229 11386 18295 11389
rect 13813 11384 18295 11386
rect 13813 11328 13818 11384
rect 13874 11328 18234 11384
rect 18290 11328 18295 11384
rect 13813 11326 18295 11328
rect 13813 11323 13879 11326
rect 18229 11323 18295 11326
rect 11053 11250 11119 11253
rect 14273 11250 14339 11253
rect 11053 11248 14339 11250
rect 11053 11192 11058 11248
rect 11114 11192 14278 11248
rect 14334 11192 14339 11248
rect 11053 11190 14339 11192
rect 11053 11187 11119 11190
rect 14273 11187 14339 11190
rect 27981 10978 28047 10981
rect 28625 10978 28691 10981
rect 27981 10976 28691 10978
rect 27981 10920 27986 10976
rect 28042 10920 28630 10976
rect 28686 10920 28691 10976
rect 27981 10918 28691 10920
rect 27981 10915 28047 10918
rect 28625 10915 28691 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 14181 10842 14247 10845
rect 15009 10842 15075 10845
rect 18321 10842 18387 10845
rect 14181 10840 18387 10842
rect 14181 10784 14186 10840
rect 14242 10784 15014 10840
rect 15070 10784 18326 10840
rect 18382 10784 18387 10840
rect 14181 10782 18387 10784
rect 14181 10779 14247 10782
rect 15009 10779 15075 10782
rect 18321 10779 18387 10782
rect 14825 10706 14891 10709
rect 20989 10706 21055 10709
rect 14825 10704 21055 10706
rect 14825 10648 14830 10704
rect 14886 10648 20994 10704
rect 21050 10648 21055 10704
rect 14825 10646 21055 10648
rect 14825 10643 14891 10646
rect 20989 10643 21055 10646
rect 10961 10570 11027 10573
rect 15561 10570 15627 10573
rect 10961 10568 15627 10570
rect 10961 10512 10966 10568
rect 11022 10512 15566 10568
rect 15622 10512 15627 10568
rect 10961 10510 15627 10512
rect 10961 10507 11027 10510
rect 15561 10507 15627 10510
rect 19425 10570 19491 10573
rect 21265 10570 21331 10573
rect 19425 10568 21331 10570
rect 19425 10512 19430 10568
rect 19486 10512 21270 10568
rect 21326 10512 21331 10568
rect 19425 10510 21331 10512
rect 19425 10507 19491 10510
rect 21265 10507 21331 10510
rect 15009 10434 15075 10437
rect 16757 10434 16823 10437
rect 15009 10432 16823 10434
rect 15009 10376 15014 10432
rect 15070 10376 16762 10432
rect 16818 10376 16823 10432
rect 15009 10374 16823 10376
rect 15009 10371 15075 10374
rect 16757 10371 16823 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 19333 10298 19399 10301
rect 25865 10298 25931 10301
rect 19333 10296 25931 10298
rect 19333 10240 19338 10296
rect 19394 10240 25870 10296
rect 25926 10240 25931 10296
rect 19333 10238 25931 10240
rect 19333 10235 19399 10238
rect 25865 10235 25931 10238
rect 19241 10162 19307 10165
rect 30557 10162 30623 10165
rect 19241 10160 30623 10162
rect 19241 10104 19246 10160
rect 19302 10104 30562 10160
rect 30618 10104 30623 10160
rect 19241 10102 30623 10104
rect 19241 10099 19307 10102
rect 30557 10099 30623 10102
rect 15101 10026 15167 10029
rect 32397 10026 32463 10029
rect 15101 10024 32463 10026
rect 15101 9968 15106 10024
rect 15162 9968 32402 10024
rect 32458 9968 32463 10024
rect 15101 9966 32463 9968
rect 15101 9963 15167 9966
rect 32397 9963 32463 9966
rect 19333 9892 19399 9893
rect 19333 9888 19380 9892
rect 19444 9890 19450 9892
rect 19333 9832 19338 9888
rect 19333 9828 19380 9832
rect 19444 9830 19490 9890
rect 19444 9828 19450 9830
rect 19333 9827 19399 9828
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 19333 9754 19399 9757
rect 20621 9754 20687 9757
rect 19333 9752 19442 9754
rect 19333 9696 19338 9752
rect 19394 9696 19442 9752
rect 19333 9691 19442 9696
rect 19382 9690 19442 9691
rect 20118 9752 20687 9754
rect 20118 9696 20626 9752
rect 20682 9696 20687 9752
rect 20118 9694 20687 9696
rect 20118 9690 20178 9694
rect 20621 9691 20687 9694
rect 19382 9630 20178 9690
rect 9857 9618 9923 9621
rect 15101 9618 15167 9621
rect 9857 9616 15167 9618
rect 9857 9560 9862 9616
rect 9918 9560 15106 9616
rect 15162 9560 15167 9616
rect 9857 9558 15167 9560
rect 9857 9555 9923 9558
rect 15101 9555 15167 9558
rect 9305 9482 9371 9485
rect 14733 9482 14799 9485
rect 9305 9480 14799 9482
rect 9305 9424 9310 9480
rect 9366 9424 14738 9480
rect 14794 9424 14799 9480
rect 9305 9422 14799 9424
rect 9305 9419 9371 9422
rect 14733 9419 14799 9422
rect 15377 9482 15443 9485
rect 15653 9482 15719 9485
rect 15377 9480 15719 9482
rect 15377 9424 15382 9480
rect 15438 9424 15658 9480
rect 15714 9424 15719 9480
rect 15377 9422 15719 9424
rect 15377 9419 15443 9422
rect 15653 9419 15719 9422
rect 26601 9482 26667 9485
rect 28165 9482 28231 9485
rect 26601 9480 28231 9482
rect 26601 9424 26606 9480
rect 26662 9424 28170 9480
rect 28226 9424 28231 9480
rect 26601 9422 28231 9424
rect 26601 9419 26667 9422
rect 28165 9419 28231 9422
rect 26509 9346 26575 9349
rect 27797 9346 27863 9349
rect 26509 9344 27863 9346
rect 26509 9288 26514 9344
rect 26570 9288 27802 9344
rect 27858 9288 27863 9344
rect 26509 9286 27863 9288
rect 26509 9283 26575 9286
rect 27797 9283 27863 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 24761 9210 24827 9213
rect 27889 9210 27955 9213
rect 24761 9208 27955 9210
rect 24761 9152 24766 9208
rect 24822 9152 27894 9208
rect 27950 9152 27955 9208
rect 24761 9150 27955 9152
rect 24761 9147 24827 9150
rect 27889 9147 27955 9150
rect 14549 9074 14615 9077
rect 15101 9074 15167 9077
rect 14549 9072 15167 9074
rect 14549 9016 14554 9072
rect 14610 9016 15106 9072
rect 15162 9016 15167 9072
rect 14549 9014 15167 9016
rect 14549 9011 14615 9014
rect 15101 9011 15167 9014
rect 26141 9074 26207 9077
rect 28809 9074 28875 9077
rect 26141 9072 28875 9074
rect 26141 9016 26146 9072
rect 26202 9016 28814 9072
rect 28870 9016 28875 9072
rect 26141 9014 28875 9016
rect 26141 9011 26207 9014
rect 28809 9011 28875 9014
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 14365 8938 14431 8941
rect 15929 8938 15995 8941
rect 14365 8936 15995 8938
rect 14365 8880 14370 8936
rect 14426 8880 15934 8936
rect 15990 8880 15995 8936
rect 14365 8878 15995 8880
rect 14365 8875 14431 8878
rect 15929 8875 15995 8878
rect 16481 8938 16547 8941
rect 30373 8938 30439 8941
rect 16481 8936 30439 8938
rect 16481 8880 16486 8936
rect 16542 8880 30378 8936
rect 30434 8880 30439 8936
rect 16481 8878 30439 8880
rect 16481 8875 16547 8878
rect 30373 8875 30439 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 15101 8802 15167 8805
rect 18137 8802 18203 8805
rect 15101 8800 18203 8802
rect 15101 8744 15106 8800
rect 15162 8744 18142 8800
rect 18198 8744 18203 8800
rect 15101 8742 18203 8744
rect 15101 8739 15167 8742
rect 18137 8739 18203 8742
rect 23749 8802 23815 8805
rect 30925 8802 30991 8805
rect 23749 8800 30991 8802
rect 23749 8744 23754 8800
rect 23810 8744 30930 8800
rect 30986 8744 30991 8800
rect 23749 8742 30991 8744
rect 23749 8739 23815 8742
rect 30925 8739 30991 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 20713 8666 20779 8669
rect 30465 8666 30531 8669
rect 20713 8664 30531 8666
rect 20713 8608 20718 8664
rect 20774 8608 30470 8664
rect 30526 8608 30531 8664
rect 20713 8606 30531 8608
rect 20713 8603 20779 8606
rect 30465 8603 30531 8606
rect 27521 8530 27587 8533
rect 28758 8530 28764 8532
rect 27521 8528 28764 8530
rect 27521 8472 27526 8528
rect 27582 8472 28764 8528
rect 27521 8470 28764 8472
rect 27521 8467 27587 8470
rect 28758 8468 28764 8470
rect 28828 8530 28834 8532
rect 29361 8530 29427 8533
rect 28828 8528 29427 8530
rect 28828 8472 29366 8528
rect 29422 8472 29427 8528
rect 28828 8470 29427 8472
rect 28828 8468 28834 8470
rect 29361 8467 29427 8470
rect 29085 8394 29151 8397
rect 26558 8392 29151 8394
rect 26558 8336 29090 8392
rect 29146 8336 29151 8392
rect 26558 8334 29151 8336
rect 26558 8261 26618 8334
rect 29085 8331 29151 8334
rect 26558 8256 26667 8261
rect 26558 8200 26606 8256
rect 26662 8200 26667 8256
rect 26558 8198 26667 8200
rect 26601 8195 26667 8198
rect 26785 8258 26851 8261
rect 29177 8258 29243 8261
rect 26785 8256 29243 8258
rect 26785 8200 26790 8256
rect 26846 8200 29182 8256
rect 29238 8200 29243 8256
rect 26785 8198 29243 8200
rect 26785 8195 26851 8198
rect 29177 8195 29243 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 24761 8122 24827 8125
rect 28993 8122 29059 8125
rect 24761 8120 29059 8122
rect 24761 8064 24766 8120
rect 24822 8064 28998 8120
rect 29054 8064 29059 8120
rect 24761 8062 29059 8064
rect 24761 8059 24827 8062
rect 28993 8059 29059 8062
rect 25405 7986 25471 7989
rect 31753 7986 31819 7989
rect 25405 7984 31819 7986
rect 25405 7928 25410 7984
rect 25466 7928 31758 7984
rect 31814 7928 31819 7984
rect 25405 7926 31819 7928
rect 25405 7923 25471 7926
rect 31753 7923 31819 7926
rect 27061 7850 27127 7853
rect 28533 7850 28599 7853
rect 27061 7848 28599 7850
rect 27061 7792 27066 7848
rect 27122 7792 28538 7848
rect 28594 7792 28599 7848
rect 27061 7790 28599 7792
rect 27061 7787 27127 7790
rect 28533 7787 28599 7790
rect 21449 7714 21515 7717
rect 28441 7714 28507 7717
rect 21449 7712 28507 7714
rect 21449 7656 21454 7712
rect 21510 7656 28446 7712
rect 28502 7656 28507 7712
rect 21449 7654 28507 7656
rect 21449 7651 21515 7654
rect 28441 7651 28507 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 20529 7578 20595 7581
rect 22369 7578 22435 7581
rect 20529 7576 22435 7578
rect 20529 7520 20534 7576
rect 20590 7520 22374 7576
rect 22430 7520 22435 7576
rect 20529 7518 22435 7520
rect 20529 7515 20595 7518
rect 22369 7515 22435 7518
rect 12249 7442 12315 7445
rect 29085 7442 29151 7445
rect 12249 7440 29151 7442
rect 12249 7384 12254 7440
rect 12310 7384 29090 7440
rect 29146 7384 29151 7440
rect 12249 7382 29151 7384
rect 12249 7379 12315 7382
rect 29085 7379 29151 7382
rect 14733 7306 14799 7309
rect 31017 7306 31083 7309
rect 14733 7304 31083 7306
rect 14733 7248 14738 7304
rect 14794 7248 31022 7304
rect 31078 7248 31083 7304
rect 14733 7246 31083 7248
rect 14733 7243 14799 7246
rect 31017 7243 31083 7246
rect 20897 7170 20963 7173
rect 28073 7170 28139 7173
rect 20897 7168 28139 7170
rect 20897 7112 20902 7168
rect 20958 7112 28078 7168
rect 28134 7112 28139 7168
rect 20897 7110 28139 7112
rect 20897 7107 20963 7110
rect 28073 7107 28139 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 20713 7034 20779 7037
rect 31017 7034 31083 7037
rect 20713 7032 31083 7034
rect 20713 6976 20718 7032
rect 20774 6976 31022 7032
rect 31078 6976 31083 7032
rect 20713 6974 31083 6976
rect 20713 6971 20779 6974
rect 31017 6971 31083 6974
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 10869 6898 10935 6901
rect 14733 6898 14799 6901
rect 10869 6896 14799 6898
rect 10869 6840 10874 6896
rect 10930 6840 14738 6896
rect 14794 6840 14799 6896
rect 10869 6838 14799 6840
rect 10869 6835 10935 6838
rect 14733 6835 14799 6838
rect 20621 6898 20687 6901
rect 22277 6898 22343 6901
rect 20621 6896 22343 6898
rect 20621 6840 20626 6896
rect 20682 6840 22282 6896
rect 22338 6840 22343 6896
rect 20621 6838 22343 6840
rect 20621 6835 20687 6838
rect 22277 6835 22343 6838
rect 23289 6898 23355 6901
rect 26785 6898 26851 6901
rect 23289 6896 26851 6898
rect 23289 6840 23294 6896
rect 23350 6840 26790 6896
rect 26846 6840 26851 6896
rect 23289 6838 26851 6840
rect 23289 6835 23355 6838
rect 26785 6835 26851 6838
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 12433 6762 12499 6765
rect 14457 6762 14523 6765
rect 12433 6760 14523 6762
rect 12433 6704 12438 6760
rect 12494 6704 14462 6760
rect 14518 6704 14523 6760
rect 12433 6702 14523 6704
rect 12433 6699 12499 6702
rect 14457 6699 14523 6702
rect 25497 6762 25563 6765
rect 30465 6762 30531 6765
rect 25497 6760 30531 6762
rect 25497 6704 25502 6760
rect 25558 6704 30470 6760
rect 30526 6704 30531 6760
rect 25497 6702 30531 6704
rect 25497 6699 25563 6702
rect 30465 6699 30531 6702
rect 20161 6626 20227 6629
rect 27797 6626 27863 6629
rect 20161 6624 27863 6626
rect 20161 6568 20166 6624
rect 20222 6568 27802 6624
rect 27858 6568 27863 6624
rect 20161 6566 27863 6568
rect 20161 6563 20227 6566
rect 27797 6563 27863 6566
rect 29177 6626 29243 6629
rect 31201 6626 31267 6629
rect 32857 6626 32923 6629
rect 29177 6624 31267 6626
rect 29177 6568 29182 6624
rect 29238 6568 31206 6624
rect 31262 6568 31267 6624
rect 29177 6566 31267 6568
rect 29177 6563 29243 6566
rect 31201 6563 31267 6566
rect 31710 6624 32923 6626
rect 31710 6568 32862 6624
rect 32918 6568 32923 6624
rect 31710 6566 32923 6568
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 22277 6490 22343 6493
rect 27613 6490 27679 6493
rect 22277 6488 27679 6490
rect 22277 6432 22282 6488
rect 22338 6432 27618 6488
rect 27674 6432 27679 6488
rect 22277 6430 27679 6432
rect 22277 6427 22343 6430
rect 27613 6427 27679 6430
rect 17585 6354 17651 6357
rect 30557 6354 30623 6357
rect 17585 6352 30623 6354
rect 17585 6296 17590 6352
rect 17646 6296 30562 6352
rect 30618 6296 30623 6352
rect 17585 6294 30623 6296
rect 17585 6291 17651 6294
rect 30557 6291 30623 6294
rect 21817 6218 21883 6221
rect 23473 6218 23539 6221
rect 24945 6218 25011 6221
rect 21817 6216 25011 6218
rect 21817 6160 21822 6216
rect 21878 6160 23478 6216
rect 23534 6160 24950 6216
rect 25006 6160 25011 6216
rect 21817 6158 25011 6160
rect 21817 6155 21883 6158
rect 23473 6155 23539 6158
rect 24945 6155 25011 6158
rect 26693 6218 26759 6221
rect 28809 6218 28875 6221
rect 31710 6218 31770 6566
rect 32857 6563 32923 6566
rect 26693 6216 31770 6218
rect 26693 6160 26698 6216
rect 26754 6160 28814 6216
rect 28870 6160 31770 6216
rect 26693 6158 31770 6160
rect 26693 6155 26759 6158
rect 28809 6155 28875 6158
rect 22185 6082 22251 6085
rect 30557 6082 30623 6085
rect 22185 6080 30623 6082
rect 22185 6024 22190 6080
rect 22246 6024 30562 6080
rect 30618 6024 30623 6080
rect 22185 6022 30623 6024
rect 22185 6019 22251 6022
rect 30557 6019 30623 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 20713 5946 20779 5949
rect 28625 5946 28691 5949
rect 20713 5944 28691 5946
rect 20713 5888 20718 5944
rect 20774 5888 28630 5944
rect 28686 5888 28691 5944
rect 20713 5886 28691 5888
rect 20713 5883 20779 5886
rect 28625 5883 28691 5886
rect 13629 5810 13695 5813
rect 25773 5810 25839 5813
rect 27705 5810 27771 5813
rect 13629 5808 22110 5810
rect 13629 5752 13634 5808
rect 13690 5752 22110 5808
rect 13629 5750 22110 5752
rect 13629 5747 13695 5750
rect 9489 5674 9555 5677
rect 15009 5674 15075 5677
rect 9489 5672 15075 5674
rect 9489 5616 9494 5672
rect 9550 5616 15014 5672
rect 15070 5616 15075 5672
rect 9489 5614 15075 5616
rect 9489 5611 9555 5614
rect 15009 5611 15075 5614
rect 16205 5674 16271 5677
rect 20253 5674 20319 5677
rect 16205 5672 20319 5674
rect 16205 5616 16210 5672
rect 16266 5616 20258 5672
rect 20314 5616 20319 5672
rect 16205 5614 20319 5616
rect 22050 5674 22110 5750
rect 25773 5808 27771 5810
rect 25773 5752 25778 5808
rect 25834 5752 27710 5808
rect 27766 5752 27771 5808
rect 25773 5750 27771 5752
rect 25773 5747 25839 5750
rect 27705 5747 27771 5750
rect 31753 5674 31819 5677
rect 22050 5672 31819 5674
rect 22050 5616 31758 5672
rect 31814 5616 31819 5672
rect 22050 5614 31819 5616
rect 16205 5611 16271 5614
rect 20253 5611 20319 5614
rect 31753 5611 31819 5614
rect 27245 5540 27311 5541
rect 27245 5536 27292 5540
rect 27356 5538 27362 5540
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 27245 5480 27250 5536
rect 27245 5476 27292 5480
rect 27356 5478 27402 5538
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 27356 5476 27362 5478
rect 27245 5475 27311 5476
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 9765 5402 9831 5405
rect 14733 5402 14799 5405
rect 9765 5400 14799 5402
rect 9765 5344 9770 5400
rect 9826 5344 14738 5400
rect 14794 5344 14799 5400
rect 9765 5342 14799 5344
rect 9765 5339 9831 5342
rect 14733 5339 14799 5342
rect 25865 5402 25931 5405
rect 33225 5402 33291 5405
rect 34145 5402 34211 5405
rect 25865 5400 34211 5402
rect 25865 5344 25870 5400
rect 25926 5344 33230 5400
rect 33286 5344 34150 5400
rect 34206 5344 34211 5400
rect 25865 5342 34211 5344
rect 25865 5339 25931 5342
rect 33225 5339 33291 5342
rect 34145 5339 34211 5342
rect 15009 5266 15075 5269
rect 33041 5266 33107 5269
rect 15009 5264 33107 5266
rect 15009 5208 15014 5264
rect 15070 5208 33046 5264
rect 33102 5208 33107 5264
rect 15009 5206 33107 5208
rect 15009 5203 15075 5206
rect 33041 5203 33107 5206
rect 14273 5130 14339 5133
rect 15377 5130 15443 5133
rect 14273 5128 15443 5130
rect 14273 5072 14278 5128
rect 14334 5072 15382 5128
rect 15438 5072 15443 5128
rect 14273 5070 15443 5072
rect 14273 5067 14339 5070
rect 15377 5067 15443 5070
rect 17861 5130 17927 5133
rect 32397 5130 32463 5133
rect 17861 5128 32463 5130
rect 17861 5072 17866 5128
rect 17922 5072 32402 5128
rect 32458 5072 32463 5128
rect 17861 5070 32463 5072
rect 17861 5067 17927 5070
rect 32397 5067 32463 5070
rect 19333 4994 19399 4997
rect 29085 4994 29151 4997
rect 19333 4992 29151 4994
rect 19333 4936 19338 4992
rect 19394 4936 29090 4992
rect 29146 4936 29151 4992
rect 19333 4934 29151 4936
rect 19333 4931 19399 4934
rect 29085 4931 29151 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1577 4858 1643 4861
rect 200 4856 1643 4858
rect 200 4800 1582 4856
rect 1638 4800 1643 4856
rect 200 4798 1643 4800
rect 200 4768 800 4798
rect 1577 4795 1643 4798
rect 10409 4858 10475 4861
rect 17309 4858 17375 4861
rect 10409 4856 17375 4858
rect 10409 4800 10414 4856
rect 10470 4800 17314 4856
rect 17370 4800 17375 4856
rect 10409 4798 17375 4800
rect 10409 4795 10475 4798
rect 17309 4795 17375 4798
rect 24301 4858 24367 4861
rect 28717 4858 28783 4861
rect 30005 4858 30071 4861
rect 24301 4856 30071 4858
rect 24301 4800 24306 4856
rect 24362 4800 28722 4856
rect 28778 4800 30010 4856
rect 30066 4800 30071 4856
rect 24301 4798 30071 4800
rect 24301 4795 24367 4798
rect 28717 4795 28783 4798
rect 30005 4795 30071 4798
rect 14273 4722 14339 4725
rect 14825 4722 14891 4725
rect 14273 4720 14891 4722
rect 14273 4664 14278 4720
rect 14334 4664 14830 4720
rect 14886 4664 14891 4720
rect 14273 4662 14891 4664
rect 14273 4659 14339 4662
rect 14825 4659 14891 4662
rect 19977 4722 20043 4725
rect 28758 4722 28764 4724
rect 19977 4720 28764 4722
rect 19977 4664 19982 4720
rect 20038 4664 28764 4720
rect 19977 4662 28764 4664
rect 19977 4659 20043 4662
rect 28758 4660 28764 4662
rect 28828 4722 28834 4724
rect 29729 4722 29795 4725
rect 28828 4720 29795 4722
rect 28828 4664 29734 4720
rect 29790 4664 29795 4720
rect 28828 4662 29795 4664
rect 28828 4660 28834 4662
rect 29729 4659 29795 4662
rect 22645 4586 22711 4589
rect 32397 4586 32463 4589
rect 22645 4584 32463 4586
rect 22645 4528 22650 4584
rect 22706 4528 32402 4584
rect 32458 4528 32463 4584
rect 22645 4526 32463 4528
rect 22645 4523 22711 4526
rect 32397 4523 32463 4526
rect 24117 4450 24183 4453
rect 27613 4450 27679 4453
rect 24117 4448 27679 4450
rect 24117 4392 24122 4448
rect 24178 4392 27618 4448
rect 27674 4392 27679 4448
rect 24117 4390 27679 4392
rect 24117 4387 24183 4390
rect 27613 4387 27679 4390
rect 29545 4450 29611 4453
rect 30649 4450 30715 4453
rect 29545 4448 30715 4450
rect 29545 4392 29550 4448
rect 29606 4392 30654 4448
rect 30710 4392 30715 4448
rect 29545 4390 30715 4392
rect 29545 4387 29611 4390
rect 30649 4387 30715 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 24669 4314 24735 4317
rect 27889 4314 27955 4317
rect 24669 4312 27955 4314
rect 24669 4256 24674 4312
rect 24730 4256 27894 4312
rect 27950 4256 27955 4312
rect 24669 4254 27955 4256
rect 24669 4251 24735 4254
rect 27889 4251 27955 4254
rect 12433 4178 12499 4181
rect 20437 4178 20503 4181
rect 22369 4178 22435 4181
rect 12433 4176 22435 4178
rect 12433 4120 12438 4176
rect 12494 4120 20442 4176
rect 20498 4120 22374 4176
rect 22430 4120 22435 4176
rect 12433 4118 22435 4120
rect 12433 4115 12499 4118
rect 20437 4115 20503 4118
rect 22369 4115 22435 4118
rect 12709 4042 12775 4045
rect 17861 4042 17927 4045
rect 12709 4040 17927 4042
rect 12709 3984 12714 4040
rect 12770 3984 17866 4040
rect 17922 3984 17927 4040
rect 12709 3982 17927 3984
rect 12709 3979 12775 3982
rect 17861 3979 17927 3982
rect 22001 4042 22067 4045
rect 29177 4042 29243 4045
rect 22001 4040 29243 4042
rect 22001 3984 22006 4040
rect 22062 3984 29182 4040
rect 29238 3984 29243 4040
rect 22001 3982 29243 3984
rect 22001 3979 22067 3982
rect 29177 3979 29243 3982
rect 13353 3906 13419 3909
rect 19149 3906 19215 3909
rect 13353 3904 19215 3906
rect 13353 3848 13358 3904
rect 13414 3848 19154 3904
rect 19210 3848 19215 3904
rect 13353 3846 19215 3848
rect 13353 3843 13419 3846
rect 19149 3843 19215 3846
rect 23657 3906 23723 3909
rect 32397 3906 32463 3909
rect 23657 3904 32463 3906
rect 23657 3848 23662 3904
rect 23718 3848 32402 3904
rect 32458 3848 32463 3904
rect 23657 3846 32463 3848
rect 23657 3843 23723 3846
rect 32397 3843 32463 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 21909 3770 21975 3773
rect 30741 3770 30807 3773
rect 21909 3768 30807 3770
rect 21909 3712 21914 3768
rect 21970 3712 30746 3768
rect 30802 3712 30807 3768
rect 21909 3710 30807 3712
rect 21909 3707 21975 3710
rect 30741 3707 30807 3710
rect 8109 3634 8175 3637
rect 31201 3634 31267 3637
rect 8109 3632 31267 3634
rect 8109 3576 8114 3632
rect 8170 3576 31206 3632
rect 31262 3576 31267 3632
rect 8109 3574 31267 3576
rect 8109 3571 8175 3574
rect 31201 3571 31267 3574
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 16205 3498 16271 3501
rect 33685 3498 33751 3501
rect 16205 3496 33751 3498
rect 16205 3440 16210 3496
rect 16266 3440 33690 3496
rect 33746 3440 33751 3496
rect 16205 3438 33751 3440
rect 16205 3435 16271 3438
rect 33685 3435 33751 3438
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 29729 3362 29795 3365
rect 33317 3362 33383 3365
rect 29729 3360 33383 3362
rect 29729 3304 29734 3360
rect 29790 3304 33322 3360
rect 33378 3304 33383 3360
rect 29729 3302 33383 3304
rect 29729 3299 29795 3302
rect 33317 3299 33383 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 12065 3226 12131 3229
rect 12617 3226 12683 3229
rect 12065 3224 12683 3226
rect 12065 3168 12070 3224
rect 12126 3168 12622 3224
rect 12678 3168 12683 3224
rect 12065 3166 12683 3168
rect 12065 3163 12131 3166
rect 12617 3163 12683 3166
rect 22093 3226 22159 3229
rect 24025 3226 24091 3229
rect 22093 3224 24091 3226
rect 22093 3168 22098 3224
rect 22154 3168 24030 3224
rect 24086 3168 24091 3224
rect 22093 3166 24091 3168
rect 22093 3163 22159 3166
rect 24025 3163 24091 3166
rect 25405 3226 25471 3229
rect 26693 3226 26759 3229
rect 31569 3226 31635 3229
rect 25405 3224 31635 3226
rect 25405 3168 25410 3224
rect 25466 3168 26698 3224
rect 26754 3168 31574 3224
rect 31630 3168 31635 3224
rect 25405 3166 31635 3168
rect 25405 3163 25471 3166
rect 26693 3163 26759 3166
rect 31569 3163 31635 3166
rect 16113 3090 16179 3093
rect 33685 3090 33751 3093
rect 16113 3088 33751 3090
rect 16113 3032 16118 3088
rect 16174 3032 33690 3088
rect 33746 3032 33751 3088
rect 16113 3030 33751 3032
rect 16113 3027 16179 3030
rect 33685 3027 33751 3030
rect 18965 2954 19031 2957
rect 32397 2954 32463 2957
rect 18965 2952 32463 2954
rect 18965 2896 18970 2952
rect 19026 2896 32402 2952
rect 32458 2896 32463 2952
rect 18965 2894 32463 2896
rect 18965 2891 19031 2894
rect 32397 2891 32463 2894
rect 20621 2818 20687 2821
rect 26601 2818 26667 2821
rect 20621 2816 26667 2818
rect 20621 2760 20626 2816
rect 20682 2760 26606 2816
rect 26662 2760 26667 2816
rect 20621 2758 26667 2760
rect 20621 2755 20687 2758
rect 26601 2755 26667 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 25957 2682 26023 2685
rect 34513 2682 34579 2685
rect 25957 2680 34579 2682
rect 25957 2624 25962 2680
rect 26018 2624 34518 2680
rect 34574 2624 34579 2680
rect 25957 2622 34579 2624
rect 25957 2619 26023 2622
rect 34513 2619 34579 2622
rect 24393 2546 24459 2549
rect 32489 2546 32555 2549
rect 24393 2544 32555 2546
rect 24393 2488 24398 2544
rect 24454 2488 32494 2544
rect 32550 2488 32555 2544
rect 24393 2486 32555 2488
rect 24393 2483 24459 2486
rect 32489 2483 32555 2486
rect 15285 2410 15351 2413
rect 32673 2410 32739 2413
rect 15285 2408 32739 2410
rect 15285 2352 15290 2408
rect 15346 2352 32678 2408
rect 32734 2352 32739 2408
rect 15285 2350 32739 2352
rect 15285 2347 15351 2350
rect 32673 2347 32739 2350
rect 23657 2274 23723 2277
rect 31661 2274 31727 2277
rect 23657 2272 31727 2274
rect 23657 2216 23662 2272
rect 23718 2216 31666 2272
rect 31722 2216 31727 2272
rect 23657 2214 31727 2216
rect 23657 2211 23723 2214
rect 31661 2211 31727 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 37641 2138 37707 2141
rect 39200 2138 39800 2168
rect 37641 2136 39800 2138
rect 37641 2080 37646 2136
rect 37702 2080 39800 2136
rect 37641 2078 39800 2080
rect 37641 2075 37707 2078
rect 39200 2048 39800 2078
rect 19149 2002 19215 2005
rect 33225 2002 33291 2005
rect 19149 2000 33291 2002
rect 19149 1944 19154 2000
rect 19210 1944 33230 2000
rect 33286 1944 33291 2000
rect 19149 1942 33291 1944
rect 19149 1939 19215 1942
rect 33225 1939 33291 1942
rect 17861 1866 17927 1869
rect 31753 1866 31819 1869
rect 17861 1864 31819 1866
rect 17861 1808 17866 1864
rect 17922 1808 31758 1864
rect 31814 1808 31819 1864
rect 17861 1806 31819 1808
rect 17861 1803 17927 1806
rect 31753 1803 31819 1806
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 38285 98 38351 101
rect 39200 98 39800 128
rect 38285 96 39800 98
rect 38285 40 38290 96
rect 38346 40 39800 96
rect 38285 38 39800 40
rect 38285 35 38351 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 16436 31724 16500 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 27292 26828 27356 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 16436 12200 16500 12204
rect 16436 12144 16486 12200
rect 16486 12144 16500 12200
rect 16436 12140 16500 12144
rect 19380 12140 19444 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19380 9888 19444 9892
rect 19380 9832 19394 9888
rect 19394 9832 19444 9888
rect 19380 9828 19444 9832
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 28764 8468 28828 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 27292 5536 27356 5540
rect 27292 5480 27306 5536
rect 27306 5480 27356 5536
rect 27292 5476 27356 5480
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 28764 4660 28828 4724
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 16435 31788 16501 31789
rect 16435 31724 16436 31788
rect 16500 31724 16501 31788
rect 16435 31723 16501 31724
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 16438 12205 16498 31723
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 27291 26892 27357 26893
rect 27291 26828 27292 26892
rect 27356 26828 27357 26892
rect 27291 26827 27357 26828
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 16435 12204 16501 12205
rect 16435 12140 16436 12204
rect 16500 12140 16501 12204
rect 16435 12139 16501 12140
rect 19379 12204 19445 12205
rect 19379 12140 19380 12204
rect 19444 12140 19445 12204
rect 19379 12139 19445 12140
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 19382 9893 19442 12139
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 9892 19445 9893
rect 19379 9828 19380 9892
rect 19444 9828 19445 9892
rect 19379 9827 19445 9828
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 27294 5541 27354 26827
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 28763 8532 28829 8533
rect 28763 8468 28764 8532
rect 28828 8468 28829 8532
rect 28763 8467 28829 8468
rect 27291 5540 27357 5541
rect 27291 5476 27292 5540
rect 27356 5476 27357 5540
rect 27291 5475 27357 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 28766 4725 28826 8467
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 28763 4724 28829 4725
rect 28763 4660 28764 4724
rect 28828 4660 28829 4724
rect 28763 4659 28829 4660
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 9476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1667941163
transform 1 0 32292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform 1 0 31648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1667941163
transform -1 0 9476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1667941163
transform -1 0 32476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform -1 0 35604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1667941163
transform 1 0 31280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1667941163
transform -1 0 32384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform -1 0 31188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform -1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 9292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform -1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1667941163
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1667941163
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1667941163
transform -1 0 31188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1667941163
transform -1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1667941163
transform -1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1667941163
transform -1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform 1 0 10488 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1667941163
transform -1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform -1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1667941163
transform 1 0 29348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 27876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform -1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform -1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform -1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A
timestamp 1667941163
transform -1 0 27324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform -1 0 34408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform -1 0 34960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1667941163
transform -1 0 25944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1667941163
transform -1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1667941163
transform -1 0 28704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1667941163
transform -1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform 1 0 9108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform -1 0 18860 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform -1 0 15456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform -1 0 20976 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform -1 0 35604 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1667941163
transform -1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform -1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1667941163
transform 1 0 27140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform -1 0 31372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform -1 0 30544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform 1 0 29992 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform 1 0 30820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform 1 0 9844 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform -1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform -1 0 31556 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform -1 0 34868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform -1 0 35052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1667941163
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1667941163
transform -1 0 33028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform -1 0 10580 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform -1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1667941163
transform -1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform 1 0 23000 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1667941163
transform -1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform -1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform 1 0 36340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform -1 0 37628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform 1 0 37076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 36616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A
timestamp 1667941163
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1667941163
transform -1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1667941163
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1667941163
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1667941163
transform 1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1667941163
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1667941163
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1667941163
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1667941163
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1667941163
transform -1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1667941163
transform 1 0 35328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1667941163
transform 1 0 34040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__A
timestamp 1667941163
transform 1 0 34868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__A
timestamp 1667941163
transform 1 0 35880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A
timestamp 1667941163
transform 1 0 35972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__A
timestamp 1667941163
transform 1 0 33488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__A
timestamp 1667941163
transform -1 0 36708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__A
timestamp 1667941163
transform 1 0 35236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__A
timestamp 1667941163
transform 1 0 33580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1667941163
transform 1 0 34132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1667941163
transform 1 0 35788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A
timestamp 1667941163
transform 1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A
timestamp 1667941163
transform 1 0 34132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1667941163
transform 1 0 36432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 32292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__D
timestamp 1667941163
transform 1 0 30912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform -1 0 6716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__RESET_B
timestamp 1667941163
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__RESET_B
timestamp 1667941163
transform -1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 27876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 20792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 31464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__D
timestamp 1667941163
transform -1 0 31648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 34224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 33028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 19136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__RESET_B
timestamp 1667941163
transform -1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__RESET_B
timestamp 1667941163
transform -1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 10212 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1667941163
transform -1 0 9844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__D
timestamp 1667941163
transform 1 0 12420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1667941163
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 12880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 31556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__RESET_B
timestamp 1667941163
transform -1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__RESET_B
timestamp 1667941163
transform -1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__RESET_B
timestamp 1667941163
transform -1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 6624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__D
timestamp 1667941163
transform 1 0 8832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 7912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__D
timestamp 1667941163
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__RESET_B
timestamp 1667941163
transform -1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__D
timestamp 1667941163
transform -1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__RESET_B
timestamp 1667941163
transform -1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 34868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 33580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__D
timestamp 1667941163
transform -1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__CLK
timestamp 1667941163
transform 1 0 30912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__CLK
timestamp 1667941163
transform 1 0 32936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__CLK
timestamp 1667941163
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__CLK
timestamp 1667941163
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__D
timestamp 1667941163
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__D
timestamp 1667941163
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__CLK
timestamp 1667941163
transform 1 0 9568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1667941163
transform -1 0 17848 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform -1 0 33580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1667941163
transform -1 0 34316 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1667941163
transform -1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1667941163
transform -1 0 5796 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform 1 0 14168 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1667941163
transform -1 0 36156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1667941163
transform -1 0 22816 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1667941163
transform -1 0 27968 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1667941163
transform 1 0 25668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1667941163
transform 1 0 2392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1667941163
transform -1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1667941163
transform 1 0 34224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1667941163
transform 1 0 21252 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A
timestamp 1667941163
transform -1 0 4876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1667941163
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1667941163
transform -1 0 10488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1667941163
transform -1 0 30912 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1667941163
transform -1 0 21160 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform -1 0 2576 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1667941163
transform -1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1667941163
transform -1 0 15640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1667941163
transform -1 0 25944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1667941163
transform -1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1667941163
transform 1 0 22632 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 37628 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 38088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 37720 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 37628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 22908 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 36248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 37628 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform 1 0 13616 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 2760 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 1748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 1748 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 37812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 1748 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 35696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 6808 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 34132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 3312 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1667941163
transform -1 0 37628 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1667941163
transform -1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform -1 0 35604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1667941163
transform 1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1667941163
transform -1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48
timestamp 1667941163
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71
timestamp 1667941163
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1667941163
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_259
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1667941163
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1667941163
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_375
timestamp 1667941163
transform 1 0 35604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_380
timestamp 1667941163
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1667941163
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1667941163
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1667941163
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1667941163
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1667941163
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1667941163
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_298
timestamp 1667941163
transform 1 0 28520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_312
timestamp 1667941163
transform 1 0 29808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1667941163
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_326
timestamp 1667941163
transform 1 0 31096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1667941163
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1667941163
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1667941163
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1667941163
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1667941163
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1667941163
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_401
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_36
timestamp 1667941163
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1667941163
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1667941163
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1667941163
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1667941163
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1667941163
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 1667941163
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1667941163
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1667941163
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1667941163
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_94
timestamp 1667941163
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_101
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_107
timestamp 1667941163
transform 1 0 10948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_111
timestamp 1667941163
transform 1 0 11316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1667941163
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1667941163
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1667941163
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1667941163
transform 1 0 27600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1667941163
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1667941163
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1667941163
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_356
timestamp 1667941163
transform 1 0 33856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1667941163
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1667941163
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1667941163
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_381
timestamp 1667941163
transform 1 0 36156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_387
timestamp 1667941163
transform 1 0 36708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_394
timestamp 1667941163
transform 1 0 37352 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_400
timestamp 1667941163
transform 1 0 37904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7
timestamp 1667941163
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_19
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_31
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1667941163
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_38
timestamp 1667941163
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1667941163
transform 1 0 5704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1667941163
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1667941163
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1667941163
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1667941163
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1667941163
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1667941163
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_104
timestamp 1667941163
transform 1 0 10672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1667941163
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_175
timestamp 1667941163
transform 1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1667941163
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1667941163
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_214
timestamp 1667941163
transform 1 0 20792 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_292
timestamp 1667941163
transform 1 0 27968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1667941163
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_324
timestamp 1667941163
transform 1 0 30912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1667941163
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1667941163
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1667941163
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_362
timestamp 1667941163
transform 1 0 34408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1667941163
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_374
timestamp 1667941163
transform 1 0 35512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1667941163
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_397
timestamp 1667941163
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1667941163
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1667941163
transform 1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1667941163
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_76
timestamp 1667941163
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1667941163
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1667941163
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_100
timestamp 1667941163
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1667941163
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1667941163
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1667941163
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1667941163
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1667941163
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_164
timestamp 1667941163
transform 1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_172
timestamp 1667941163
transform 1 0 16928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_220
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_226
timestamp 1667941163
transform 1 0 21896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1667941163
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_259
timestamp 1667941163
transform 1 0 24932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1667941163
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1667941163
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1667941163
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1667941163
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_328
timestamp 1667941163
transform 1 0 31280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_342
timestamp 1667941163
transform 1 0 32568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1667941163
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_355
timestamp 1667941163
transform 1 0 33764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1667941163
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_369
timestamp 1667941163
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_375
timestamp 1667941163
transform 1 0 35604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1667941163
transform 1 0 36156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_387
timestamp 1667941163
transform 1 0 36708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_393
timestamp 1667941163
transform 1 0 37260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_28
timestamp 1667941163
transform 1 0 3680 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_40
timestamp 1667941163
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1667941163
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1667941163
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1667941163
transform 1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1667941163
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1667941163
transform 1 0 8464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1667941163
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1667941163
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1667941163
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1667941163
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1667941163
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1667941163
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp 1667941163
transform 1 0 24380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1667941163
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_263
timestamp 1667941163
transform 1 0 25300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1667941163
transform 1 0 25944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_274
timestamp 1667941163
transform 1 0 26312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_287
timestamp 1667941163
transform 1 0 27508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1667941163
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1667941163
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_308
timestamp 1667941163
transform 1 0 29440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1667941163
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_322
timestamp 1667941163
transform 1 0 30728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_342
timestamp 1667941163
transform 1 0 32568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_355
timestamp 1667941163
transform 1 0 33764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1667941163
transform 1 0 34868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_379
timestamp 1667941163
transform 1 0 35972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_399
timestamp 1667941163
transform 1 0 37812 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1667941163
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1667941163
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_35
timestamp 1667941163
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 1667941163
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_76
timestamp 1667941163
transform 1 0 8096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1667941163
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp 1667941163
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1667941163
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1667941163
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1667941163
transform 1 0 11316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1667941163
transform 1 0 11868 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1667941163
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_167
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1667941163
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_202
timestamp 1667941163
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1667941163
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_216
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_296
timestamp 1667941163
transform 1 0 28336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_314
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp 1667941163
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_335
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_342
timestamp 1667941163
transform 1 0 32568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_349
timestamp 1667941163
transform 1 0 33212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_355
timestamp 1667941163
transform 1 0 33764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1667941163
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_369
timestamp 1667941163
transform 1 0 35052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1667941163
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_379
timestamp 1667941163
transform 1 0 35972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_382
timestamp 1667941163
transform 1 0 36248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_388
timestamp 1667941163
transform 1 0 36800 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_394
timestamp 1667941163
transform 1 0 37352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1667941163
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1667941163
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1667941163
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1667941163
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1667941163
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_90
timestamp 1667941163
transform 1 0 9384 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1667941163
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1667941163
transform 1 0 10672 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_121
timestamp 1667941163
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1667941163
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1667941163
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_158
timestamp 1667941163
transform 1 0 15640 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_162
timestamp 1667941163
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1667941163
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_271
timestamp 1667941163
transform 1 0 26036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_297
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1667941163
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_308
timestamp 1667941163
transform 1 0 29440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_315
timestamp 1667941163
transform 1 0 30084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_322
timestamp 1667941163
transform 1 0 30728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_348
timestamp 1667941163
transform 1 0 33120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_354
timestamp 1667941163
transform 1 0 33672 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_360
timestamp 1667941163
transform 1 0 34224 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_372
timestamp 1667941163
transform 1 0 35328 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1667941163
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_397
timestamp 1667941163
transform 1 0 37628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_89
timestamp 1667941163
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1667941163
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1667941163
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1667941163
transform 1 0 10948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1667941163
transform 1 0 11500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 1667941163
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1667941163
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1667941163
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1667941163
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1667941163
transform 1 0 21252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_223
timestamp 1667941163
transform 1 0 21620 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_278
timestamp 1667941163
transform 1 0 26680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1667941163
transform 1 0 27324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1667941163
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1667941163
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_314
timestamp 1667941163
transform 1 0 29992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1667941163
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_335
timestamp 1667941163
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_341
timestamp 1667941163
transform 1 0 32476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_347
timestamp 1667941163
transform 1 0 33028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1667941163
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1667941163
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1667941163
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_91
timestamp 1667941163
transform 1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_97
timestamp 1667941163
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1667941163
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1667941163
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_173
timestamp 1667941163
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1667941163
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1667941163
transform 1 0 18308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1667941163
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_218
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1667941163
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_262
timestamp 1667941163
transform 1 0 25208 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_268
timestamp 1667941163
transform 1 0 25760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_292
timestamp 1667941163
transform 1 0 27968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_299
timestamp 1667941163
transform 1 0 28612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_306
timestamp 1667941163
transform 1 0 29256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1667941163
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1667941163
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_327
timestamp 1667941163
transform 1 0 31188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1667941163
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_341
timestamp 1667941163
transform 1 0 32476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_353
timestamp 1667941163
transform 1 0 33580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1667941163
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1667941163
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1667941163
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1667941163
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1667941163
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1667941163
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp 1667941163
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1667941163
transform 1 0 11500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_147
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1667941163
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1667941163
transform 1 0 21528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_226
timestamp 1667941163
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_284
timestamp 1667941163
transform 1 0 27232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_297
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 29992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_328
timestamp 1667941163
transform 1 0 31280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1667941163
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_340
timestamp 1667941163
transform 1 0 32384 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_352
timestamp 1667941163
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1667941163
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1667941163
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1667941163
transform 1 0 10120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1667941163
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1667941163
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1667941163
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1667941163
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_250
timestamp 1667941163
transform 1 0 24104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1667941163
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_292
timestamp 1667941163
transform 1 0 27968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1667941163
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1667941163
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1667941163
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_326
timestamp 1667941163
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1667941163
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_341
timestamp 1667941163
transform 1 0 32476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_353
timestamp 1667941163
transform 1 0 33580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_365
timestamp 1667941163
transform 1 0 34684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_377
timestamp 1667941163
transform 1 0 35788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1667941163
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1667941163
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1667941163
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1667941163
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_131
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_164
timestamp 1667941163
transform 1 0 16192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1667941163
transform 1 0 16744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1667941163
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_215
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_244
timestamp 1667941163
transform 1 0 23552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1667941163
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_257
timestamp 1667941163
transform 1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1667941163
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_281
timestamp 1667941163
transform 1 0 26956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_293
timestamp 1667941163
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1667941163
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_320
timestamp 1667941163
transform 1 0 30544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_326
timestamp 1667941163
transform 1 0 31096 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_332
timestamp 1667941163
transform 1 0 31648 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_344
timestamp 1667941163
transform 1 0 32752 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_356
timestamp 1667941163
transform 1 0 33856 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1667941163
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_90
timestamp 1667941163
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1667941163
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_122
timestamp 1667941163
transform 1 0 12328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1667941163
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_160
timestamp 1667941163
transform 1 0 15824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1667941163
transform 1 0 18032 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1667941163
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_248
timestamp 1667941163
transform 1 0 23920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_252
timestamp 1667941163
transform 1 0 24288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_262
timestamp 1667941163
transform 1 0 25208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1667941163
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1667941163
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1667941163
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1667941163
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_321
timestamp 1667941163
transform 1 0 30636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 1667941163
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_92
timestamp 1667941163
transform 1 0 9568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1667941163
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1667941163
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1667941163
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1667941163
transform 1 0 12788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1667941163
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1667941163
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_202
timestamp 1667941163
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_208
timestamp 1667941163
transform 1 0 20240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_222
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_235
timestamp 1667941163
transform 1 0 22724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_268
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_275
timestamp 1667941163
transform 1 0 26404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_279
timestamp 1667941163
transform 1 0 26772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1667941163
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_327
timestamp 1667941163
transform 1 0 31188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_339
timestamp 1667941163
transform 1 0 32292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_351
timestamp 1667941163
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1667941163
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1667941163
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1667941163
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1667941163
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1667941163
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1667941163
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1667941163
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1667941163
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1667941163
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1667941163
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1667941163
transform 1 0 23184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1667941163
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_256
timestamp 1667941163
transform 1 0 24656 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_265
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_269
timestamp 1667941163
transform 1 0 25852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1667941163
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_296
timestamp 1667941163
transform 1 0 28336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1667941163
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_324
timestamp 1667941163
transform 1 0 30912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1667941163
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_402
timestamp 1667941163
transform 1 0 38088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_406
timestamp 1667941163
transform 1 0 38456 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_91
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_98
timestamp 1667941163
transform 1 0 10120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1667941163
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1667941163
transform 1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1667941163
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1667941163
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1667941163
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1667941163
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_231
timestamp 1667941163
transform 1 0 22356 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 1667941163
transform 1 0 23460 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_263
timestamp 1667941163
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1667941163
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_284
timestamp 1667941163
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1667941163
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_327
timestamp 1667941163
transform 1 0 31188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_339
timestamp 1667941163
transform 1 0 32292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_351
timestamp 1667941163
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1667941163
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1667941163
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_92
timestamp 1667941163
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1667941163
transform 1 0 15364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1667941163
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1667941163
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_229
timestamp 1667941163
transform 1 0 22172 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1667941163
transform 1 0 24840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_262
timestamp 1667941163
transform 1 0 25208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 1667941163
transform 1 0 26036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1667941163
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1667941163
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_313
timestamp 1667941163
transform 1 0 29900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1667941163
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1667941163
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_401
timestamp 1667941163
transform 1 0 37996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_71
timestamp 1667941163
transform 1 0 7636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_89
timestamp 1667941163
transform 1 0 9292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1667941163
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_116
timestamp 1667941163
transform 1 0 11776 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_129
timestamp 1667941163
transform 1 0 12972 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1667941163
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1667941163
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1667941163
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1667941163
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_231
timestamp 1667941163
transform 1 0 22356 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_276
timestamp 1667941163
transform 1 0 26496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_283
timestamp 1667941163
transform 1 0 27140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1667941163
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1667941163
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1667941163
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_320
timestamp 1667941163
transform 1 0 30544 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_332
timestamp 1667941163
transform 1 0 31648 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_344
timestamp 1667941163
transform 1 0 32752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_356
timestamp 1667941163
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1667941163
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1667941163
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_80
timestamp 1667941163
transform 1 0 8464 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1667941163
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1667941163
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1667941163
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1667941163
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1667941163
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_151
timestamp 1667941163
transform 1 0 14996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_180
timestamp 1667941163
transform 1 0 17664 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_195
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1667941163
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1667941163
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_267
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1667941163
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp 1667941163
transform 1 0 28612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_303
timestamp 1667941163
transform 1 0 28980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_313
timestamp 1667941163
transform 1 0 29900 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_316
timestamp 1667941163
transform 1 0 30176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1667941163
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_10
timestamp 1667941163
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_16
timestamp 1667941163
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_91
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1667941163
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1667941163
transform 1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_124
timestamp 1667941163
transform 1 0 12512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1667941163
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1667941163
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1667941163
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_178
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_184
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1667941163
transform 1 0 20424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1667941163
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_287
timestamp 1667941163
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1667941163
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_101
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_104
timestamp 1667941163
transform 1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1667941163
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_187
timestamp 1667941163
transform 1 0 18308 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_203
timestamp 1667941163
transform 1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_209
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_244
timestamp 1667941163
transform 1 0 23552 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_264
timestamp 1667941163
transform 1 0 25392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1667941163
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_285
timestamp 1667941163
transform 1 0 27324 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_291
timestamp 1667941163
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_303
timestamp 1667941163
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_315
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_327
timestamp 1667941163
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_401
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_7
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1667941163
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_104
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_152
timestamp 1667941163
transform 1 0 15088 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_169
timestamp 1667941163
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1667941163
transform 1 0 17020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_183
timestamp 1667941163
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1667941163
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1667941163
transform 1 0 20240 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_272
timestamp 1667941163
transform 1 0 26128 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_285
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1667941163
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1667941163
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_16
timestamp 1667941163
transform 1 0 2576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_28
timestamp 1667941163
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1667941163
transform 1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 1667941163
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1667941163
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_97
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1667941163
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_122
timestamp 1667941163
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1667941163
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1667941163
transform 1 0 19504 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1667941163
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1667941163
transform 1 0 10856 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_112
timestamp 1667941163
transform 1 0 11408 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_169
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1667941163
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1667941163
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_275
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_287
timestamp 1667941163
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1667941163
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_325
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_329
timestamp 1667941163
transform 1 0 31372 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_341
timestamp 1667941163
transform 1 0 32476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_353
timestamp 1667941163
transform 1 0 33580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1667941163
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1667941163
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_134
timestamp 1667941163
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1667941163
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1667941163
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1667941163
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1667941163
transform 1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1667941163
transform 1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1667941163
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1667941163
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_257
timestamp 1667941163
transform 1 0 24748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_264
timestamp 1667941163
transform 1 0 25392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1667941163
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_348
timestamp 1667941163
transform 1 0 33120 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_360
timestamp 1667941163
transform 1 0 34224 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_372
timestamp 1667941163
transform 1 0 35328 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_161
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1667941163
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_202
timestamp 1667941163
transform 1 0 19688 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_214
timestamp 1667941163
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_222
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1667941163
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_264
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_276
timestamp 1667941163
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_288
timestamp 1667941163
transform 1 0 27600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1667941163
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1667941163
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 1667941163
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_182
timestamp 1667941163
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1667941163
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1667941163
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_263
timestamp 1667941163
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1667941163
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_207
timestamp 1667941163
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_224
timestamp 1667941163
transform 1 0 21712 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_239
timestamp 1667941163
transform 1 0 23092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1667941163
transform 1 0 25300 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_269
timestamp 1667941163
transform 1 0 25852 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_281
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1667941163
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1667941163
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1667941163
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_274
timestamp 1667941163
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1667941163
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1667941163
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1667941163
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_349
timestamp 1667941163
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1667941163
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_285
timestamp 1667941163
transform 1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_293
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1667941163
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_395
timestamp 1667941163
transform 1 0 37444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_398
timestamp 1667941163
transform 1 0 37720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_7
timestamp 1667941163
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1667941163
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_397
timestamp 1667941163
transform 1 0 37628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_402
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1667941163
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_74
timestamp 1667941163
transform 1 0 7912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1667941163
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_399
timestamp 1667941163
transform 1 0 37812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1667941163
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1667941163
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_402
timestamp 1667941163
transform 1 0 38088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1667941163
transform 1 0 38456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_10
timestamp 1667941163
transform 1 0 2024 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_16
timestamp 1667941163
transform 1 0 2576 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1667941163
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_269
timestamp 1667941163
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_281
timestamp 1667941163
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_293
timestamp 1667941163
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1667941163
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1667941163
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1667941163
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_211
timestamp 1667941163
transform 1 0 20516 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_215
timestamp 1667941163
transform 1 0 20884 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_397
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1667941163
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_356
timestamp 1667941163
transform 1 0 33856 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_362
timestamp 1667941163
transform 1 0 34408 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_374
timestamp 1667941163
transform 1 0 35512 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1667941163
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_401
timestamp 1667941163
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_404
timestamp 1667941163
transform 1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1667941163
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_152
timestamp 1667941163
transform 1 0 15088 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_176
timestamp 1667941163
transform 1 0 17296 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1667941163
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1667941163
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_205
timestamp 1667941163
transform 1 0 19964 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_211
timestamp 1667941163
transform 1 0 20516 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_223
timestamp 1667941163
transform 1 0 21620 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_235
timestamp 1667941163
transform 1 0 22724 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1667941163
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_397
timestamp 1667941163
transform 1 0 37628 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_402
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1667941163
transform 1 0 38456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1667941163
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_153
timestamp 1667941163
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_156
timestamp 1667941163
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_187
timestamp 1667941163
transform 1 0 18308 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_229
timestamp 1667941163
transform 1 0 22172 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1667941163
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_21
timestamp 1667941163
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_33
timestamp 1667941163
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1667941163
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1667941163
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_323
timestamp 1667941163
transform 1 0 30820 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_212
timestamp 1667941163
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1667941163
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_321
timestamp 1667941163
transform 1 0 30636 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1667941163
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1667941163
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1667941163
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_197
timestamp 1667941163
transform 1 0 19228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_201
timestamp 1667941163
transform 1 0 19596 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1667941163
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1667941163
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_324
timestamp 1667941163
transform 1 0 30912 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_336
timestamp 1667941163
transform 1 0 32016 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_348
timestamp 1667941163
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1667941163
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_7
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_19
timestamp 1667941163
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_31
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_43
timestamp 1667941163
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1667941163
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_93
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_103
timestamp 1667941163
transform 1 0 10580 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_115
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_127
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1667941163
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_236
timestamp 1667941163
transform 1 0 22816 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_248
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_260
timestamp 1667941163
transform 1 0 25024 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1667941163
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_7
timestamp 1667941163
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1667941163
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_45
timestamp 1667941163
transform 1 0 5244 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_51
timestamp 1667941163
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_63
timestamp 1667941163
transform 1 0 6900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_75
timestamp 1667941163
transform 1 0 8004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_96
timestamp 1667941163
transform 1 0 9936 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_102
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_114
timestamp 1667941163
transform 1 0 11592 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_126
timestamp 1667941163
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1667941163
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1667941163
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_182
timestamp 1667941163
transform 1 0 17848 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_397
timestamp 1667941163
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_18
timestamp 1667941163
transform 1 0 2760 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_24
timestamp 1667941163
transform 1 0 3312 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_36
timestamp 1667941163
transform 1 0 4416 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1667941163
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_133
timestamp 1667941163
transform 1 0 13340 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1667941163
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_155
timestamp 1667941163
transform 1 0 15364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_213
timestamp 1667941163
transform 1 0 20700 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1667941163
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1667941163
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1667941163
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_248
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1667941163
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1667941163
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_292
timestamp 1667941163
transform 1 0 27968 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_304
timestamp 1667941163
transform 1 0 29072 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_316
timestamp 1667941163
transform 1 0 30176 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1667941163
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_397
timestamp 1667941163
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_14
timestamp 1667941163
transform 1 0 2392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1667941163
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_91
timestamp 1667941163
transform 1 0 9476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_99
timestamp 1667941163
transform 1 0 10212 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_134
timestamp 1667941163
transform 1 0 13432 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1667941163
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_211
timestamp 1667941163
transform 1 0 20516 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_378
timestamp 1667941163
transform 1 0 35880 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _216_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform 1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform -1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform 1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform -1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 29808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 29624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 29992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform 1 0 26404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 30360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 30360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform 1 0 29808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform -1 0 30912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 28796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 11224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform 1 0 20976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform -1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform 1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 26404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 25944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 18400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 12328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform 1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 21344 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform -1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform -1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 12328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform 1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform 1 0 24748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform 1 0 22448 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 27140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 14720 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform -1 0 26588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform -1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform 1 0 29624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 28980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform -1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform -1 0 29072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform 1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform -1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform -1 0 23920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform -1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform 1 0 28704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform -1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform 1 0 27508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform -1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform -1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform -1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform -1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 13524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform -1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform -1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform -1 0 13156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform -1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform -1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform -1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform -1 0 18308 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform 1 0 10580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform -1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform 1 0 37812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 21528 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform -1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform 1 0 10212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform -1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform 1 0 30544 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 29348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform -1 0 29992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform -1 0 28704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform 1 0 13156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform -1 0 31004 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform -1 0 28980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform -1 0 10028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform -1 0 27232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1667941163
transform -1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform -1 0 30452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform -1 0 28060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform -1 0 25760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform 1 0 7636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform -1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 19596 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform -1 0 33120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform -1 0 33212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform -1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform -1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1667941163
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform -1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform 1 0 31096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _398_
timestamp 1667941163
transform -1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform -1 0 28980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform -1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform -1 0 28796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform -1 0 30544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1667941163
transform -1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform -1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform -1 0 32568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform -1 0 30084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _409_
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform -1 0 31280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 30728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform -1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1667941163
transform -1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform -1 0 29992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _420_
timestamp 1667941163
transform -1 0 37352 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform -1 0 33212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform -1 0 31924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform -1 0 31280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1667941163
transform -1 0 29624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform -1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 31280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform -1 0 29992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 30728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform -1 0 31280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _431_
timestamp 1667941163
transform -1 0 36984 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform -1 0 30544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform -1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1667941163
transform -1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform -1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform -1 0 31924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _442_
timestamp 1667941163
transform -1 0 7636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1667941163
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 3496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _453_
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform -1 0 33212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform -1 0 30912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 31096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1667941163
transform -1 0 24748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1667941163
transform -1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1667941163
transform -1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1667941163
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1667941163
transform -1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1667941163
transform -1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _475_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24104 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform -1 0 18860 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _479_
timestamp 1667941163
transform 1 0 14076 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1667941163
transform 1 0 11868 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _481_
timestamp 1667941163
transform -1 0 21528 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform 1 0 19228 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform -1 0 21528 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _485_
timestamp 1667941163
transform 1 0 20976 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1667941163
transform 1 0 24472 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _487_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform 1 0 19688 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _491_
timestamp 1667941163
transform -1 0 21528 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _492_
timestamp 1667941163
transform -1 0 23644 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _493_
timestamp 1667941163
transform 1 0 22080 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform -1 0 13708 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform -1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _497_
timestamp 1667941163
transform 1 0 18676 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _498_
timestamp 1667941163
transform 1 0 15640 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _499_
timestamp 1667941163
transform -1 0 23644 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform -1 0 20608 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _503_
timestamp 1667941163
transform -1 0 23920 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _505_
timestamp 1667941163
transform 1 0 17296 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform -1 0 18952 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _509_
timestamp 1667941163
transform -1 0 15824 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _510_
timestamp 1667941163
transform -1 0 14076 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _511_
timestamp 1667941163
transform -1 0 16376 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform -1 0 14168 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _515_
timestamp 1667941163
transform -1 0 15640 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _516_
timestamp 1667941163
transform -1 0 16192 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1667941163
transform -1 0 16376 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform -1 0 14168 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _521_
timestamp 1667941163
transform -1 0 15824 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _522_
timestamp 1667941163
transform 1 0 14536 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1667941163
transform 1 0 14352 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 26036 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform 1 0 22080 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _527_
timestamp 1667941163
transform 1 0 21988 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _528_
timestamp 1667941163
transform 1 0 17572 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _529_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _530_
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _531_
timestamp 1667941163
transform 1 0 24196 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 1667941163
transform 1 0 19504 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _533_
timestamp 1667941163
transform 1 0 17020 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _534_
timestamp 1667941163
transform 1 0 17204 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _535_
timestamp 1667941163
transform -1 0 22632 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _547_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18492 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1667941163
transform -1 0 34224 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1667941163
transform -1 0 21344 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1667941163
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1667941163
transform -1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform -1 0 5244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1667941163
transform -1 0 38088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1667941163
transform -1 0 28520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform -1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1667941163
transform 1 0 37812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1667941163
transform -1 0 22264 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1667941163
transform -1 0 27416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _563_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24104 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1667941163
transform 1 0 7636 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _566_
timestamp 1667941163
transform 1 0 33580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform 1 0 20608 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform -1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform 1 0 4048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1667941163
transform 1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 9660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1667941163
transform -1 0 30360 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform -1 0 20608 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform -1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _576_
timestamp 1667941163
transform -1 0 27508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _578_
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _579_
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _580_
timestamp 1667941163
transform 1 0 23736 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _581_
timestamp 1667941163
transform -1 0 25300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _582_
timestamp 1667941163
transform 1 0 24472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _583_
timestamp 1667941163
transform -1 0 38088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _586_
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _587_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16008 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _589__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _590_
timestamp 1667941163
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _592_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _593_
timestamp 1667941163
transform -1 0 22724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _596_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _597_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _598_
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _600_
timestamp 1667941163
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _601_
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _601__92
timestamp 1667941163
transform -1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _602_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _603_
timestamp 1667941163
transform -1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _604_
timestamp 1667941163
transform 1 0 20424 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _605_
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _606_
timestamp 1667941163
transform 1 0 12144 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform -1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _608_
timestamp 1667941163
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _609_
timestamp 1667941163
transform 1 0 26312 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _610_
timestamp 1667941163
transform 1 0 22908 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform 1 0 20516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _612_
timestamp 1667941163
transform -1 0 24380 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _612__93
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _613_
timestamp 1667941163
transform -1 0 26496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _614_
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _615_
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _616_
timestamp 1667941163
transform -1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _617_
timestamp 1667941163
transform -1 0 24840 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _618_
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _619_
timestamp 1667941163
transform -1 0 26496 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _620_
timestamp 1667941163
transform -1 0 24196 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _621_
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _622_
timestamp 1667941163
transform -1 0 27232 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _623_
timestamp 1667941163
transform -1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _624__94
timestamp 1667941163
transform 1 0 29716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _624_
timestamp 1667941163
transform -1 0 25852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _625_
timestamp 1667941163
transform -1 0 26680 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform -1 0 26680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _627_
timestamp 1667941163
transform -1 0 25484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _628_
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _629_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _630_
timestamp 1667941163
transform -1 0 29164 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform -1 0 27968 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _632_
timestamp 1667941163
transform -1 0 24288 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _633_
timestamp 1667941163
transform -1 0 21528 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _634_
timestamp 1667941163
transform 1 0 15364 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636__95
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform -1 0 27968 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _639_
timestamp 1667941163
transform -1 0 26312 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform -1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _641_
timestamp 1667941163
transform 1 0 17756 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform -1 0 18952 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _643_
timestamp 1667941163
transform -1 0 25392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform -1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform -1 0 25392 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform -1 0 18860 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _647_
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _648__96
timestamp 1667941163
transform -1 0 18584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _648_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _649_
timestamp 1667941163
transform -1 0 25116 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _650_
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _651_
timestamp 1667941163
transform -1 0 25300 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _652_
timestamp 1667941163
transform 1 0 22356 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform -1 0 24104 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _654_
timestamp 1667941163
transform -1 0 19688 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _655_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _656_
timestamp 1667941163
transform -1 0 23828 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 19504 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform 1 0 18216 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform 1 0 12696 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _660__97
timestamp 1667941163
transform -1 0 13156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _661_
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform -1 0 22540 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _667_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _668_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _669_
timestamp 1667941163
transform -1 0 12420 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform -1 0 11224 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform -1 0 13524 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _672__98
timestamp 1667941163
transform -1 0 10672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 11040 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform 1 0 11776 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform -1 0 17204 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _675_
timestamp 1667941163
transform -1 0 20240 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _676_
timestamp 1667941163
transform -1 0 17480 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform -1 0 13616 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform 1 0 11868 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform 1 0 15824 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _680_
timestamp 1667941163
transform -1 0 19780 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform -1 0 16008 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform -1 0 15916 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _683_
timestamp 1667941163
transform -1 0 20332 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _684__99
timestamp 1667941163
transform -1 0 11224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform -1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform -1 0 24104 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform -1 0 13800 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform 1 0 17020 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 21804 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 29716 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform 1 0 28520 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _695_
timestamp 1667941163
transform 1 0 27324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _696__100
timestamp 1667941163
transform 1 0 30360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _696_
timestamp 1667941163
transform -1 0 28796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform -1 0 27968 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform 1 0 28244 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _699_
timestamp 1667941163
transform -1 0 26680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _700_
timestamp 1667941163
transform -1 0 28336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _702_
timestamp 1667941163
transform -1 0 26680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 26864 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _704_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _705_
timestamp 1667941163
transform -1 0 27600 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _706_
timestamp 1667941163
transform -1 0 23184 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _708_
timestamp 1667941163
transform 1 0 21896 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _708__101
timestamp 1667941163
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _709_
timestamp 1667941163
transform -1 0 27876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _710_
timestamp 1667941163
transform -1 0 25760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _711_
timestamp 1667941163
transform -1 0 25208 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _712_
timestamp 1667941163
transform -1 0 28428 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _713_
timestamp 1667941163
transform 1 0 19412 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _714_
timestamp 1667941163
transform -1 0 21528 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _715_
timestamp 1667941163
transform -1 0 26036 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _716_
timestamp 1667941163
transform 1 0 19504 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform -1 0 38364 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 38088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform -1 0 35880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform -1 0 38364 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 20608 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform 1 0 2024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 13800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform -1 0 38364 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 2760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform -1 0 38364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform -1 0 38364 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1667941163
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform -1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform -1 0 38364 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1667941163
transform -1 0 38364 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform -1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform -1 0 15916 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform -1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 10764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 24104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform -1 0 12696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 36984 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 30820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform -1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 9476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 78 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 79 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 80 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 pReset
port 81 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 prog_clk
port 82 nsew signal input
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
port 83 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_
port 86 nsew signal tristate
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_
port 87 nsew signal tristate
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_
port 88 nsew signal tristate
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_
port 89 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_
port 90 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 vssd1
port 92 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 28106 3978 28106 3978 0 _000_
rlabel metal1 30452 6086 30452 6086 0 _001_
rlabel metal1 19143 6698 19143 6698 0 _002_
rlabel metal1 16153 8874 16153 8874 0 _003_
rlabel metal1 18913 8874 18913 8874 0 _004_
rlabel metal1 27876 5338 27876 5338 0 _005_
rlabel metal2 19366 5287 19366 5287 0 _006_
rlabel metal2 17894 5729 17894 5729 0 _007_
rlabel metal2 5474 2108 5474 2108 0 _008_
rlabel metal2 16514 6936 16514 6936 0 _009_
rlabel metal1 13945 7786 13945 7786 0 _010_
rlabel metal1 20799 7786 20799 7786 0 _011_
rlabel metal1 30774 5202 30774 5202 0 _012_
rlabel via2 32430 4539 32430 4539 0 _013_
rlabel metal2 31786 6052 31786 6052 0 _014_
rlabel metal1 30406 5882 30406 5882 0 _015_
rlabel metal1 29670 4794 29670 4794 0 _016_
rlabel metal3 26220 1972 26220 1972 0 _017_
rlabel metal3 30268 2652 30268 2652 0 _018_
rlabel metal3 28474 2516 28474 2516 0 _019_
rlabel metal3 27692 2244 27692 2244 0 _020_
rlabel metal2 20654 7701 20654 7701 0 _021_
rlabel metal2 22862 7310 22862 7310 0 _022_
rlabel metal2 30406 5440 30406 5440 0 _023_
rlabel metal1 12282 7337 12282 7337 0 _024_
rlabel via2 15134 9979 15134 9979 0 _025_
rlabel metal1 16567 6698 16567 6698 0 _026_
rlabel metal2 21942 7888 21942 7888 0 _027_
rlabel metal1 17395 7786 17395 7786 0 _028_
rlabel metal1 23697 5610 23697 5610 0 _029_
rlabel metal1 21114 9588 21114 9588 0 _030_
rlabel metal1 21489 6766 21489 6766 0 _031_
rlabel metal1 18959 9962 18959 9962 0 _032_
rlabel metal1 23552 9690 23552 9690 0 _033_
rlabel metal2 27922 6800 27922 6800 0 _034_
rlabel metal2 19458 8772 19458 8772 0 _035_
rlabel metal2 17894 2091 17894 2091 0 _036_
rlabel metal1 16107 3094 16107 3094 0 _037_
rlabel metal1 13577 5610 13577 5610 0 _038_
rlabel metal2 14766 8449 14766 8449 0 _039_
rlabel metal1 6440 6426 6440 6426 0 _040_
rlabel metal2 13662 7684 13662 7684 0 _041_
rlabel metal2 10994 3332 10994 3332 0 _042_
rlabel metal2 12558 3196 12558 3196 0 _043_
rlabel metal1 9890 2482 9890 2482 0 _044_
rlabel metal1 6302 5814 6302 5814 0 _045_
rlabel metal1 4416 5882 4416 5882 0 _046_
rlabel metal1 19189 3434 19189 3434 0 _047_
rlabel metal2 9798 5729 9798 5729 0 _048_
rlabel metal2 12466 5406 12466 5406 0 _049_
rlabel metal2 19182 3927 19182 3927 0 _050_
rlabel via2 15042 5253 15042 5253 0 _051_
rlabel metal1 16245 5610 16245 5610 0 _052_
rlabel metal1 16061 3434 16061 3434 0 _053_
rlabel metal1 27278 3128 27278 3128 0 _054_
rlabel metal2 30958 3332 30958 3332 0 _055_
rlabel metal1 23506 2489 23506 2489 0 _056_
rlabel metal1 24847 4522 24847 4522 0 _057_
rlabel metal2 18998 3519 18998 3519 0 _058_
rlabel metal1 21121 4522 21121 4522 0 _059_
rlabel metal1 24288 5338 24288 5338 0 _060_
rlabel metal1 30498 5066 30498 5066 0 _061_
rlabel metal1 21673 2346 21673 2346 0 _062_
rlabel metal1 18446 4699 18446 4699 0 _063_
rlabel metal2 19826 4930 19826 4930 0 _064_
rlabel metal2 21850 3570 21850 3570 0 _065_
rlabel metal1 16238 2958 16238 2958 0 _066_
rlabel metal1 28888 4114 28888 4114 0 _067_
rlabel metal1 35374 3026 35374 3026 0 _068_
rlabel metal1 33166 3468 33166 3468 0 _069_
rlabel metal1 28014 6324 28014 6324 0 _070_
rlabel metal2 9154 6494 9154 6494 0 _071_
rlabel metal1 8326 2312 8326 2312 0 _072_
rlabel metal1 18584 15674 18584 15674 0 _073_
rlabel metal1 20378 15130 20378 15130 0 _074_
rlabel metal1 16422 16490 16422 16490 0 _075_
rlabel metal1 18400 14586 18400 14586 0 _076_
rlabel metal1 17158 15062 17158 15062 0 _077_
rlabel metal1 14076 13974 14076 13974 0 _078_
rlabel metal1 21482 14280 21482 14280 0 _079_
rlabel metal1 24334 7514 24334 7514 0 _080_
rlabel metal2 24702 14926 24702 14926 0 _081_
rlabel metal1 13708 13430 13708 13430 0 _082_
rlabel metal1 15686 15130 15686 15130 0 _083_
rlabel metal1 21850 13226 21850 13226 0 _084_
rlabel metal1 16100 8058 16100 8058 0 _085_
rlabel metal2 14030 13838 14030 13838 0 _086_
rlabel metal1 15686 10710 15686 10710 0 _087_
rlabel metal2 13478 9894 13478 9894 0 _088_
rlabel metal1 10856 9622 10856 9622 0 _089_
rlabel metal1 14122 9146 14122 9146 0 _090_
rlabel metal1 20562 11322 20562 11322 0 _091_
rlabel metal1 20286 13498 20286 13498 0 _092_
rlabel metal1 22540 11798 22540 11798 0 _093_
rlabel metal1 11500 11322 11500 11322 0 _094_
rlabel metal1 16744 12886 16744 12886 0 _095_
rlabel metal1 20424 12342 20424 12342 0 _096_
rlabel metal1 26956 13226 26956 13226 0 _097_
rlabel metal1 23782 13158 23782 13158 0 _098_
rlabel metal1 20608 12410 20608 12410 0 _099_
rlabel metal1 24058 11322 24058 11322 0 _100_
rlabel metal1 26910 12682 26910 12682 0 _101_
rlabel metal2 25530 11900 25530 11900 0 _102_
rlabel metal1 23184 12750 23184 12750 0 _103_
rlabel metal1 25530 12818 25530 12818 0 _104_
rlabel metal1 24840 13974 24840 13974 0 _105_
rlabel metal2 23046 13906 23046 13906 0 _106_
rlabel metal1 27232 13498 27232 13498 0 _107_
rlabel metal2 23966 12308 23966 12308 0 _108_
rlabel metal1 28244 5882 28244 5882 0 _109_
rlabel metal2 29762 8024 29762 8024 0 _110_
rlabel metal1 26956 6766 26956 6766 0 _111_
rlabel metal1 27278 8058 27278 8058 0 _112_
rlabel metal1 26450 7480 26450 7480 0 _113_
rlabel metal1 27002 5882 27002 5882 0 _114_
rlabel metal2 25346 8670 25346 8670 0 _115_
rlabel metal1 22954 11084 22954 11084 0 _116_
rlabel metal2 30130 10302 30130 10302 0 _117_
rlabel metal1 29026 7514 29026 7514 0 _118_
rlabel metal1 28060 9622 28060 9622 0 _119_
rlabel metal1 24380 8058 24380 8058 0 _120_
rlabel metal2 19458 10387 19458 10387 0 _121_
rlabel metal1 13846 9384 13846 9384 0 _122_
rlabel metal1 15318 12410 15318 12410 0 _123_
rlabel metal2 13662 16082 13662 16082 0 _124_
rlabel metal1 28934 4182 28934 4182 0 _125_
rlabel metal2 27002 3672 27002 3672 0 _126_
rlabel metal1 27738 12954 27738 12954 0 _127_
rlabel metal1 26082 12138 26082 12138 0 _128_
rlabel metal2 14490 8160 14490 8160 0 _129_
rlabel metal1 18262 13158 18262 13158 0 _130_
rlabel metal1 26220 12954 26220 12954 0 _131_
rlabel metal2 18814 13566 18814 13566 0 _132_
rlabel metal2 27278 14059 27278 14059 0 _133_
rlabel metal1 18400 14042 18400 14042 0 _134_
rlabel metal1 20792 15674 20792 15674 0 _135_
rlabel metal1 19504 16762 19504 16762 0 _136_
rlabel metal1 25070 16218 25070 16218 0 _137_
rlabel metal1 22954 16218 22954 16218 0 _138_
rlabel metal1 24978 15130 24978 15130 0 _139_
rlabel metal2 23230 16830 23230 16830 0 _140_
rlabel metal1 25254 17102 25254 17102 0 _141_
rlabel metal2 19366 16626 19366 16626 0 _142_
rlabel metal1 24702 16218 24702 16218 0 _143_
rlabel metal2 22770 15198 22770 15198 0 _144_
rlabel metal1 19458 5882 19458 5882 0 _145_
rlabel metal2 13018 10336 13018 10336 0 _146_
rlabel metal1 11224 9146 11224 9146 0 _147_
rlabel metal2 14490 14178 14490 14178 0 _148_
rlabel metal2 18262 15470 18262 15470 0 _149_
rlabel metal2 14674 15912 14674 15912 0 _150_
rlabel metal1 21666 15674 21666 15674 0 _151_
rlabel metal2 19642 15640 19642 15640 0 _152_
rlabel metal1 16652 10166 16652 10166 0 _153_
rlabel metal2 16054 16184 16054 16184 0 _154_
rlabel metal1 16330 14042 16330 14042 0 _155_
rlabel via1 22218 16405 22218 16405 0 _156_
rlabel metal1 11776 8058 11776 8058 0 _157_
rlabel metal2 11086 8738 11086 8738 0 _158_
rlabel metal2 11086 13736 11086 13736 0 _159_
rlabel metal2 11270 14552 11270 14552 0 _160_
rlabel metal1 10810 10710 10810 10710 0 _161_
rlabel metal2 14674 11662 14674 11662 0 _162_
rlabel metal2 20010 15198 20010 15198 0 _163_
rlabel metal2 17250 13583 17250 13583 0 _164_
rlabel metal2 9982 11560 9982 11560 0 _165_
rlabel metal1 11270 12886 11270 12886 0 _166_
rlabel metal1 13984 13498 13984 13498 0 _167_
rlabel metal1 19458 13974 19458 13974 0 _168_
rlabel metal1 16008 6426 16008 6426 0 _169_
rlabel metal1 15548 12886 15548 12886 0 _170_
rlabel metal1 19458 9962 19458 9962 0 _171_
rlabel metal1 14214 11832 14214 11832 0 _172_
rlabel metal1 25622 11322 25622 11322 0 _173_
rlabel metal1 23874 9928 23874 9928 0 _174_
rlabel metal1 17158 12138 17158 12138 0 _175_
rlabel metal2 12926 9928 12926 9928 0 _176_
rlabel metal1 13110 11016 13110 11016 0 _177_
rlabel metal2 15134 14008 15134 14008 0 _178_
rlabel metal2 16606 8772 16606 8772 0 _179_
rlabel metal1 21344 10778 21344 10778 0 _180_
rlabel metal2 29946 7106 29946 7106 0 _181_
rlabel metal1 27232 4998 27232 4998 0 _182_
rlabel metal2 27554 9248 27554 9248 0 _183_
rlabel metal2 28566 10540 28566 10540 0 _184_
rlabel metal1 28474 5814 28474 5814 0 _185_
rlabel metal1 28566 5338 28566 5338 0 _186_
rlabel metal1 28152 10234 28152 10234 0 _187_
rlabel metal2 28106 10948 28106 10948 0 _188_
rlabel metal1 26956 5814 26956 5814 0 _189_
rlabel metal1 29762 8058 29762 8058 0 _190_
rlabel metal2 27094 10234 27094 10234 0 _191_
rlabel metal1 26910 10608 26910 10608 0 _192_
rlabel metal2 27370 4114 27370 4114 0 _193_
rlabel metal1 25116 8058 25116 8058 0 _194_
rlabel metal1 13708 9078 13708 9078 0 _195_
rlabel metal1 20010 7276 20010 7276 0 _196_
rlabel metal1 27646 2924 27646 2924 0 _197_
rlabel metal1 26036 2482 26036 2482 0 _198_
rlabel metal1 26864 8602 26864 8602 0 _199_
rlabel metal1 28428 7514 28428 7514 0 _200_
rlabel metal1 18630 7514 18630 7514 0 _201_
rlabel metal2 21114 10642 21114 10642 0 _202_
rlabel metal2 31234 2108 31234 2108 0 _203_
rlabel metal2 19734 9010 19734 9010 0 _204_
rlabel metal2 38318 26741 38318 26741 0 ccff_head
rlabel metal2 38226 36907 38226 36907 0 ccff_tail
rlabel metal1 38456 36822 38456 36822 0 chany_bottom_in[0]
rlabel metal1 38180 4590 38180 4590 0 chany_bottom_in[10]
rlabel via2 38318 19805 38318 19805 0 chany_bottom_in[11]
rlabel metal1 35282 37434 35282 37434 0 chany_bottom_in[12]
rlabel via2 1702 3485 1702 3485 0 chany_bottom_in[13]
rlabel metal2 1610 19023 1610 19023 0 chany_bottom_in[14]
rlabel metal1 32568 2414 32568 2414 0 chany_bottom_in[15]
rlabel metal3 38786 12308 38786 12308 0 chany_bottom_in[16]
rlabel metal2 20654 38260 20654 38260 0 chany_bottom_in[17]
rlabel metal1 2070 37230 2070 37230 0 chany_bottom_in[18]
rlabel metal1 36018 2414 36018 2414 0 chany_bottom_in[1]
rlabel metal2 14858 823 14858 823 0 chany_bottom_in[2]
rlabel via2 1610 4811 1610 4811 0 chany_bottom_in[3]
rlabel metal2 38226 33439 38226 33439 0 chany_bottom_in[4]
rlabel metal1 13616 37434 13616 37434 0 chany_bottom_in[5]
rlabel metal2 2898 38029 2898 38029 0 chany_bottom_in[6]
rlabel metal2 1702 33439 1702 33439 0 chany_bottom_in[7]
rlabel metal2 38226 5559 38226 5559 0 chany_bottom_in[8]
rlabel metal2 3450 2176 3450 2176 0 chany_bottom_in[9]
rlabel metal2 38226 28815 38226 28815 0 chany_bottom_out[0]
rlabel metal1 16882 37094 16882 37094 0 chany_bottom_out[10]
rlabel metal2 38226 32113 38226 32113 0 chany_bottom_out[11]
rlabel metal3 1188 27948 1188 27948 0 chany_bottom_out[12]
rlabel metal1 24334 37094 24334 37094 0 chany_bottom_out[13]
rlabel via2 38226 30005 38226 30005 0 chany_bottom_out[14]
rlabel metal1 874 36346 874 36346 0 chany_bottom_out[15]
rlabel metal3 1188 1428 1188 1428 0 chany_bottom_out[16]
rlabel metal3 1188 15708 1188 15708 0 chany_bottom_out[17]
rlabel metal1 8786 2822 8786 2822 0 chany_bottom_out[18]
rlabel metal1 19550 37094 19550 37094 0 chany_bottom_out[1]
rlabel metal1 15594 37094 15594 37094 0 chany_bottom_out[2]
rlabel metal2 38226 8857 38226 8857 0 chany_bottom_out[3]
rlabel metal1 25346 37094 25346 37094 0 chany_bottom_out[4]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[5]
rlabel metal2 34822 1520 34822 1520 0 chany_bottom_out[6]
rlabel metal3 1188 17748 1188 17748 0 chany_bottom_out[7]
rlabel via2 38226 35445 38226 35445 0 chany_bottom_out[8]
rlabel metal2 25162 1520 25162 1520 0 chany_bottom_out[9]
rlabel via2 1610 21131 1610 21131 0 chany_top_in[0]
rlabel metal1 37582 2482 37582 2482 0 chany_top_in[10]
rlabel via2 38318 15691 38318 15691 0 chany_top_in[11]
rlabel metal2 4554 1299 4554 1299 0 chany_top_in[12]
rlabel metal2 1702 13787 1702 13787 0 chany_top_in[13]
rlabel via2 1610 31365 1610 31365 0 chany_top_in[14]
rlabel metal1 28750 2448 28750 2448 0 chany_top_in[15]
rlabel metal2 1610 29903 1610 29903 0 chany_top_in[16]
rlabel metal2 7130 38260 7130 38260 0 chany_top_in[17]
rlabel metal1 3634 2414 3634 2414 0 chany_top_in[18]
rlabel metal2 11086 3468 11086 3468 0 chany_top_in[1]
rlabel metal1 33902 2414 33902 2414 0 chany_top_in[2]
rlabel via2 38318 14365 38318 14365 0 chany_top_in[3]
rlabel via2 38318 6885 38318 6885 0 chany_top_in[4]
rlabel metal3 1142 6868 1142 6868 0 chany_top_in[5]
rlabel via2 1702 36771 1702 36771 0 chany_top_in[6]
rlabel metal3 38786 68 38786 68 0 chany_top_in[7]
rlabel via2 1702 8891 1702 8891 0 chany_top_in[8]
rlabel metal2 38318 11033 38318 11033 0 chany_top_in[9]
rlabel metal3 1188 24548 1188 24548 0 chany_top_out[0]
rlabel metal2 29670 1520 29670 1520 0 chany_top_out[10]
rlabel via2 38226 24565 38226 24565 0 chany_top_out[11]
rlabel metal1 10442 37094 10442 37094 0 chany_top_out[12]
rlabel metal1 5336 37094 5336 37094 0 chany_top_out[13]
rlabel metal2 18078 1299 18078 1299 0 chany_top_out[14]
rlabel metal2 46 1656 46 1656 0 chany_top_out[15]
rlabel metal1 23552 3366 23552 3366 0 chany_top_out[16]
rlabel metal2 12374 37094 12374 37094 0 chany_top_out[17]
rlabel metal1 22172 37094 22172 37094 0 chany_top_out[18]
rlabel metal1 33672 37094 33672 37094 0 chany_top_out[1]
rlabel metal3 1188 26588 1188 26588 0 chany_top_out[2]
rlabel metal3 1188 22508 1188 22508 0 chany_top_out[3]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[4]
rlabel metal1 37536 37094 37536 37094 0 chany_top_out[5]
rlabel metal1 29486 37094 29486 37094 0 chany_top_out[6]
rlabel metal1 16928 3910 16928 3910 0 chany_top_out[7]
rlabel metal2 36754 38131 36754 38131 0 chany_top_out[8]
rlabel metal2 38226 3417 38226 3417 0 chany_top_out[9]
rlabel metal3 1188 10268 1188 10268 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal2 38226 21233 38226 21233 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal2 6486 1520 6486 1520 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal1 15870 14994 15870 14994 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal2 14444 13396 14444 13396 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 17434 15470 17434 15470 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal1 21344 7378 21344 7378 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal2 24886 4930 24886 4930 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal1 23598 8942 23598 8942 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal2 18630 7480 18630 7480 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal1 13662 14994 13662 14994 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal1 15364 2482 15364 2482 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal1 16836 2482 16836 2482 0 mem_left_ipin_1.DFFR_3_.Q
rlabel via1 16514 6154 16514 6154 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal2 18906 6630 18906 6630 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal2 21942 2873 21942 2873 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal2 26266 8874 26266 8874 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 22540 9078 22540 9078 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal2 21850 5627 21850 5627 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal1 19688 6358 19688 6358 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal2 22402 5610 22402 5610 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal1 29118 7378 29118 7378 0 mem_left_ipin_3.DFFR_0_.Q
rlabel metal1 29486 7378 29486 7378 0 mem_left_ipin_3.DFFR_1_.Q
rlabel metal1 19964 8330 19964 8330 0 mem_left_ipin_3.DFFR_2_.Q
rlabel metal1 22310 3128 22310 3128 0 mem_left_ipin_3.DFFR_3_.Q
rlabel metal1 25024 3434 25024 3434 0 mem_left_ipin_3.DFFR_4_.Q
rlabel metal1 26358 3400 26358 3400 0 mem_left_ipin_3.DFFR_5_.Q
rlabel metal2 20838 14722 20838 14722 0 mem_left_ipin_4.DFFR_0_.Q
rlabel metal1 14122 12920 14122 12920 0 mem_left_ipin_4.DFFR_1_.Q
rlabel metal1 14122 15470 14122 15470 0 mem_left_ipin_4.DFFR_2_.Q
rlabel metal1 15962 6834 15962 6834 0 mem_left_ipin_4.DFFR_3_.Q
rlabel metal1 13478 10030 13478 10030 0 mem_left_ipin_4.DFFR_4_.Q
rlabel metal1 12650 9486 12650 9486 0 mem_left_ipin_4.DFFR_5_.Q
rlabel metal1 19228 14994 19228 14994 0 mem_left_ipin_5.DFFR_0_.Q
rlabel metal1 23552 9622 23552 9622 0 mem_left_ipin_5.DFFR_1_.Q
rlabel metal1 20884 10234 20884 10234 0 mem_left_ipin_5.DFFR_2_.Q
rlabel metal2 18906 10302 18906 10302 0 mem_left_ipin_5.DFFR_3_.Q
rlabel metal1 20755 9350 20755 9350 0 mem_left_ipin_5.DFFR_4_.Q
rlabel metal1 18722 9350 18722 9350 0 mem_left_ipin_5.DFFR_5_.Q
rlabel metal2 16238 16252 16238 16252 0 mem_left_ipin_6.DFFR_0_.Q
rlabel metal1 17802 16048 17802 16048 0 mem_left_ipin_6.DFFR_1_.Q
rlabel metal2 12282 14212 12282 14212 0 mem_left_ipin_6.DFFR_2_.Q
rlabel metal1 13800 5814 13800 5814 0 mem_left_ipin_6.DFFR_3_.Q
rlabel metal1 18860 2346 18860 2346 0 mem_left_ipin_6.DFFR_4_.Q
rlabel metal1 17020 2550 17020 2550 0 mem_left_ipin_6.DFFR_5_.Q
rlabel metal2 8970 4828 8970 4828 0 mem_left_ipin_7.DFFR_0_.Q
rlabel metal1 10764 14042 10764 14042 0 mem_left_ipin_7.DFFR_1_.Q
rlabel metal1 12006 14994 12006 14994 0 mem_left_ipin_7.DFFR_2_.Q
rlabel metal1 12144 2550 12144 2550 0 mem_left_ipin_7.DFFR_3_.Q
rlabel metal1 13662 3570 13662 3570 0 mem_left_ipin_7.DFFR_4_.Q
rlabel metal2 13570 3298 13570 3298 0 mem_left_ipin_7.DFFR_5_.Q
rlabel metal1 14398 14994 14398 14994 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal1 17342 7446 17342 7446 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 14582 5134 14582 5134 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal1 11960 5270 11960 5270 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal2 16054 5168 16054 5168 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal2 14582 4250 14582 4250 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal1 29946 7786 29946 7786 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal2 30406 9299 30406 9299 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal1 22908 2482 22908 2482 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal1 24196 2482 24196 2482 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 27922 4250 27922 4250 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal1 24794 2958 24794 2958 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 31418 2414 31418 2414 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal2 33350 3451 33350 3451 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 19826 2312 19826 2312 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal1 21252 2550 21252 2550 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal2 25990 4998 25990 4998 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal2 21482 16218 21482 16218 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 20424 16082 20424 16082 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 19964 26282 19964 26282 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal2 15962 14892 15962 14892 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 18262 26758 18262 26758 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal2 10718 15844 10718 15844 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 15824 26758 15824 26758 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal1 14076 13838 14076 13838 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal1 20516 15878 20516 15878 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 17710 14212 17710 14212 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17526 14688 17526 14688 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 37490 21862 37490 21862 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 21666 11832 21666 11832 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 17526 12920 17526 12920 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal1 13892 10574 13892 10574 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal1 15318 10574 15318 10574 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal1 12144 12750 12144 12750 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal1 13478 13838 13478 13838 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal2 21206 13192 21206 13192 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16882 9486 16882 9486 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 12742 11492 12742 11492 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 31050 2482 31050 2482 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 24978 12750 24978 12750 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal1 26588 12206 26588 12206 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal1 26312 12818 26312 12818 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal1 26910 10098 26910 10098 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal2 21574 14042 21574 14042 0 mux_left_ipin_2.INVTX1_6_.out
rlabel metal1 20424 13362 20424 13362 0 mux_left_ipin_2.INVTX1_7_.out
rlabel metal1 24656 12954 24656 12954 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 26082 12954 26082 12954 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 22172 13362 22172 13362 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 30912 28050 30912 28050 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17986 12750 17986 12750 0 mux_left_ipin_3.INVTX1_2_.out
rlabel metal2 28842 13396 28842 13396 0 mux_left_ipin_3.INVTX1_3_.out
rlabel metal1 28382 7310 28382 7310 0 mux_left_ipin_3.INVTX1_4_.out
rlabel metal2 28382 5100 28382 5100 0 mux_left_ipin_3.INVTX1_5_.out
rlabel metal1 29210 8942 29210 8942 0 mux_left_ipin_3.INVTX1_6_.out
rlabel metal2 26910 7650 26910 7650 0 mux_left_ipin_3.INVTX1_7_.out
rlabel metal2 23598 10948 23598 10948 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 27922 8398 27922 8398 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 27370 8806 27370 8806 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 31188 29138 31188 29138 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 24702 15538 24702 15538 0 mux_left_ipin_4.INVTX1_2_.out
rlabel metal1 25208 13362 25208 13362 0 mux_left_ipin_4.INVTX1_3_.out
rlabel metal1 29072 2958 29072 2958 0 mux_left_ipin_4.INVTX1_4_.out
rlabel metal1 26036 2414 26036 2414 0 mux_left_ipin_4.INVTX1_5_.out
rlabel metal1 20286 13158 20286 13158 0 mux_left_ipin_4.INVTX1_6_.out
rlabel metal2 7774 13328 7774 13328 0 mux_left_ipin_4.INVTX1_7_.out
rlabel metal1 18446 12886 18446 12886 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21735 10098 21735 10098 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15962 13804 15962 13804 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel via2 10534 31773 10534 31773 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22310 27302 22310 27302 0 mux_left_ipin_5.INVTX1_2_.out
rlabel metal1 23506 16966 23506 16966 0 mux_left_ipin_5.INVTX1_3_.out
rlabel metal2 33074 18394 33074 18394 0 mux_left_ipin_5.INVTX1_4_.out
rlabel metal2 32982 16660 32982 16660 0 mux_left_ipin_5.INVTX1_5_.out
rlabel metal1 19412 30022 19412 30022 0 mux_left_ipin_5.INVTX1_6_.out
rlabel metal2 15502 16116 15502 16116 0 mux_left_ipin_5.INVTX1_7_.out
rlabel metal2 23966 17510 23966 17510 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 25208 16490 25208 16490 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19550 17850 19550 17850 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14766 26350 14766 26350 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 21528 16490 21528 16490 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 17250 13770 17250 13770 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 15042 15028 15042 15028 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 20102 10982 20102 10982 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19412 13838 19412 13838 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16422 11084 16422 11084 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 12650 13838 12650 13838 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 12650 12002 12650 12002 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 13754 11050 13754 11050 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20378 10608 20378 10608 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15778 12716 15778 12716 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 15272 11118 15272 11118 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 25622 10778 25622 10778 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 27186 8772 27186 8772 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 27922 9894 27922 9894 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 29900 9622 29900 9622 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 20148 9078 20148 9078 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 25208 4454 25208 4454 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19964 11730 19964 11730 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 12466 3927 12466 3927 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 37720 26894 37720 26894 0 net1
rlabel metal1 20148 37162 20148 37162 0 net10
rlabel metal1 29578 10098 29578 10098 0 net100
rlabel metal2 18906 8874 18906 8874 0 net101
rlabel metal2 20562 37128 20562 37128 0 net11
rlabel metal1 34040 25874 34040 25874 0 net12
rlabel metal1 9154 21862 9154 21862 0 net13
rlabel metal1 1932 5202 1932 5202 0 net14
rlabel via1 26197 33286 26197 33286 0 net15
rlabel metal1 22816 27438 22816 27438 0 net16
rlabel metal2 2990 37536 2990 37536 0 net17
rlabel metal1 9844 13226 9844 13226 0 net18
rlabel metal1 37766 24922 37766 24922 0 net19
rlabel metal1 21114 24786 21114 24786 0 net2
rlabel metal1 10074 2550 10074 2550 0 net20
rlabel metal2 1886 20910 1886 20910 0 net21
rlabel metal2 37766 2176 37766 2176 0 net22
rlabel metal2 37858 20672 37858 20672 0 net23
rlabel metal1 2208 23086 2208 23086 0 net24
rlabel metal1 20700 29138 20700 29138 0 net25
rlabel metal1 16560 31858 16560 31858 0 net26
rlabel metal2 25530 28798 25530 28798 0 net27
rlabel metal2 2530 13022 2530 13022 0 net28
rlabel metal1 4554 14994 4554 14994 0 net29
rlabel metal2 38134 3808 38134 3808 0 net3
rlabel metal1 10166 3026 10166 3026 0 net30
rlabel metal1 17986 33966 17986 33966 0 net31
rlabel metal1 22494 32402 22494 32402 0 net32
rlabel metal1 36961 12886 36961 12886 0 net33
rlabel metal1 36984 7378 36984 7378 0 net34
rlabel metal1 25024 24174 25024 24174 0 net35
rlabel metal2 1794 36448 1794 36448 0 net36
rlabel metal1 15042 15028 15042 15028 0 net37
rlabel metal2 1886 10030 1886 10030 0 net38
rlabel metal1 28888 3502 28888 3502 0 net39
rlabel metal2 38134 19210 38134 19210 0 net4
rlabel metal2 8050 3094 8050 3094 0 net40
rlabel metal1 37812 36142 37812 36142 0 net41
rlabel metal2 34178 26758 34178 26758 0 net42
rlabel metal1 17388 37230 17388 37230 0 net43
rlabel metal1 38134 25466 38134 25466 0 net44
rlabel metal1 1840 23290 1840 23290 0 net45
rlabel metal1 22586 29274 22586 29274 0 net46
rlabel metal2 38042 30532 38042 30532 0 net47
rlabel metal1 3680 36142 3680 36142 0 net48
rlabel metal2 1886 4963 1886 4963 0 net49
rlabel metal1 20470 36686 20470 36686 0 net5
rlabel metal2 4094 15606 4094 15606 0 net50
rlabel metal2 8970 3196 8970 3196 0 net51
rlabel metal1 18952 37230 18952 37230 0 net52
rlabel metal2 15870 34714 15870 34714 0 net53
rlabel metal2 38042 9690 38042 9690 0 net54
rlabel metal1 25300 36686 25300 36686 0 net55
rlabel metal2 25254 30770 25254 30770 0 net56
rlabel metal1 35328 2414 35328 2414 0 net57
rlabel metal2 1886 16558 1886 16558 0 net58
rlabel metal1 37766 35666 37766 35666 0 net59
rlabel metal1 5014 32810 5014 32810 0 net6
rlabel metal1 26726 2414 26726 2414 0 net60
rlabel metal1 2162 24786 2162 24786 0 net61
rlabel metal1 29348 2414 29348 2414 0 net62
rlabel metal1 38088 21114 38088 21114 0 net63
rlabel metal1 12144 36890 12144 36890 0 net64
rlabel metal1 5244 33082 5244 33082 0 net65
rlabel metal2 12650 3451 12650 3451 0 net66
rlabel metal1 4048 2482 4048 2482 0 net67
rlabel metal1 24058 3434 24058 3434 0 net68
rlabel metal1 14720 36890 14720 36890 0 net69
rlabel metal1 1932 19346 1932 19346 0 net7
rlabel metal2 21298 37060 21298 37060 0 net70
rlabel metal2 33626 31620 33626 31620 0 net71
rlabel metal1 4370 26962 4370 26962 0 net72
rlabel metal1 1840 22610 1840 22610 0 net73
rlabel metal1 2162 2414 2162 2414 0 net74
rlabel metal2 37490 36958 37490 36958 0 net75
rlabel metal1 25254 36584 25254 36584 0 net76
rlabel metal1 12834 3978 12834 3978 0 net77
rlabel metal1 37398 26554 37398 26554 0 net78
rlabel metal1 38042 3570 38042 3570 0 net79
rlabel metal1 33534 5134 33534 5134 0 net8
rlabel metal2 9430 10438 9430 10438 0 net80
rlabel metal2 38042 18598 38042 18598 0 net81
rlabel metal1 6854 2448 6854 2448 0 net82
rlabel metal1 37996 22746 37996 22746 0 net83
rlabel metal2 30590 2142 30590 2142 0 net84
rlabel metal1 31510 37162 31510 37162 0 net85
rlabel metal1 30820 29274 30820 29274 0 net86
rlabel metal1 4278 37196 4278 37196 0 net87
rlabel metal1 11914 26554 11914 26554 0 net88
rlabel metal2 27186 2244 27186 2244 0 net89
rlabel metal1 36110 12750 36110 12750 0 net9
rlabel metal1 3726 12818 3726 12818 0 net90
rlabel metal1 16652 14926 16652 14926 0 net91
rlabel metal1 11500 10574 11500 10574 0 net92
rlabel metal2 25254 14688 25254 14688 0 net93
rlabel metal2 29762 9282 29762 9282 0 net94
rlabel metal2 14858 16864 14858 16864 0 net95
rlabel metal2 19458 18020 19458 18020 0 net96
rlabel metal1 13754 14314 13754 14314 0 net97
rlabel metal1 10902 14314 10902 14314 0 net98
rlabel metal1 11178 12716 11178 12716 0 net99
rlabel metal2 12926 823 12926 823 0 pReset
rlabel metal1 7222 2618 7222 2618 0 prog_clk
rlabel metal2 38226 23341 38226 23341 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 21298 2064 21298 2064 0 right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 32384 37094 32384 37094 0 right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 30498 37094 30498 37094 0 right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 4002 37094 4002 37094 0 right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal1 8832 37094 8832 37094 0 right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal2 26450 1520 26450 1520 0 right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal3 1188 12308 1188 12308 0 right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
