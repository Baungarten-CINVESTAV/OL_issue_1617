VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_4__4_
  CLASS BLOCK ;
  FOREIGN sb_4__4_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 30.640 199.000 31.240 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 166.640 199.000 167.240 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 199.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 199.000 191.040 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 61.240 4.000 61.840 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1.000 174.250 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.640 4.000 184.240 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 196.000 190.350 199.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1.000 145.270 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 37.440 4.000 38.040 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 153.040 4.000 153.640 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1.000 51.890 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1.000 22.910 4.000 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 102.040 4.000 102.640 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 88.440 4.000 89.040 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.840 199.000 143.440 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 196.000 90.530 199.000 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1.000 167.810 4.000 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.840 4.000 126.440 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 159.840 4.000 160.440 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1.000 113.070 4.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1.000 74.430 4.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1.000 196.790 4.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 6.840 4.000 7.440 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.040 199.000 102.640 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 196.000 122.730 199.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 199.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 199.000 184.240 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 1.000 84.090 4.000 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 78.240 4.000 78.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 173.440 199.000 174.040 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 199.000 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.240 199.000 44.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 199.000 61.840 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 196.000 84.090 199.000 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 196.000 51.890 199.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1.000 45.450 4.000 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 199.000 150.240 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1.000 190.350 4.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 199.000 78.840 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 196.000 145.270 199.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 199.000 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 199.000 7.440 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.840 199.000 160.440 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 196.000 183.910 199.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 196.000 106.630 199.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 95.240 4.000 95.840 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 199.000 38.040 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 112.240 4.000 112.840 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 13.640 4.000 14.240 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 196.000 129.170 199.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 142.840 4.000 143.440 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1.000 151.710 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 196.000 167.810 199.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 47.640 4.000 48.240 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1.000 13.250 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1.000 58.330 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 85.040 199.000 85.640 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 199.000 55.040 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 30.640 4.000 31.240 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 166.640 4.000 167.240 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 199.000 14.240 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 199.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 199.000 72.040 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 199.000 126.440 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1.000 158.150 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 199.000 136.640 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 196.000 29.350 199.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 119.040 4.000 119.640 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1.000 96.970 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1.000 119.510 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 196.000 39.010 199.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 199.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 23.840 4.000 24.440 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 196.000 0.370 199.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1.000 29.350 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1.000 6.810 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 196.000 174.250 199.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 196.000 138.830 199.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1.000 90.530 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 199.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 199.000 21.040 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 196.000 6.810 199.000 ;
    END
  END chany_bottom_out[9]
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 199.000 109.440 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1.000 35.790 4.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1.000 67.990 4.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 71.440 4.000 72.040 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 199.000 119.640 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1.000 106.630 4.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 196.000 161.370 199.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 196.000 151.710 199.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 199.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 196.000 45.450 199.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1.000 135.610 4.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.440 4.000 55.040 ;
    END
  END prog_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 176.840 4.000 177.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 199.000 95.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 0.070 10.640 196.810 187.920 ;
      LAYER met2 ;
        RECT 0.650 195.720 6.250 196.000 ;
        RECT 7.090 195.720 15.910 196.000 ;
        RECT 16.750 195.720 22.350 196.000 ;
        RECT 23.190 195.720 28.790 196.000 ;
        RECT 29.630 195.720 38.450 196.000 ;
        RECT 39.290 195.720 44.890 196.000 ;
        RECT 45.730 195.720 51.330 196.000 ;
        RECT 52.170 195.720 60.990 196.000 ;
        RECT 61.830 195.720 67.430 196.000 ;
        RECT 68.270 195.720 77.090 196.000 ;
        RECT 77.930 195.720 83.530 196.000 ;
        RECT 84.370 195.720 89.970 196.000 ;
        RECT 90.810 195.720 99.630 196.000 ;
        RECT 100.470 195.720 106.070 196.000 ;
        RECT 106.910 195.720 112.510 196.000 ;
        RECT 113.350 195.720 122.170 196.000 ;
        RECT 123.010 195.720 128.610 196.000 ;
        RECT 129.450 195.720 138.270 196.000 ;
        RECT 139.110 195.720 144.710 196.000 ;
        RECT 145.550 195.720 151.150 196.000 ;
        RECT 151.990 195.720 160.810 196.000 ;
        RECT 161.650 195.720 167.250 196.000 ;
        RECT 168.090 195.720 173.690 196.000 ;
        RECT 174.530 195.720 183.350 196.000 ;
        RECT 184.190 195.720 189.790 196.000 ;
        RECT 190.630 195.720 196.230 196.000 ;
        RECT 0.100 4.280 196.780 195.720 ;
        RECT 0.650 4.000 6.250 4.280 ;
        RECT 7.090 4.000 12.690 4.280 ;
        RECT 13.530 4.000 22.350 4.280 ;
        RECT 23.190 4.000 28.790 4.280 ;
        RECT 29.630 4.000 35.230 4.280 ;
        RECT 36.070 4.000 44.890 4.280 ;
        RECT 45.730 4.000 51.330 4.280 ;
        RECT 52.170 4.000 57.770 4.280 ;
        RECT 58.610 4.000 67.430 4.280 ;
        RECT 68.270 4.000 73.870 4.280 ;
        RECT 74.710 4.000 83.530 4.280 ;
        RECT 84.370 4.000 89.970 4.280 ;
        RECT 90.810 4.000 96.410 4.280 ;
        RECT 97.250 4.000 106.070 4.280 ;
        RECT 106.910 4.000 112.510 4.280 ;
        RECT 113.350 4.000 118.950 4.280 ;
        RECT 119.790 4.000 128.610 4.280 ;
        RECT 129.450 4.000 135.050 4.280 ;
        RECT 135.890 4.000 144.710 4.280 ;
        RECT 145.550 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.590 4.280 ;
        RECT 158.430 4.000 167.250 4.280 ;
        RECT 168.090 4.000 173.690 4.280 ;
        RECT 174.530 4.000 180.130 4.280 ;
        RECT 180.970 4.000 189.790 4.280 ;
        RECT 190.630 4.000 196.230 4.280 ;
      LAYER met3 ;
        RECT 4.400 190.040 195.600 190.905 ;
        RECT 4.000 184.640 196.000 190.040 ;
        RECT 4.400 183.240 195.600 184.640 ;
        RECT 4.000 177.840 196.000 183.240 ;
        RECT 4.400 176.440 196.000 177.840 ;
        RECT 4.000 174.440 196.000 176.440 ;
        RECT 4.000 173.040 195.600 174.440 ;
        RECT 4.000 167.640 196.000 173.040 ;
        RECT 4.400 166.240 195.600 167.640 ;
        RECT 4.000 160.840 196.000 166.240 ;
        RECT 4.400 159.440 195.600 160.840 ;
        RECT 4.000 154.040 196.000 159.440 ;
        RECT 4.400 152.640 196.000 154.040 ;
        RECT 4.000 150.640 196.000 152.640 ;
        RECT 4.000 149.240 195.600 150.640 ;
        RECT 4.000 143.840 196.000 149.240 ;
        RECT 4.400 142.440 195.600 143.840 ;
        RECT 4.000 137.040 196.000 142.440 ;
        RECT 4.400 135.640 195.600 137.040 ;
        RECT 4.000 126.840 196.000 135.640 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 4.000 120.040 196.000 125.440 ;
        RECT 4.400 118.640 195.600 120.040 ;
        RECT 4.000 113.240 196.000 118.640 ;
        RECT 4.400 111.840 196.000 113.240 ;
        RECT 4.000 109.840 196.000 111.840 ;
        RECT 4.000 108.440 195.600 109.840 ;
        RECT 4.000 103.040 196.000 108.440 ;
        RECT 4.400 101.640 195.600 103.040 ;
        RECT 4.000 96.240 196.000 101.640 ;
        RECT 4.400 94.840 195.600 96.240 ;
        RECT 4.000 89.440 196.000 94.840 ;
        RECT 4.400 88.040 196.000 89.440 ;
        RECT 4.000 86.040 196.000 88.040 ;
        RECT 4.000 84.640 195.600 86.040 ;
        RECT 4.000 79.240 196.000 84.640 ;
        RECT 4.400 77.840 195.600 79.240 ;
        RECT 4.000 72.440 196.000 77.840 ;
        RECT 4.400 71.040 195.600 72.440 ;
        RECT 4.000 62.240 196.000 71.040 ;
        RECT 4.400 60.840 195.600 62.240 ;
        RECT 4.000 55.440 196.000 60.840 ;
        RECT 4.400 54.040 195.600 55.440 ;
        RECT 4.000 48.640 196.000 54.040 ;
        RECT 4.400 47.240 196.000 48.640 ;
        RECT 4.000 45.240 196.000 47.240 ;
        RECT 4.000 43.840 195.600 45.240 ;
        RECT 4.000 38.440 196.000 43.840 ;
        RECT 4.400 37.040 195.600 38.440 ;
        RECT 4.000 31.640 196.000 37.040 ;
        RECT 4.400 30.240 195.600 31.640 ;
        RECT 4.000 24.840 196.000 30.240 ;
        RECT 4.400 23.440 196.000 24.840 ;
        RECT 4.000 21.440 196.000 23.440 ;
        RECT 4.000 20.040 195.600 21.440 ;
        RECT 4.000 14.640 196.000 20.040 ;
        RECT 4.400 13.240 195.600 14.640 ;
        RECT 4.000 7.840 196.000 13.240 ;
        RECT 4.400 6.975 195.600 7.840 ;
      LAYER met4 ;
        RECT 10.415 19.895 20.640 158.945 ;
        RECT 23.040 19.895 77.905 158.945 ;
  END
END sb_4__4_
END LIBRARY

