magic
tech sky130A
magscale 1 2
timestamp 1672604766
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 14 2128 582820 701808
<< metal2 >>
rect 662 703200 718 703800
rect 4526 703200 4582 703800
rect 8390 703200 8446 703800
rect 12254 703200 12310 703800
rect 16118 703200 16174 703800
rect 19982 703200 20038 703800
rect 23846 703200 23902 703800
rect 27710 703200 27766 703800
rect 31574 703200 31630 703800
rect 35438 703200 35494 703800
rect 39946 703200 40002 703800
rect 43810 703200 43866 703800
rect 47674 703200 47730 703800
rect 51538 703200 51594 703800
rect 55402 703200 55458 703800
rect 59266 703200 59322 703800
rect 63130 703200 63186 703800
rect 66994 703200 67050 703800
rect 70858 703200 70914 703800
rect 74722 703200 74778 703800
rect 79230 703200 79286 703800
rect 83094 703200 83150 703800
rect 86958 703200 87014 703800
rect 90822 703200 90878 703800
rect 94686 703200 94742 703800
rect 98550 703200 98606 703800
rect 102414 703200 102470 703800
rect 106278 703200 106334 703800
rect 110142 703200 110198 703800
rect 114006 703200 114062 703800
rect 118514 703200 118570 703800
rect 122378 703200 122434 703800
rect 126242 703200 126298 703800
rect 130106 703200 130162 703800
rect 133970 703200 134026 703800
rect 137834 703200 137890 703800
rect 141698 703200 141754 703800
rect 145562 703200 145618 703800
rect 149426 703200 149482 703800
rect 153290 703200 153346 703800
rect 157798 703200 157854 703800
rect 161662 703200 161718 703800
rect 165526 703200 165582 703800
rect 169390 703200 169446 703800
rect 173254 703200 173310 703800
rect 177118 703200 177174 703800
rect 180982 703200 181038 703800
rect 184846 703200 184902 703800
rect 188710 703200 188766 703800
rect 193218 703200 193274 703800
rect 197082 703200 197138 703800
rect 200946 703200 201002 703800
rect 204810 703200 204866 703800
rect 208674 703200 208730 703800
rect 212538 703200 212594 703800
rect 216402 703200 216458 703800
rect 220266 703200 220322 703800
rect 224130 703200 224186 703800
rect 227994 703200 228050 703800
rect 232502 703200 232558 703800
rect 236366 703200 236422 703800
rect 240230 703200 240286 703800
rect 244094 703200 244150 703800
rect 247958 703200 248014 703800
rect 251822 703200 251878 703800
rect 255686 703200 255742 703800
rect 259550 703200 259606 703800
rect 263414 703200 263470 703800
rect 267278 703200 267334 703800
rect 271786 703200 271842 703800
rect 275650 703200 275706 703800
rect 279514 703200 279570 703800
rect 283378 703200 283434 703800
rect 287242 703200 287298 703800
rect 291106 703200 291162 703800
rect 294970 703200 295026 703800
rect 298834 703200 298890 703800
rect 302698 703200 302754 703800
rect 306562 703200 306618 703800
rect 311070 703200 311126 703800
rect 314934 703200 314990 703800
rect 318798 703200 318854 703800
rect 322662 703200 322718 703800
rect 326526 703200 326582 703800
rect 330390 703200 330446 703800
rect 334254 703200 334310 703800
rect 338118 703200 338174 703800
rect 341982 703200 342038 703800
rect 345846 703200 345902 703800
rect 350354 703200 350410 703800
rect 354218 703200 354274 703800
rect 358082 703200 358138 703800
rect 361946 703200 362002 703800
rect 365810 703200 365866 703800
rect 369674 703200 369730 703800
rect 373538 703200 373594 703800
rect 377402 703200 377458 703800
rect 381266 703200 381322 703800
rect 385130 703200 385186 703800
rect 389638 703200 389694 703800
rect 393502 703200 393558 703800
rect 397366 703200 397422 703800
rect 401230 703200 401286 703800
rect 405094 703200 405150 703800
rect 408958 703200 409014 703800
rect 412822 703200 412878 703800
rect 416686 703200 416742 703800
rect 420550 703200 420606 703800
rect 424414 703200 424470 703800
rect 428922 703200 428978 703800
rect 432786 703200 432842 703800
rect 436650 703200 436706 703800
rect 440514 703200 440570 703800
rect 444378 703200 444434 703800
rect 448242 703200 448298 703800
rect 452106 703200 452162 703800
rect 455970 703200 456026 703800
rect 459834 703200 459890 703800
rect 463698 703200 463754 703800
rect 468206 703200 468262 703800
rect 472070 703200 472126 703800
rect 475934 703200 475990 703800
rect 479798 703200 479854 703800
rect 483662 703200 483718 703800
rect 487526 703200 487582 703800
rect 491390 703200 491446 703800
rect 495254 703200 495310 703800
rect 499118 703200 499174 703800
rect 502982 703200 503038 703800
rect 507490 703200 507546 703800
rect 511354 703200 511410 703800
rect 515218 703200 515274 703800
rect 519082 703200 519138 703800
rect 522946 703200 523002 703800
rect 526810 703200 526866 703800
rect 530674 703200 530730 703800
rect 534538 703200 534594 703800
rect 538402 703200 538458 703800
rect 542266 703200 542322 703800
rect 546774 703200 546830 703800
rect 550638 703200 550694 703800
rect 554502 703200 554558 703800
rect 558366 703200 558422 703800
rect 562230 703200 562286 703800
rect 566094 703200 566150 703800
rect 569958 703200 570014 703800
rect 573822 703200 573878 703800
rect 577686 703200 577742 703800
rect 581550 703200 581606 703800
rect 18 200 74 800
rect 3882 200 3938 800
rect 7746 200 7802 800
rect 11610 200 11666 800
rect 15474 200 15530 800
rect 19338 200 19394 800
rect 23202 200 23258 800
rect 27066 200 27122 800
rect 30930 200 30986 800
rect 34794 200 34850 800
rect 39302 200 39358 800
rect 43166 200 43222 800
rect 47030 200 47086 800
rect 50894 200 50950 800
rect 54758 200 54814 800
rect 58622 200 58678 800
rect 62486 200 62542 800
rect 66350 200 66406 800
rect 70214 200 70270 800
rect 74078 200 74134 800
rect 78586 200 78642 800
rect 82450 200 82506 800
rect 86314 200 86370 800
rect 90178 200 90234 800
rect 94042 200 94098 800
rect 97906 200 97962 800
rect 101770 200 101826 800
rect 105634 200 105690 800
rect 109498 200 109554 800
rect 113362 200 113418 800
rect 117870 200 117926 800
rect 121734 200 121790 800
rect 125598 200 125654 800
rect 129462 200 129518 800
rect 133326 200 133382 800
rect 137190 200 137246 800
rect 141054 200 141110 800
rect 144918 200 144974 800
rect 148782 200 148838 800
rect 152646 200 152702 800
rect 157154 200 157210 800
rect 161018 200 161074 800
rect 164882 200 164938 800
rect 168746 200 168802 800
rect 172610 200 172666 800
rect 176474 200 176530 800
rect 180338 200 180394 800
rect 184202 200 184258 800
rect 188066 200 188122 800
rect 191930 200 191986 800
rect 196438 200 196494 800
rect 200302 200 200358 800
rect 204166 200 204222 800
rect 208030 200 208086 800
rect 211894 200 211950 800
rect 215758 200 215814 800
rect 219622 200 219678 800
rect 223486 200 223542 800
rect 227350 200 227406 800
rect 231214 200 231270 800
rect 235722 200 235778 800
rect 239586 200 239642 800
rect 243450 200 243506 800
rect 247314 200 247370 800
rect 251178 200 251234 800
rect 255042 200 255098 800
rect 258906 200 258962 800
rect 262770 200 262826 800
rect 266634 200 266690 800
rect 270498 200 270554 800
rect 275006 200 275062 800
rect 278870 200 278926 800
rect 282734 200 282790 800
rect 286598 200 286654 800
rect 290462 200 290518 800
rect 294326 200 294382 800
rect 298190 200 298246 800
rect 302054 200 302110 800
rect 305918 200 305974 800
rect 309782 200 309838 800
rect 314290 200 314346 800
rect 318154 200 318210 800
rect 322018 200 322074 800
rect 325882 200 325938 800
rect 329746 200 329802 800
rect 333610 200 333666 800
rect 337474 200 337530 800
rect 341338 200 341394 800
rect 345202 200 345258 800
rect 349066 200 349122 800
rect 353574 200 353630 800
rect 357438 200 357494 800
rect 361302 200 361358 800
rect 365166 200 365222 800
rect 369030 200 369086 800
rect 372894 200 372950 800
rect 376758 200 376814 800
rect 380622 200 380678 800
rect 384486 200 384542 800
rect 388350 200 388406 800
rect 392858 200 392914 800
rect 396722 200 396778 800
rect 400586 200 400642 800
rect 404450 200 404506 800
rect 408314 200 408370 800
rect 412178 200 412234 800
rect 416042 200 416098 800
rect 419906 200 419962 800
rect 423770 200 423826 800
rect 427634 200 427690 800
rect 432142 200 432198 800
rect 436006 200 436062 800
rect 439870 200 439926 800
rect 443734 200 443790 800
rect 447598 200 447654 800
rect 451462 200 451518 800
rect 455326 200 455382 800
rect 459190 200 459246 800
rect 463054 200 463110 800
rect 466918 200 466974 800
rect 471426 200 471482 800
rect 475290 200 475346 800
rect 479154 200 479210 800
rect 483018 200 483074 800
rect 486882 200 486938 800
rect 490746 200 490802 800
rect 494610 200 494666 800
rect 498474 200 498530 800
rect 502338 200 502394 800
rect 506202 200 506258 800
rect 510710 200 510766 800
rect 514574 200 514630 800
rect 518438 200 518494 800
rect 522302 200 522358 800
rect 526166 200 526222 800
rect 530030 200 530086 800
rect 533894 200 533950 800
rect 537758 200 537814 800
rect 541622 200 541678 800
rect 545486 200 545542 800
rect 549994 200 550050 800
rect 553858 200 553914 800
rect 557722 200 557778 800
rect 561586 200 561642 800
rect 565450 200 565506 800
rect 569314 200 569370 800
rect 573178 200 573234 800
rect 577042 200 577098 800
rect 580906 200 580962 800
<< obsm2 >>
rect 20 703856 582658 703882
rect 20 703144 606 703856
rect 774 703144 4470 703856
rect 4638 703144 8334 703856
rect 8502 703144 12198 703856
rect 12366 703144 16062 703856
rect 16230 703144 19926 703856
rect 20094 703144 23790 703856
rect 23958 703144 27654 703856
rect 27822 703144 31518 703856
rect 31686 703144 35382 703856
rect 35550 703144 39890 703856
rect 40058 703144 43754 703856
rect 43922 703144 47618 703856
rect 47786 703144 51482 703856
rect 51650 703144 55346 703856
rect 55514 703144 59210 703856
rect 59378 703144 63074 703856
rect 63242 703144 66938 703856
rect 67106 703144 70802 703856
rect 70970 703144 74666 703856
rect 74834 703144 79174 703856
rect 79342 703144 83038 703856
rect 83206 703144 86902 703856
rect 87070 703144 90766 703856
rect 90934 703144 94630 703856
rect 94798 703144 98494 703856
rect 98662 703144 102358 703856
rect 102526 703144 106222 703856
rect 106390 703144 110086 703856
rect 110254 703144 113950 703856
rect 114118 703144 118458 703856
rect 118626 703144 122322 703856
rect 122490 703144 126186 703856
rect 126354 703144 130050 703856
rect 130218 703144 133914 703856
rect 134082 703144 137778 703856
rect 137946 703144 141642 703856
rect 141810 703144 145506 703856
rect 145674 703144 149370 703856
rect 149538 703144 153234 703856
rect 153402 703144 157742 703856
rect 157910 703144 161606 703856
rect 161774 703144 165470 703856
rect 165638 703144 169334 703856
rect 169502 703144 173198 703856
rect 173366 703144 177062 703856
rect 177230 703144 180926 703856
rect 181094 703144 184790 703856
rect 184958 703144 188654 703856
rect 188822 703144 193162 703856
rect 193330 703144 197026 703856
rect 197194 703144 200890 703856
rect 201058 703144 204754 703856
rect 204922 703144 208618 703856
rect 208786 703144 212482 703856
rect 212650 703144 216346 703856
rect 216514 703144 220210 703856
rect 220378 703144 224074 703856
rect 224242 703144 227938 703856
rect 228106 703144 232446 703856
rect 232614 703144 236310 703856
rect 236478 703144 240174 703856
rect 240342 703144 244038 703856
rect 244206 703144 247902 703856
rect 248070 703144 251766 703856
rect 251934 703144 255630 703856
rect 255798 703144 259494 703856
rect 259662 703144 263358 703856
rect 263526 703144 267222 703856
rect 267390 703144 271730 703856
rect 271898 703144 275594 703856
rect 275762 703144 279458 703856
rect 279626 703144 283322 703856
rect 283490 703144 287186 703856
rect 287354 703144 291050 703856
rect 291218 703144 294914 703856
rect 295082 703144 298778 703856
rect 298946 703144 302642 703856
rect 302810 703144 306506 703856
rect 306674 703144 311014 703856
rect 311182 703144 314878 703856
rect 315046 703144 318742 703856
rect 318910 703144 322606 703856
rect 322774 703144 326470 703856
rect 326638 703144 330334 703856
rect 330502 703144 334198 703856
rect 334366 703144 338062 703856
rect 338230 703144 341926 703856
rect 342094 703144 345790 703856
rect 345958 703144 350298 703856
rect 350466 703144 354162 703856
rect 354330 703144 358026 703856
rect 358194 703144 361890 703856
rect 362058 703144 365754 703856
rect 365922 703144 369618 703856
rect 369786 703144 373482 703856
rect 373650 703144 377346 703856
rect 377514 703144 381210 703856
rect 381378 703144 385074 703856
rect 385242 703144 389582 703856
rect 389750 703144 393446 703856
rect 393614 703144 397310 703856
rect 397478 703144 401174 703856
rect 401342 703144 405038 703856
rect 405206 703144 408902 703856
rect 409070 703144 412766 703856
rect 412934 703144 416630 703856
rect 416798 703144 420494 703856
rect 420662 703144 424358 703856
rect 424526 703144 428866 703856
rect 429034 703144 432730 703856
rect 432898 703144 436594 703856
rect 436762 703144 440458 703856
rect 440626 703144 444322 703856
rect 444490 703144 448186 703856
rect 448354 703144 452050 703856
rect 452218 703144 455914 703856
rect 456082 703144 459778 703856
rect 459946 703144 463642 703856
rect 463810 703144 468150 703856
rect 468318 703144 472014 703856
rect 472182 703144 475878 703856
rect 476046 703144 479742 703856
rect 479910 703144 483606 703856
rect 483774 703144 487470 703856
rect 487638 703144 491334 703856
rect 491502 703144 495198 703856
rect 495366 703144 499062 703856
rect 499230 703144 502926 703856
rect 503094 703144 507434 703856
rect 507602 703144 511298 703856
rect 511466 703144 515162 703856
rect 515330 703144 519026 703856
rect 519194 703144 522890 703856
rect 523058 703144 526754 703856
rect 526922 703144 530618 703856
rect 530786 703144 534482 703856
rect 534650 703144 538346 703856
rect 538514 703144 542210 703856
rect 542378 703144 546718 703856
rect 546886 703144 550582 703856
rect 550750 703144 554446 703856
rect 554614 703144 558310 703856
rect 558478 703144 562174 703856
rect 562342 703144 566038 703856
rect 566206 703144 569902 703856
rect 570070 703144 573766 703856
rect 573934 703144 577630 703856
rect 577798 703144 581494 703856
rect 581662 703144 582658 703856
rect 20 856 582658 703144
rect 130 734 3826 856
rect 3994 734 7690 856
rect 7858 734 11554 856
rect 11722 734 15418 856
rect 15586 734 19282 856
rect 19450 734 23146 856
rect 23314 734 27010 856
rect 27178 734 30874 856
rect 31042 734 34738 856
rect 34906 734 39246 856
rect 39414 734 43110 856
rect 43278 734 46974 856
rect 47142 734 50838 856
rect 51006 734 54702 856
rect 54870 734 58566 856
rect 58734 734 62430 856
rect 62598 734 66294 856
rect 66462 734 70158 856
rect 70326 734 74022 856
rect 74190 734 78530 856
rect 78698 734 82394 856
rect 82562 734 86258 856
rect 86426 734 90122 856
rect 90290 734 93986 856
rect 94154 734 97850 856
rect 98018 734 101714 856
rect 101882 734 105578 856
rect 105746 734 109442 856
rect 109610 734 113306 856
rect 113474 734 117814 856
rect 117982 734 121678 856
rect 121846 734 125542 856
rect 125710 734 129406 856
rect 129574 734 133270 856
rect 133438 734 137134 856
rect 137302 734 140998 856
rect 141166 734 144862 856
rect 145030 734 148726 856
rect 148894 734 152590 856
rect 152758 734 157098 856
rect 157266 734 160962 856
rect 161130 734 164826 856
rect 164994 734 168690 856
rect 168858 734 172554 856
rect 172722 734 176418 856
rect 176586 734 180282 856
rect 180450 734 184146 856
rect 184314 734 188010 856
rect 188178 734 191874 856
rect 192042 734 196382 856
rect 196550 734 200246 856
rect 200414 734 204110 856
rect 204278 734 207974 856
rect 208142 734 211838 856
rect 212006 734 215702 856
rect 215870 734 219566 856
rect 219734 734 223430 856
rect 223598 734 227294 856
rect 227462 734 231158 856
rect 231326 734 235666 856
rect 235834 734 239530 856
rect 239698 734 243394 856
rect 243562 734 247258 856
rect 247426 734 251122 856
rect 251290 734 254986 856
rect 255154 734 258850 856
rect 259018 734 262714 856
rect 262882 734 266578 856
rect 266746 734 270442 856
rect 270610 734 274950 856
rect 275118 734 278814 856
rect 278982 734 282678 856
rect 282846 734 286542 856
rect 286710 734 290406 856
rect 290574 734 294270 856
rect 294438 734 298134 856
rect 298302 734 301998 856
rect 302166 734 305862 856
rect 306030 734 309726 856
rect 309894 734 314234 856
rect 314402 734 318098 856
rect 318266 734 321962 856
rect 322130 734 325826 856
rect 325994 734 329690 856
rect 329858 734 333554 856
rect 333722 734 337418 856
rect 337586 734 341282 856
rect 341450 734 345146 856
rect 345314 734 349010 856
rect 349178 734 353518 856
rect 353686 734 357382 856
rect 357550 734 361246 856
rect 361414 734 365110 856
rect 365278 734 368974 856
rect 369142 734 372838 856
rect 373006 734 376702 856
rect 376870 734 380566 856
rect 380734 734 384430 856
rect 384598 734 388294 856
rect 388462 734 392802 856
rect 392970 734 396666 856
rect 396834 734 400530 856
rect 400698 734 404394 856
rect 404562 734 408258 856
rect 408426 734 412122 856
rect 412290 734 415986 856
rect 416154 734 419850 856
rect 420018 734 423714 856
rect 423882 734 427578 856
rect 427746 734 432086 856
rect 432254 734 435950 856
rect 436118 734 439814 856
rect 439982 734 443678 856
rect 443846 734 447542 856
rect 447710 734 451406 856
rect 451574 734 455270 856
rect 455438 734 459134 856
rect 459302 734 462998 856
rect 463166 734 466862 856
rect 467030 734 471370 856
rect 471538 734 475234 856
rect 475402 734 479098 856
rect 479266 734 482962 856
rect 483130 734 486826 856
rect 486994 734 490690 856
rect 490858 734 494554 856
rect 494722 734 498418 856
rect 498586 734 502282 856
rect 502450 734 506146 856
rect 506314 734 510654 856
rect 510822 734 514518 856
rect 514686 734 518382 856
rect 518550 734 522246 856
rect 522414 734 526110 856
rect 526278 734 529974 856
rect 530142 734 533838 856
rect 534006 734 537702 856
rect 537870 734 541566 856
rect 541734 734 545430 856
rect 545598 734 549938 856
rect 550106 734 553802 856
rect 553970 734 557666 856
rect 557834 734 561530 856
rect 561698 734 565394 856
rect 565562 734 569258 856
rect 569426 734 573122 856
rect 573290 734 576986 856
rect 577154 734 580850 856
rect 581018 734 582658 856
<< metal3 >>
rect 583200 701768 583800 701888
rect 200 700408 800 700528
rect 583200 697688 583800 697808
rect 200 696328 800 696448
rect 583200 693608 583800 693728
rect 200 692248 800 692368
rect 583200 689528 583800 689648
rect 200 688168 800 688288
rect 583200 685448 583800 685568
rect 200 684088 800 684208
rect 583200 681368 583800 681488
rect 200 680008 800 680128
rect 583200 677288 583800 677408
rect 200 675928 800 676048
rect 583200 673208 583800 673328
rect 200 671848 800 671968
rect 583200 669128 583800 669248
rect 200 667768 800 667888
rect 583200 665048 583800 665168
rect 200 663688 800 663808
rect 583200 660288 583800 660408
rect 200 658928 800 659048
rect 583200 656208 583800 656328
rect 200 654848 800 654968
rect 583200 652128 583800 652248
rect 200 650768 800 650888
rect 583200 648048 583800 648168
rect 200 646688 800 646808
rect 583200 643968 583800 644088
rect 200 642608 800 642728
rect 583200 639888 583800 640008
rect 200 638528 800 638648
rect 583200 635808 583800 635928
rect 200 634448 800 634568
rect 583200 631728 583800 631848
rect 200 630368 800 630488
rect 583200 627648 583800 627768
rect 200 626288 800 626408
rect 583200 623568 583800 623688
rect 200 622208 800 622328
rect 583200 618808 583800 618928
rect 200 617448 800 617568
rect 583200 614728 583800 614848
rect 200 613368 800 613488
rect 583200 610648 583800 610768
rect 200 609288 800 609408
rect 583200 606568 583800 606688
rect 200 605208 800 605328
rect 583200 602488 583800 602608
rect 200 601128 800 601248
rect 583200 598408 583800 598528
rect 200 597048 800 597168
rect 583200 594328 583800 594448
rect 200 592968 800 593088
rect 583200 590248 583800 590368
rect 200 588888 800 589008
rect 583200 586168 583800 586288
rect 200 584808 800 584928
rect 583200 582088 583800 582208
rect 200 580728 800 580848
rect 583200 577328 583800 577448
rect 200 575968 800 576088
rect 583200 573248 583800 573368
rect 200 571888 800 572008
rect 583200 569168 583800 569288
rect 200 567808 800 567928
rect 583200 565088 583800 565208
rect 200 563728 800 563848
rect 583200 561008 583800 561128
rect 200 559648 800 559768
rect 583200 556928 583800 557048
rect 200 555568 800 555688
rect 583200 552848 583800 552968
rect 200 551488 800 551608
rect 583200 548768 583800 548888
rect 200 547408 800 547528
rect 583200 544688 583800 544808
rect 200 543328 800 543448
rect 583200 540608 583800 540728
rect 200 539248 800 539368
rect 583200 535848 583800 535968
rect 200 534488 800 534608
rect 583200 531768 583800 531888
rect 200 530408 800 530528
rect 583200 527688 583800 527808
rect 200 526328 800 526448
rect 583200 523608 583800 523728
rect 200 522248 800 522368
rect 583200 519528 583800 519648
rect 200 518168 800 518288
rect 583200 515448 583800 515568
rect 200 514088 800 514208
rect 583200 511368 583800 511488
rect 200 510008 800 510128
rect 583200 507288 583800 507408
rect 200 505928 800 506048
rect 583200 503208 583800 503328
rect 200 501848 800 501968
rect 583200 499128 583800 499248
rect 200 497768 800 497888
rect 583200 494368 583800 494488
rect 200 493008 800 493128
rect 583200 490288 583800 490408
rect 200 488928 800 489048
rect 583200 486208 583800 486328
rect 200 484848 800 484968
rect 583200 482128 583800 482248
rect 200 480768 800 480888
rect 583200 478048 583800 478168
rect 200 476688 800 476808
rect 583200 473968 583800 474088
rect 200 472608 800 472728
rect 583200 469888 583800 470008
rect 200 468528 800 468648
rect 583200 465808 583800 465928
rect 200 464448 800 464568
rect 583200 461728 583800 461848
rect 200 460368 800 460488
rect 583200 457648 583800 457768
rect 200 456288 800 456408
rect 583200 452888 583800 453008
rect 200 451528 800 451648
rect 583200 448808 583800 448928
rect 200 447448 800 447568
rect 583200 444728 583800 444848
rect 200 443368 800 443488
rect 583200 440648 583800 440768
rect 200 439288 800 439408
rect 583200 436568 583800 436688
rect 200 435208 800 435328
rect 583200 432488 583800 432608
rect 200 431128 800 431248
rect 583200 428408 583800 428528
rect 200 427048 800 427168
rect 583200 424328 583800 424448
rect 200 422968 800 423088
rect 583200 420248 583800 420368
rect 200 418888 800 419008
rect 583200 416168 583800 416288
rect 200 414808 800 414928
rect 583200 411408 583800 411528
rect 200 410048 800 410168
rect 583200 407328 583800 407448
rect 200 405968 800 406088
rect 583200 403248 583800 403368
rect 200 401888 800 402008
rect 583200 399168 583800 399288
rect 200 397808 800 397928
rect 583200 395088 583800 395208
rect 200 393728 800 393848
rect 583200 391008 583800 391128
rect 200 389648 800 389768
rect 583200 386928 583800 387048
rect 200 385568 800 385688
rect 583200 382848 583800 382968
rect 200 381488 800 381608
rect 583200 378768 583800 378888
rect 200 377408 800 377528
rect 583200 374688 583800 374808
rect 200 373328 800 373448
rect 583200 369928 583800 370048
rect 200 368568 800 368688
rect 583200 365848 583800 365968
rect 200 364488 800 364608
rect 583200 361768 583800 361888
rect 200 360408 800 360528
rect 583200 357688 583800 357808
rect 200 356328 800 356448
rect 583200 353608 583800 353728
rect 200 352248 800 352368
rect 583200 349528 583800 349648
rect 200 348168 800 348288
rect 583200 345448 583800 345568
rect 200 344088 800 344208
rect 583200 341368 583800 341488
rect 200 340008 800 340128
rect 583200 337288 583800 337408
rect 200 335928 800 336048
rect 583200 333208 583800 333328
rect 200 331848 800 331968
rect 583200 328448 583800 328568
rect 200 327088 800 327208
rect 583200 324368 583800 324488
rect 200 323008 800 323128
rect 583200 320288 583800 320408
rect 200 318928 800 319048
rect 583200 316208 583800 316328
rect 200 314848 800 314968
rect 583200 312128 583800 312248
rect 200 310768 800 310888
rect 583200 308048 583800 308168
rect 200 306688 800 306808
rect 583200 303968 583800 304088
rect 200 302608 800 302728
rect 583200 299888 583800 300008
rect 200 298528 800 298648
rect 583200 295808 583800 295928
rect 200 294448 800 294568
rect 583200 291728 583800 291848
rect 200 290368 800 290488
rect 583200 286968 583800 287088
rect 200 285608 800 285728
rect 583200 282888 583800 283008
rect 200 281528 800 281648
rect 583200 278808 583800 278928
rect 200 277448 800 277568
rect 583200 274728 583800 274848
rect 200 273368 800 273488
rect 583200 270648 583800 270768
rect 200 269288 800 269408
rect 583200 266568 583800 266688
rect 200 265208 800 265328
rect 583200 262488 583800 262608
rect 200 261128 800 261248
rect 583200 258408 583800 258528
rect 200 257048 800 257168
rect 583200 254328 583800 254448
rect 200 252968 800 253088
rect 583200 249568 583800 249688
rect 200 248888 800 249008
rect 583200 245488 583800 245608
rect 200 244128 800 244248
rect 583200 241408 583800 241528
rect 200 240048 800 240168
rect 583200 237328 583800 237448
rect 200 235968 800 236088
rect 583200 233248 583800 233368
rect 200 231888 800 232008
rect 583200 229168 583800 229288
rect 200 227808 800 227928
rect 583200 225088 583800 225208
rect 200 223728 800 223848
rect 583200 221008 583800 221128
rect 200 219648 800 219768
rect 583200 216928 583800 217048
rect 200 215568 800 215688
rect 583200 212848 583800 212968
rect 200 211488 800 211608
rect 583200 208088 583800 208208
rect 200 207408 800 207528
rect 583200 204008 583800 204128
rect 200 202648 800 202768
rect 583200 199928 583800 200048
rect 200 198568 800 198688
rect 583200 195848 583800 195968
rect 200 194488 800 194608
rect 583200 191768 583800 191888
rect 200 190408 800 190528
rect 583200 187688 583800 187808
rect 200 186328 800 186448
rect 583200 183608 583800 183728
rect 200 182248 800 182368
rect 583200 179528 583800 179648
rect 200 178168 800 178288
rect 583200 175448 583800 175568
rect 200 174088 800 174208
rect 583200 171368 583800 171488
rect 200 170008 800 170128
rect 583200 166608 583800 166728
rect 200 165928 800 166048
rect 583200 162528 583800 162648
rect 200 161168 800 161288
rect 583200 158448 583800 158568
rect 200 157088 800 157208
rect 583200 154368 583800 154488
rect 200 153008 800 153128
rect 583200 150288 583800 150408
rect 200 148928 800 149048
rect 583200 146208 583800 146328
rect 200 144848 800 144968
rect 583200 142128 583800 142248
rect 200 140768 800 140888
rect 583200 138048 583800 138168
rect 200 136688 800 136808
rect 583200 133968 583800 134088
rect 200 132608 800 132728
rect 583200 129888 583800 130008
rect 200 128528 800 128648
rect 583200 125128 583800 125248
rect 200 124448 800 124568
rect 583200 121048 583800 121168
rect 200 119688 800 119808
rect 583200 116968 583800 117088
rect 200 115608 800 115728
rect 583200 112888 583800 113008
rect 200 111528 800 111648
rect 583200 108808 583800 108928
rect 200 107448 800 107568
rect 583200 104728 583800 104848
rect 200 103368 800 103488
rect 583200 100648 583800 100768
rect 200 99288 800 99408
rect 583200 96568 583800 96688
rect 200 95208 800 95328
rect 583200 92488 583800 92608
rect 200 91128 800 91248
rect 583200 88408 583800 88528
rect 200 87048 800 87168
rect 583200 83648 583800 83768
rect 200 82968 800 83088
rect 583200 79568 583800 79688
rect 200 78208 800 78328
rect 583200 75488 583800 75608
rect 200 74128 800 74248
rect 583200 71408 583800 71528
rect 200 70048 800 70168
rect 583200 67328 583800 67448
rect 200 65968 800 66088
rect 583200 63248 583800 63368
rect 200 61888 800 62008
rect 583200 59168 583800 59288
rect 200 57808 800 57928
rect 583200 55088 583800 55208
rect 200 53728 800 53848
rect 583200 51008 583800 51128
rect 200 49648 800 49768
rect 583200 46928 583800 47048
rect 200 45568 800 45688
rect 583200 42168 583800 42288
rect 200 41488 800 41608
rect 583200 38088 583800 38208
rect 200 36728 800 36848
rect 583200 34008 583800 34128
rect 200 32648 800 32768
rect 583200 29928 583800 30048
rect 200 28568 800 28688
rect 583200 25848 583800 25968
rect 200 24488 800 24608
rect 583200 21768 583800 21888
rect 200 20408 800 20528
rect 583200 17688 583800 17808
rect 200 16328 800 16448
rect 583200 13608 583800 13728
rect 200 12248 800 12368
rect 583200 9528 583800 9648
rect 200 8168 800 8288
rect 583200 5448 583800 5568
rect 200 4088 800 4208
rect 583200 688 583800 808
<< obsm3 >>
rect 800 701688 583120 701793
rect 800 700608 583200 701688
rect 880 700328 583200 700608
rect 800 697888 583200 700328
rect 800 697608 583120 697888
rect 800 696528 583200 697608
rect 880 696248 583200 696528
rect 800 693808 583200 696248
rect 800 693528 583120 693808
rect 800 692448 583200 693528
rect 880 692168 583200 692448
rect 800 689728 583200 692168
rect 800 689448 583120 689728
rect 800 688368 583200 689448
rect 880 688088 583200 688368
rect 800 685648 583200 688088
rect 800 685368 583120 685648
rect 800 684288 583200 685368
rect 880 684008 583200 684288
rect 800 681568 583200 684008
rect 800 681288 583120 681568
rect 800 680208 583200 681288
rect 880 679928 583200 680208
rect 800 677488 583200 679928
rect 800 677208 583120 677488
rect 800 676128 583200 677208
rect 880 675848 583200 676128
rect 800 673408 583200 675848
rect 800 673128 583120 673408
rect 800 672048 583200 673128
rect 880 671768 583200 672048
rect 800 669328 583200 671768
rect 800 669048 583120 669328
rect 800 667968 583200 669048
rect 880 667688 583200 667968
rect 800 665248 583200 667688
rect 800 664968 583120 665248
rect 800 663888 583200 664968
rect 880 663608 583200 663888
rect 800 660488 583200 663608
rect 800 660208 583120 660488
rect 800 659128 583200 660208
rect 880 658848 583200 659128
rect 800 656408 583200 658848
rect 800 656128 583120 656408
rect 800 655048 583200 656128
rect 880 654768 583200 655048
rect 800 652328 583200 654768
rect 800 652048 583120 652328
rect 800 650968 583200 652048
rect 880 650688 583200 650968
rect 800 648248 583200 650688
rect 800 647968 583120 648248
rect 800 646888 583200 647968
rect 880 646608 583200 646888
rect 800 644168 583200 646608
rect 800 643888 583120 644168
rect 800 642808 583200 643888
rect 880 642528 583200 642808
rect 800 640088 583200 642528
rect 800 639808 583120 640088
rect 800 638728 583200 639808
rect 880 638448 583200 638728
rect 800 636008 583200 638448
rect 800 635728 583120 636008
rect 800 634648 583200 635728
rect 880 634368 583200 634648
rect 800 631928 583200 634368
rect 800 631648 583120 631928
rect 800 630568 583200 631648
rect 880 630288 583200 630568
rect 800 627848 583200 630288
rect 800 627568 583120 627848
rect 800 626488 583200 627568
rect 880 626208 583200 626488
rect 800 623768 583200 626208
rect 800 623488 583120 623768
rect 800 622408 583200 623488
rect 880 622128 583200 622408
rect 800 619008 583200 622128
rect 800 618728 583120 619008
rect 800 617648 583200 618728
rect 880 617368 583200 617648
rect 800 614928 583200 617368
rect 800 614648 583120 614928
rect 800 613568 583200 614648
rect 880 613288 583200 613568
rect 800 610848 583200 613288
rect 800 610568 583120 610848
rect 800 609488 583200 610568
rect 880 609208 583200 609488
rect 800 606768 583200 609208
rect 800 606488 583120 606768
rect 800 605408 583200 606488
rect 880 605128 583200 605408
rect 800 602688 583200 605128
rect 800 602408 583120 602688
rect 800 601328 583200 602408
rect 880 601048 583200 601328
rect 800 598608 583200 601048
rect 800 598328 583120 598608
rect 800 597248 583200 598328
rect 880 596968 583200 597248
rect 800 594528 583200 596968
rect 800 594248 583120 594528
rect 800 593168 583200 594248
rect 880 592888 583200 593168
rect 800 590448 583200 592888
rect 800 590168 583120 590448
rect 800 589088 583200 590168
rect 880 588808 583200 589088
rect 800 586368 583200 588808
rect 800 586088 583120 586368
rect 800 585008 583200 586088
rect 880 584728 583200 585008
rect 800 582288 583200 584728
rect 800 582008 583120 582288
rect 800 580928 583200 582008
rect 880 580648 583200 580928
rect 800 577528 583200 580648
rect 800 577248 583120 577528
rect 800 576168 583200 577248
rect 880 575888 583200 576168
rect 800 573448 583200 575888
rect 800 573168 583120 573448
rect 800 572088 583200 573168
rect 880 571808 583200 572088
rect 800 569368 583200 571808
rect 800 569088 583120 569368
rect 800 568008 583200 569088
rect 880 567728 583200 568008
rect 800 565288 583200 567728
rect 800 565008 583120 565288
rect 800 563928 583200 565008
rect 880 563648 583200 563928
rect 800 561208 583200 563648
rect 800 560928 583120 561208
rect 800 559848 583200 560928
rect 880 559568 583200 559848
rect 800 557128 583200 559568
rect 800 556848 583120 557128
rect 800 555768 583200 556848
rect 880 555488 583200 555768
rect 800 553048 583200 555488
rect 800 552768 583120 553048
rect 800 551688 583200 552768
rect 880 551408 583200 551688
rect 800 548968 583200 551408
rect 800 548688 583120 548968
rect 800 547608 583200 548688
rect 880 547328 583200 547608
rect 800 544888 583200 547328
rect 800 544608 583120 544888
rect 800 543528 583200 544608
rect 880 543248 583200 543528
rect 800 540808 583200 543248
rect 800 540528 583120 540808
rect 800 539448 583200 540528
rect 880 539168 583200 539448
rect 800 536048 583200 539168
rect 800 535768 583120 536048
rect 800 534688 583200 535768
rect 880 534408 583200 534688
rect 800 531968 583200 534408
rect 800 531688 583120 531968
rect 800 530608 583200 531688
rect 880 530328 583200 530608
rect 800 527888 583200 530328
rect 800 527608 583120 527888
rect 800 526528 583200 527608
rect 880 526248 583200 526528
rect 800 523808 583200 526248
rect 800 523528 583120 523808
rect 800 522448 583200 523528
rect 880 522168 583200 522448
rect 800 519728 583200 522168
rect 800 519448 583120 519728
rect 800 518368 583200 519448
rect 880 518088 583200 518368
rect 800 515648 583200 518088
rect 800 515368 583120 515648
rect 800 514288 583200 515368
rect 880 514008 583200 514288
rect 800 511568 583200 514008
rect 800 511288 583120 511568
rect 800 510208 583200 511288
rect 880 509928 583200 510208
rect 800 507488 583200 509928
rect 800 507208 583120 507488
rect 800 506128 583200 507208
rect 880 505848 583200 506128
rect 800 503408 583200 505848
rect 800 503128 583120 503408
rect 800 502048 583200 503128
rect 880 501768 583200 502048
rect 800 499328 583200 501768
rect 800 499048 583120 499328
rect 800 497968 583200 499048
rect 880 497688 583200 497968
rect 800 494568 583200 497688
rect 800 494288 583120 494568
rect 800 493208 583200 494288
rect 880 492928 583200 493208
rect 800 490488 583200 492928
rect 800 490208 583120 490488
rect 800 489128 583200 490208
rect 880 488848 583200 489128
rect 800 486408 583200 488848
rect 800 486128 583120 486408
rect 800 485048 583200 486128
rect 880 484768 583200 485048
rect 800 482328 583200 484768
rect 800 482048 583120 482328
rect 800 480968 583200 482048
rect 880 480688 583200 480968
rect 800 478248 583200 480688
rect 800 477968 583120 478248
rect 800 476888 583200 477968
rect 880 476608 583200 476888
rect 800 474168 583200 476608
rect 800 473888 583120 474168
rect 800 472808 583200 473888
rect 880 472528 583200 472808
rect 800 470088 583200 472528
rect 800 469808 583120 470088
rect 800 468728 583200 469808
rect 880 468448 583200 468728
rect 800 466008 583200 468448
rect 800 465728 583120 466008
rect 800 464648 583200 465728
rect 880 464368 583200 464648
rect 800 461928 583200 464368
rect 800 461648 583120 461928
rect 800 460568 583200 461648
rect 880 460288 583200 460568
rect 800 457848 583200 460288
rect 800 457568 583120 457848
rect 800 456488 583200 457568
rect 880 456208 583200 456488
rect 800 453088 583200 456208
rect 800 452808 583120 453088
rect 800 451728 583200 452808
rect 880 451448 583200 451728
rect 800 449008 583200 451448
rect 800 448728 583120 449008
rect 800 447648 583200 448728
rect 880 447368 583200 447648
rect 800 444928 583200 447368
rect 800 444648 583120 444928
rect 800 443568 583200 444648
rect 880 443288 583200 443568
rect 800 440848 583200 443288
rect 800 440568 583120 440848
rect 800 439488 583200 440568
rect 880 439208 583200 439488
rect 800 436768 583200 439208
rect 800 436488 583120 436768
rect 800 435408 583200 436488
rect 880 435128 583200 435408
rect 800 432688 583200 435128
rect 800 432408 583120 432688
rect 800 431328 583200 432408
rect 880 431048 583200 431328
rect 800 428608 583200 431048
rect 800 428328 583120 428608
rect 800 427248 583200 428328
rect 880 426968 583200 427248
rect 800 424528 583200 426968
rect 800 424248 583120 424528
rect 800 423168 583200 424248
rect 880 422888 583200 423168
rect 800 420448 583200 422888
rect 800 420168 583120 420448
rect 800 419088 583200 420168
rect 880 418808 583200 419088
rect 800 416368 583200 418808
rect 800 416088 583120 416368
rect 800 415008 583200 416088
rect 880 414728 583200 415008
rect 800 411608 583200 414728
rect 800 411328 583120 411608
rect 800 410248 583200 411328
rect 880 409968 583200 410248
rect 800 407528 583200 409968
rect 800 407248 583120 407528
rect 800 406168 583200 407248
rect 880 405888 583200 406168
rect 800 403448 583200 405888
rect 800 403168 583120 403448
rect 800 402088 583200 403168
rect 880 401808 583200 402088
rect 800 399368 583200 401808
rect 800 399088 583120 399368
rect 800 398008 583200 399088
rect 880 397728 583200 398008
rect 800 395288 583200 397728
rect 800 395008 583120 395288
rect 800 393928 583200 395008
rect 880 393648 583200 393928
rect 800 391208 583200 393648
rect 800 390928 583120 391208
rect 800 389848 583200 390928
rect 880 389568 583200 389848
rect 800 387128 583200 389568
rect 800 386848 583120 387128
rect 800 385768 583200 386848
rect 880 385488 583200 385768
rect 800 383048 583200 385488
rect 800 382768 583120 383048
rect 800 381688 583200 382768
rect 880 381408 583200 381688
rect 800 378968 583200 381408
rect 800 378688 583120 378968
rect 800 377608 583200 378688
rect 880 377328 583200 377608
rect 800 374888 583200 377328
rect 800 374608 583120 374888
rect 800 373528 583200 374608
rect 880 373248 583200 373528
rect 800 370128 583200 373248
rect 800 369848 583120 370128
rect 800 368768 583200 369848
rect 880 368488 583200 368768
rect 800 366048 583200 368488
rect 800 365768 583120 366048
rect 800 364688 583200 365768
rect 880 364408 583200 364688
rect 800 361968 583200 364408
rect 800 361688 583120 361968
rect 800 360608 583200 361688
rect 880 360328 583200 360608
rect 800 357888 583200 360328
rect 800 357608 583120 357888
rect 800 356528 583200 357608
rect 880 356248 583200 356528
rect 800 353808 583200 356248
rect 800 353528 583120 353808
rect 800 352448 583200 353528
rect 880 352168 583200 352448
rect 800 349728 583200 352168
rect 800 349448 583120 349728
rect 800 348368 583200 349448
rect 880 348088 583200 348368
rect 800 345648 583200 348088
rect 800 345368 583120 345648
rect 800 344288 583200 345368
rect 880 344008 583200 344288
rect 800 341568 583200 344008
rect 800 341288 583120 341568
rect 800 340208 583200 341288
rect 880 339928 583200 340208
rect 800 337488 583200 339928
rect 800 337208 583120 337488
rect 800 336128 583200 337208
rect 880 335848 583200 336128
rect 800 333408 583200 335848
rect 800 333128 583120 333408
rect 800 332048 583200 333128
rect 880 331768 583200 332048
rect 800 328648 583200 331768
rect 800 328368 583120 328648
rect 800 327288 583200 328368
rect 880 327008 583200 327288
rect 800 324568 583200 327008
rect 800 324288 583120 324568
rect 800 323208 583200 324288
rect 880 322928 583200 323208
rect 800 320488 583200 322928
rect 800 320208 583120 320488
rect 800 319128 583200 320208
rect 880 318848 583200 319128
rect 800 316408 583200 318848
rect 800 316128 583120 316408
rect 800 315048 583200 316128
rect 880 314768 583200 315048
rect 800 312328 583200 314768
rect 800 312048 583120 312328
rect 800 310968 583200 312048
rect 880 310688 583200 310968
rect 800 308248 583200 310688
rect 800 307968 583120 308248
rect 800 306888 583200 307968
rect 880 306608 583200 306888
rect 800 304168 583200 306608
rect 800 303888 583120 304168
rect 800 302808 583200 303888
rect 880 302528 583200 302808
rect 800 300088 583200 302528
rect 800 299808 583120 300088
rect 800 298728 583200 299808
rect 880 298448 583200 298728
rect 800 296008 583200 298448
rect 800 295728 583120 296008
rect 800 294648 583200 295728
rect 880 294368 583200 294648
rect 800 291928 583200 294368
rect 800 291648 583120 291928
rect 800 290568 583200 291648
rect 880 290288 583200 290568
rect 800 287168 583200 290288
rect 800 286888 583120 287168
rect 800 285808 583200 286888
rect 880 285528 583200 285808
rect 800 283088 583200 285528
rect 800 282808 583120 283088
rect 800 281728 583200 282808
rect 880 281448 583200 281728
rect 800 279008 583200 281448
rect 800 278728 583120 279008
rect 800 277648 583200 278728
rect 880 277368 583200 277648
rect 800 274928 583200 277368
rect 800 274648 583120 274928
rect 800 273568 583200 274648
rect 880 273288 583200 273568
rect 800 270848 583200 273288
rect 800 270568 583120 270848
rect 800 269488 583200 270568
rect 880 269208 583200 269488
rect 800 266768 583200 269208
rect 800 266488 583120 266768
rect 800 265408 583200 266488
rect 880 265128 583200 265408
rect 800 262688 583200 265128
rect 800 262408 583120 262688
rect 800 261328 583200 262408
rect 880 261048 583200 261328
rect 800 258608 583200 261048
rect 800 258328 583120 258608
rect 800 257248 583200 258328
rect 880 256968 583200 257248
rect 800 254528 583200 256968
rect 800 254248 583120 254528
rect 800 253168 583200 254248
rect 880 252888 583200 253168
rect 800 249768 583200 252888
rect 800 249488 583120 249768
rect 800 249088 583200 249488
rect 880 248808 583200 249088
rect 800 245688 583200 248808
rect 800 245408 583120 245688
rect 800 244328 583200 245408
rect 880 244048 583200 244328
rect 800 241608 583200 244048
rect 800 241328 583120 241608
rect 800 240248 583200 241328
rect 880 239968 583200 240248
rect 800 237528 583200 239968
rect 800 237248 583120 237528
rect 800 236168 583200 237248
rect 880 235888 583200 236168
rect 800 233448 583200 235888
rect 800 233168 583120 233448
rect 800 232088 583200 233168
rect 880 231808 583200 232088
rect 800 229368 583200 231808
rect 800 229088 583120 229368
rect 800 228008 583200 229088
rect 880 227728 583200 228008
rect 800 225288 583200 227728
rect 800 225008 583120 225288
rect 800 223928 583200 225008
rect 880 223648 583200 223928
rect 800 221208 583200 223648
rect 800 220928 583120 221208
rect 800 219848 583200 220928
rect 880 219568 583200 219848
rect 800 217128 583200 219568
rect 800 216848 583120 217128
rect 800 215768 583200 216848
rect 880 215488 583200 215768
rect 800 213048 583200 215488
rect 800 212768 583120 213048
rect 800 211688 583200 212768
rect 880 211408 583200 211688
rect 800 208288 583200 211408
rect 800 208008 583120 208288
rect 800 207608 583200 208008
rect 880 207328 583200 207608
rect 800 204208 583200 207328
rect 800 203928 583120 204208
rect 800 202848 583200 203928
rect 880 202568 583200 202848
rect 800 200128 583200 202568
rect 800 199848 583120 200128
rect 800 198768 583200 199848
rect 880 198488 583200 198768
rect 800 196048 583200 198488
rect 800 195768 583120 196048
rect 800 194688 583200 195768
rect 880 194408 583200 194688
rect 800 191968 583200 194408
rect 800 191688 583120 191968
rect 800 190608 583200 191688
rect 880 190328 583200 190608
rect 800 187888 583200 190328
rect 800 187608 583120 187888
rect 800 186528 583200 187608
rect 880 186248 583200 186528
rect 800 183808 583200 186248
rect 800 183528 583120 183808
rect 800 182448 583200 183528
rect 880 182168 583200 182448
rect 800 179728 583200 182168
rect 800 179448 583120 179728
rect 800 178368 583200 179448
rect 880 178088 583200 178368
rect 800 175648 583200 178088
rect 800 175368 583120 175648
rect 800 174288 583200 175368
rect 880 174008 583200 174288
rect 800 171568 583200 174008
rect 800 171288 583120 171568
rect 800 170208 583200 171288
rect 880 169928 583200 170208
rect 800 166808 583200 169928
rect 800 166528 583120 166808
rect 800 166128 583200 166528
rect 880 165848 583200 166128
rect 800 162728 583200 165848
rect 800 162448 583120 162728
rect 800 161368 583200 162448
rect 880 161088 583200 161368
rect 800 158648 583200 161088
rect 800 158368 583120 158648
rect 800 157288 583200 158368
rect 880 157008 583200 157288
rect 800 154568 583200 157008
rect 800 154288 583120 154568
rect 800 153208 583200 154288
rect 880 152928 583200 153208
rect 800 150488 583200 152928
rect 800 150208 583120 150488
rect 800 149128 583200 150208
rect 880 148848 583200 149128
rect 800 146408 583200 148848
rect 800 146128 583120 146408
rect 800 145048 583200 146128
rect 880 144768 583200 145048
rect 800 142328 583200 144768
rect 800 142048 583120 142328
rect 800 140968 583200 142048
rect 880 140688 583200 140968
rect 800 138248 583200 140688
rect 800 137968 583120 138248
rect 800 136888 583200 137968
rect 880 136608 583200 136888
rect 800 134168 583200 136608
rect 800 133888 583120 134168
rect 800 132808 583200 133888
rect 880 132528 583200 132808
rect 800 130088 583200 132528
rect 800 129808 583120 130088
rect 800 128728 583200 129808
rect 880 128448 583200 128728
rect 800 125328 583200 128448
rect 800 125048 583120 125328
rect 800 124648 583200 125048
rect 880 124368 583200 124648
rect 800 121248 583200 124368
rect 800 120968 583120 121248
rect 800 119888 583200 120968
rect 880 119608 583200 119888
rect 800 117168 583200 119608
rect 800 116888 583120 117168
rect 800 115808 583200 116888
rect 880 115528 583200 115808
rect 800 113088 583200 115528
rect 800 112808 583120 113088
rect 800 111728 583200 112808
rect 880 111448 583200 111728
rect 800 109008 583200 111448
rect 800 108728 583120 109008
rect 800 107648 583200 108728
rect 880 107368 583200 107648
rect 800 104928 583200 107368
rect 800 104648 583120 104928
rect 800 103568 583200 104648
rect 880 103288 583200 103568
rect 800 100848 583200 103288
rect 800 100568 583120 100848
rect 800 99488 583200 100568
rect 880 99208 583200 99488
rect 800 96768 583200 99208
rect 800 96488 583120 96768
rect 800 95408 583200 96488
rect 880 95128 583200 95408
rect 800 92688 583200 95128
rect 800 92408 583120 92688
rect 800 91328 583200 92408
rect 880 91048 583200 91328
rect 800 88608 583200 91048
rect 800 88328 583120 88608
rect 800 87248 583200 88328
rect 880 86968 583200 87248
rect 800 83848 583200 86968
rect 800 83568 583120 83848
rect 800 83168 583200 83568
rect 880 82888 583200 83168
rect 800 79768 583200 82888
rect 800 79488 583120 79768
rect 800 78408 583200 79488
rect 880 78128 583200 78408
rect 800 75688 583200 78128
rect 800 75408 583120 75688
rect 800 74328 583200 75408
rect 880 74048 583200 74328
rect 800 71608 583200 74048
rect 800 71328 583120 71608
rect 800 70248 583200 71328
rect 880 69968 583200 70248
rect 800 67528 583200 69968
rect 800 67248 583120 67528
rect 800 66168 583200 67248
rect 880 65888 583200 66168
rect 800 63448 583200 65888
rect 800 63168 583120 63448
rect 800 62088 583200 63168
rect 880 61808 583200 62088
rect 800 59368 583200 61808
rect 800 59088 583120 59368
rect 800 58008 583200 59088
rect 880 57728 583200 58008
rect 800 55288 583200 57728
rect 800 55008 583120 55288
rect 800 53928 583200 55008
rect 880 53648 583200 53928
rect 800 51208 583200 53648
rect 800 50928 583120 51208
rect 800 49848 583200 50928
rect 880 49568 583200 49848
rect 800 47128 583200 49568
rect 800 46848 583120 47128
rect 800 45768 583200 46848
rect 880 45488 583200 45768
rect 800 42368 583200 45488
rect 800 42088 583120 42368
rect 800 41688 583200 42088
rect 880 41408 583200 41688
rect 800 38288 583200 41408
rect 800 38008 583120 38288
rect 800 36928 583200 38008
rect 880 36648 583200 36928
rect 800 34208 583200 36648
rect 800 33928 583120 34208
rect 800 32848 583200 33928
rect 880 32568 583200 32848
rect 800 30128 583200 32568
rect 800 29848 583120 30128
rect 800 28768 583200 29848
rect 880 28488 583200 28768
rect 800 26048 583200 28488
rect 800 25768 583120 26048
rect 800 24688 583200 25768
rect 880 24408 583200 24688
rect 800 21968 583200 24408
rect 800 21688 583120 21968
rect 800 20608 583200 21688
rect 880 20328 583200 20608
rect 800 17888 583200 20328
rect 800 17608 583120 17888
rect 800 16528 583200 17608
rect 880 16248 583200 16528
rect 800 13808 583200 16248
rect 800 13528 583120 13808
rect 800 12448 583200 13528
rect 880 12168 583200 12448
rect 800 9728 583200 12168
rect 800 9448 583120 9728
rect 800 8368 583200 9448
rect 880 8088 583200 8368
rect 800 5648 583200 8088
rect 800 5368 583120 5648
rect 800 4288 583200 5368
rect 880 4008 583200 4288
rect 800 2143 583200 4008
<< metal4 >>
rect -5036 -3964 -4716 707900
rect -4376 -3304 -4056 707240
rect -3716 -2644 -3396 706580
rect -3056 -1984 -2736 705920
rect -2396 -1324 -2076 705260
rect -1736 -664 -1416 704600
rect -1076 -4 -756 703940
rect -416 656 -96 703280
rect 4900 54352 5220 649584
rect 8344 -3964 8664 707900
rect 9004 -3964 9324 707900
rect 9664 -3964 9984 707900
rect 10324 -3964 10644 707900
rect 10984 -3964 11304 707900
rect 11644 -3964 11964 707900
rect 12304 -3964 12624 707900
rect 12964 -3964 13284 707900
rect 22344 646209 22664 707900
rect 23004 646209 23324 707900
rect 23664 646209 23984 707900
rect 24324 646209 24644 707900
rect 24984 646209 25304 707900
rect 25644 646209 25964 707900
rect 26304 646209 26624 707900
rect 26964 646209 27284 707900
rect 36344 646209 36664 707900
rect 37004 646209 37324 707900
rect 37664 646209 37984 707900
rect 38324 646209 38644 707900
rect 38984 646209 39304 707900
rect 39644 646209 39964 707900
rect 40304 646209 40624 707900
rect 40964 646209 41284 707900
rect 50344 646209 50664 707900
rect 51004 646209 51324 707900
rect 51664 646209 51984 707900
rect 52324 646209 52644 707900
rect 52984 646209 53304 707900
rect 53644 646209 53964 707900
rect 54304 646209 54624 707900
rect 54964 646209 55284 707900
rect 64344 646209 64664 707900
rect 65004 646209 65324 707900
rect 65664 646209 65984 707900
rect 66324 646209 66644 707900
rect 66984 646209 67304 707900
rect 67644 646209 67964 707900
rect 68304 646209 68624 707900
rect 68964 646209 69284 707900
rect 78344 646209 78664 707900
rect 79004 646209 79324 707900
rect 79664 646209 79984 707900
rect 80324 646209 80644 707900
rect 80984 646209 81304 707900
rect 81644 646209 81964 707900
rect 82304 646209 82624 707900
rect 82964 646209 83284 707900
rect 92344 646209 92664 707900
rect 93004 646209 93324 707900
rect 93664 646209 93984 707900
rect 94324 646209 94644 707900
rect 94984 646209 95304 707900
rect 95644 646209 95964 707900
rect 96304 646209 96624 707900
rect 96964 646209 97284 707900
rect 106344 646209 106664 707900
rect 107004 646209 107324 707900
rect 107664 646209 107984 707900
rect 108324 646209 108644 707900
rect 108984 646209 109304 707900
rect 109644 646209 109964 707900
rect 110304 646209 110624 707900
rect 110964 646209 111284 707900
rect 120344 646209 120664 707900
rect 121004 646209 121324 707900
rect 121664 646209 121984 707900
rect 122324 646209 122644 707900
rect 122984 646209 123304 707900
rect 123644 646209 123964 707900
rect 124304 646209 124624 707900
rect 124964 646209 125284 707900
rect 134344 646209 134664 707900
rect 135004 646209 135324 707900
rect 135664 646209 135984 707900
rect 136324 646209 136644 707900
rect 136984 646209 137304 707900
rect 137644 646209 137964 707900
rect 138304 646209 138624 707900
rect 138964 646209 139284 707900
rect 148344 646209 148664 707900
rect 149004 646209 149324 707900
rect 149664 646209 149984 707900
rect 150324 646209 150644 707900
rect 150984 646209 151304 707900
rect 151644 646209 151964 707900
rect 152304 646209 152624 707900
rect 152964 646209 153284 707900
rect 162344 646209 162664 707900
rect 163004 646209 163324 707900
rect 163664 646209 163984 707900
rect 164324 646209 164644 707900
rect 164984 646209 165304 707900
rect 165644 646209 165964 707900
rect 166304 646209 166624 707900
rect 166964 646209 167284 707900
rect 176344 646209 176664 707900
rect 177004 646209 177324 707900
rect 177664 646209 177984 707900
rect 178324 646209 178644 707900
rect 178984 646209 179304 707900
rect 179644 646209 179964 707900
rect 180304 646209 180624 707900
rect 180964 646209 181284 707900
rect 190344 646209 190664 707900
rect 191004 646209 191324 707900
rect 191664 646209 191984 707900
rect 192324 646209 192644 707900
rect 192984 646209 193304 707900
rect 193644 646209 193964 707900
rect 194304 646209 194624 707900
rect 194964 646209 195284 707900
rect 204344 646209 204664 707900
rect 205004 646209 205324 707900
rect 205664 646209 205984 707900
rect 206324 646209 206644 707900
rect 206984 646209 207304 707900
rect 207644 646209 207964 707900
rect 208304 646209 208624 707900
rect 208964 646209 209284 707900
rect 218344 646209 218664 707900
rect 219004 646209 219324 707900
rect 219664 646209 219984 707900
rect 220324 646209 220644 707900
rect 220984 646209 221304 707900
rect 221644 646209 221964 707900
rect 222304 646209 222624 707900
rect 222964 646209 223284 707900
rect 232344 646209 232664 707900
rect 233004 646209 233324 707900
rect 233664 646209 233984 707900
rect 234324 646209 234644 707900
rect 234984 646209 235304 707900
rect 235644 646209 235964 707900
rect 236304 646209 236624 707900
rect 236964 646209 237284 707900
rect 246344 646209 246664 707900
rect 247004 646209 247324 707900
rect 247664 646209 247984 707900
rect 248324 646209 248644 707900
rect 248984 646209 249304 707900
rect 249644 646209 249964 707900
rect 250304 646209 250624 707900
rect 250964 646209 251284 707900
rect 260344 646209 260664 707900
rect 261004 646209 261324 707900
rect 261664 646209 261984 707900
rect 262324 646209 262644 707900
rect 262984 646209 263304 707900
rect 263644 646209 263964 707900
rect 264304 646209 264624 707900
rect 264964 646209 265284 707900
rect 274344 646209 274664 707900
rect 275004 646209 275324 707900
rect 275664 646209 275984 707900
rect 276324 646209 276644 707900
rect 276984 646209 277304 707900
rect 277644 646209 277964 707900
rect 278304 646209 278624 707900
rect 278964 646209 279284 707900
rect 288344 646209 288664 707900
rect 289004 646209 289324 707900
rect 289664 646209 289984 707900
rect 290324 646209 290644 707900
rect 290984 646209 291304 707900
rect 291644 646209 291964 707900
rect 292304 646209 292624 707900
rect 292964 646209 293284 707900
rect 302344 646209 302664 707900
rect 303004 646209 303324 707900
rect 303664 646209 303984 707900
rect 304324 646209 304644 707900
rect 304984 646209 305304 707900
rect 305644 646209 305964 707900
rect 306304 646209 306624 707900
rect 306964 646209 307284 707900
rect 316344 646209 316664 707900
rect 317004 646209 317324 707900
rect 317664 646209 317984 707900
rect 318324 646209 318644 707900
rect 318984 646209 319304 707900
rect 319644 646209 319964 707900
rect 320304 646209 320624 707900
rect 320964 646209 321284 707900
rect 330344 646209 330664 707900
rect 331004 646209 331324 707900
rect 331664 646209 331984 707900
rect 332324 646209 332644 707900
rect 332984 646209 333304 707900
rect 333644 646209 333964 707900
rect 334304 646209 334624 707900
rect 334964 646209 335284 707900
rect 344344 646209 344664 707900
rect 345004 646209 345324 707900
rect 345664 646209 345984 707900
rect 346324 646209 346644 707900
rect 346984 646209 347304 707900
rect 347644 646209 347964 707900
rect 348304 646209 348624 707900
rect 348964 646209 349284 707900
rect 358344 646209 358664 707900
rect 359004 646209 359324 707900
rect 359664 646209 359984 707900
rect 360324 646209 360644 707900
rect 360984 646209 361304 707900
rect 361644 646209 361964 707900
rect 362304 646209 362624 707900
rect 362964 646209 363284 707900
rect 372344 646209 372664 707900
rect 373004 646209 373324 707900
rect 373664 646209 373984 707900
rect 374324 646209 374644 707900
rect 374984 646209 375304 707900
rect 375644 646209 375964 707900
rect 376304 646209 376624 707900
rect 376964 646209 377284 707900
rect 386344 646209 386664 707900
rect 387004 646209 387324 707900
rect 387664 646209 387984 707900
rect 388324 646209 388644 707900
rect 388984 646209 389304 707900
rect 389644 646209 389964 707900
rect 390304 646209 390624 707900
rect 390964 646209 391284 707900
rect 400344 646209 400664 707900
rect 401004 646209 401324 707900
rect 401664 646209 401984 707900
rect 402324 646209 402644 707900
rect 402984 646209 403304 707900
rect 403644 646209 403964 707900
rect 404304 646209 404624 707900
rect 404964 646209 405284 707900
rect 414344 646209 414664 707900
rect 415004 646209 415324 707900
rect 415664 646209 415984 707900
rect 416324 646209 416644 707900
rect 416984 646209 417304 707900
rect 417644 646209 417964 707900
rect 418304 646209 418624 707900
rect 418964 646209 419284 707900
rect 428344 646209 428664 707900
rect 429004 646209 429324 707900
rect 429664 646209 429984 707900
rect 430324 646209 430644 707900
rect 430984 646209 431304 707900
rect 431644 646209 431964 707900
rect 432304 646209 432624 707900
rect 432964 646209 433284 707900
rect 442344 646209 442664 707900
rect 443004 646209 443324 707900
rect 443664 646209 443984 707900
rect 444324 646209 444644 707900
rect 444984 646209 445304 707900
rect 445644 646209 445964 707900
rect 446304 646209 446624 707900
rect 446964 646209 447284 707900
rect 456344 646209 456664 707900
rect 457004 646209 457324 707900
rect 457664 646209 457984 707900
rect 458324 646209 458644 707900
rect 458984 646209 459304 707900
rect 459644 646209 459964 707900
rect 460304 646209 460624 707900
rect 460964 646209 461284 707900
rect 470344 646209 470664 707900
rect 471004 646209 471324 707900
rect 471664 646209 471984 707900
rect 472324 646209 472644 707900
rect 472984 646209 473304 707900
rect 473644 646209 473964 707900
rect 474304 646209 474624 707900
rect 474964 646209 475284 707900
rect 484344 646209 484664 707900
rect 485004 646209 485324 707900
rect 485664 646209 485984 707900
rect 486324 646209 486644 707900
rect 486984 646209 487304 707900
rect 487644 646209 487964 707900
rect 488304 646209 488624 707900
rect 488964 646209 489284 707900
rect 498344 646209 498664 707900
rect 499004 646209 499324 707900
rect 499664 646209 499984 707900
rect 500324 646209 500644 707900
rect 500984 646209 501304 707900
rect 501644 646209 501964 707900
rect 502304 646209 502624 707900
rect 502964 646209 503284 707900
rect 512344 646209 512664 707900
rect 513004 646209 513324 707900
rect 513664 646209 513984 707900
rect 514324 646209 514644 707900
rect 514984 646209 515304 707900
rect 515644 646209 515964 707900
rect 516304 646209 516624 707900
rect 516964 646209 517284 707900
rect 526344 646209 526664 707900
rect 527004 646209 527324 707900
rect 527664 646209 527984 707900
rect 528324 646209 528644 707900
rect 528984 646209 529304 707900
rect 529644 646209 529964 707900
rect 530304 646209 530624 707900
rect 530964 646209 531284 707900
rect 540344 646209 540664 707900
rect 541004 646209 541324 707900
rect 541664 646209 541984 707900
rect 542324 646209 542644 707900
rect 542984 646209 543304 707900
rect 543644 646209 543964 707900
rect 544304 646209 544624 707900
rect 544964 646209 545284 707900
rect 554344 646209 554664 707900
rect 555004 646209 555324 707900
rect 555664 646209 555984 707900
rect 556324 646209 556644 707900
rect 556984 646209 557304 707900
rect 557644 646209 557964 707900
rect 558304 646209 558624 707900
rect 558964 646209 559284 707900
rect 22344 -3964 22664 56679
rect 23004 -3964 23324 56679
rect 23664 -3964 23984 56679
rect 24324 -3964 24644 56679
rect 24984 -3964 25304 56679
rect 25644 -3964 25964 56679
rect 26304 -3964 26624 56679
rect 26964 -3964 27284 56679
rect 36344 -3964 36664 56679
rect 37004 -3964 37324 56679
rect 37664 -3964 37984 56679
rect 38324 -3964 38644 56679
rect 38984 -3964 39304 56679
rect 39644 -3964 39964 56679
rect 40304 -3964 40624 56679
rect 40964 -3964 41284 56679
rect 50344 -3964 50664 56679
rect 51004 -3964 51324 56679
rect 51664 -3964 51984 56679
rect 52324 -3964 52644 56679
rect 52984 -3964 53304 56679
rect 53644 -3964 53964 56679
rect 54304 -3964 54624 56679
rect 54964 -3964 55284 56679
rect 64344 -3964 64664 56679
rect 65004 -3964 65324 56679
rect 65664 -3964 65984 56679
rect 66324 -3964 66644 56679
rect 66984 -3964 67304 56679
rect 67644 -3964 67964 56679
rect 68304 -3964 68624 56679
rect 68964 -3964 69284 56679
rect 78344 -3964 78664 56679
rect 79004 -3964 79324 56679
rect 79664 -3964 79984 56679
rect 80324 -3964 80644 56679
rect 80984 -3964 81304 56679
rect 81644 -3964 81964 56679
rect 82304 -3964 82624 56679
rect 82964 -3964 83284 56679
rect 92344 -3964 92664 56679
rect 93004 -3964 93324 56679
rect 93664 -3964 93984 56679
rect 94324 -3964 94644 56679
rect 94984 -3964 95304 56679
rect 95644 -3964 95964 56679
rect 96304 -3964 96624 56679
rect 96964 -3964 97284 56679
rect 106344 -3964 106664 56679
rect 107004 -3964 107324 56679
rect 107664 -3964 107984 56679
rect 108324 -3964 108644 56679
rect 108984 -3964 109304 56679
rect 109644 -3964 109964 56679
rect 110304 -3964 110624 56679
rect 110964 -3964 111284 56679
rect 120344 -3964 120664 56679
rect 121004 -3964 121324 56679
rect 121664 -3964 121984 56679
rect 122324 -3964 122644 56679
rect 122984 -3964 123304 56679
rect 123644 -3964 123964 56679
rect 124304 -3964 124624 56679
rect 124964 -3964 125284 56679
rect 134344 -3964 134664 56679
rect 135004 -3964 135324 56679
rect 135664 -3964 135984 56679
rect 136324 -3964 136644 56679
rect 136984 -3964 137304 56679
rect 137644 -3964 137964 56679
rect 138304 -3964 138624 56679
rect 138964 -3964 139284 56679
rect 148344 -3964 148664 56679
rect 149004 -3964 149324 56679
rect 149664 -3964 149984 56679
rect 150324 -3964 150644 56679
rect 150984 -3964 151304 56679
rect 151644 -3964 151964 56679
rect 152304 -3964 152624 56679
rect 152964 -3964 153284 56679
rect 162344 -3964 162664 56679
rect 163004 -3964 163324 56679
rect 163664 -3964 163984 56679
rect 164324 -3964 164644 56679
rect 164984 -3964 165304 56679
rect 165644 -3964 165964 56679
rect 166304 -3964 166624 56679
rect 166964 -3964 167284 56679
rect 176344 -3964 176664 56679
rect 177004 -3964 177324 56679
rect 177664 -3964 177984 56679
rect 178324 -3964 178644 56679
rect 178984 -3964 179304 56679
rect 179644 -3964 179964 56679
rect 180304 -3964 180624 56679
rect 180964 -3964 181284 56679
rect 190344 -3964 190664 56679
rect 191004 -3964 191324 56679
rect 191664 -3964 191984 56679
rect 192324 -3964 192644 56679
rect 192984 -3964 193304 56679
rect 193644 -3964 193964 56679
rect 194304 -3964 194624 56679
rect 194964 -3964 195284 56679
rect 204344 -3964 204664 56679
rect 205004 -3964 205324 56679
rect 205664 -3964 205984 56679
rect 206324 -3964 206644 56679
rect 206984 -3964 207304 56679
rect 207644 -3964 207964 56679
rect 208304 -3964 208624 56679
rect 208964 -3964 209284 56679
rect 218344 -3964 218664 56679
rect 219004 -3964 219324 56679
rect 219664 -3964 219984 56679
rect 220324 -3964 220644 56679
rect 220984 -3964 221304 56679
rect 221644 -3964 221964 56679
rect 222304 -3964 222624 56679
rect 222964 -3964 223284 56679
rect 232344 -3964 232664 56679
rect 233004 -3964 233324 56679
rect 233664 -3964 233984 56679
rect 234324 -3964 234644 56679
rect 234984 -3964 235304 56679
rect 235644 -3964 235964 56679
rect 236304 -3964 236624 56679
rect 236964 -3964 237284 56679
rect 246344 -3964 246664 56679
rect 247004 -3964 247324 56679
rect 247664 -3964 247984 56679
rect 248324 -3964 248644 56679
rect 248984 -3964 249304 56679
rect 249644 -3964 249964 56679
rect 250304 -3964 250624 56679
rect 250964 -3964 251284 56679
rect 260344 -3964 260664 56679
rect 261004 -3964 261324 56679
rect 261664 -3964 261984 56679
rect 262324 -3964 262644 56679
rect 262984 -3964 263304 56679
rect 263644 -3964 263964 56679
rect 264304 -3964 264624 56679
rect 264964 -3964 265284 56679
rect 274344 -3964 274664 56679
rect 275004 -3964 275324 56679
rect 275664 -3964 275984 56679
rect 276324 -3964 276644 56679
rect 276984 -3964 277304 56679
rect 277644 -3964 277964 56679
rect 278304 -3964 278624 56679
rect 278964 -3964 279284 56679
rect 288344 -3964 288664 56679
rect 289004 -3964 289324 56679
rect 289664 -3964 289984 56679
rect 290324 -3964 290644 56679
rect 290984 -3964 291304 56679
rect 291644 -3964 291964 56679
rect 292304 -3964 292624 56679
rect 292964 -3964 293284 56679
rect 302344 -3964 302664 56679
rect 303004 -3964 303324 56679
rect 303664 -3964 303984 56679
rect 304324 -3964 304644 56679
rect 304984 -3964 305304 56679
rect 305644 -3964 305964 56679
rect 306304 -3964 306624 56679
rect 306964 -3964 307284 56679
rect 316344 -3964 316664 56679
rect 317004 -3964 317324 56679
rect 317664 -3964 317984 56679
rect 318324 -3964 318644 56679
rect 318984 -3964 319304 56679
rect 319644 -3964 319964 56679
rect 320304 -3964 320624 56679
rect 320964 -3964 321284 56679
rect 330344 -3964 330664 56679
rect 331004 -3964 331324 56679
rect 331664 -3964 331984 56679
rect 332324 -3964 332644 56679
rect 332984 -3964 333304 56679
rect 333644 -3964 333964 56679
rect 334304 -3964 334624 56679
rect 334964 -3964 335284 56679
rect 344344 -3964 344664 56679
rect 345004 -3964 345324 56679
rect 345664 -3964 345984 56679
rect 346324 -3964 346644 56679
rect 346984 -3964 347304 56679
rect 347644 -3964 347964 56679
rect 348304 -3964 348624 56679
rect 348964 -3964 349284 56679
rect 358344 -3964 358664 56679
rect 359004 -3964 359324 56679
rect 359664 -3964 359984 56679
rect 360324 -3964 360644 56679
rect 360984 -3964 361304 56679
rect 361644 -3964 361964 56679
rect 362304 -3964 362624 56679
rect 362964 -3964 363284 56679
rect 372344 -3964 372664 56679
rect 373004 -3964 373324 56679
rect 373664 -3964 373984 56679
rect 374324 -3964 374644 56679
rect 374984 -3964 375304 56679
rect 375644 -3964 375964 56679
rect 376304 -3964 376624 56679
rect 376964 -3964 377284 56679
rect 386344 -3964 386664 56679
rect 387004 -3964 387324 56679
rect 387664 -3964 387984 56679
rect 388324 -3964 388644 56679
rect 388984 -3964 389304 56679
rect 389644 -3964 389964 56679
rect 390304 -3964 390624 56679
rect 390964 -3964 391284 56679
rect 400344 -3964 400664 56679
rect 401004 -3964 401324 56679
rect 401664 -3964 401984 56679
rect 402324 -3964 402644 56679
rect 402984 -3964 403304 56679
rect 403644 -3964 403964 56679
rect 404304 -3964 404624 56679
rect 404964 -3964 405284 56679
rect 414344 -3964 414664 56679
rect 415004 -3964 415324 56679
rect 415664 -3964 415984 56679
rect 416324 -3964 416644 56679
rect 416984 -3964 417304 56679
rect 417644 -3964 417964 56679
rect 418304 -3964 418624 56679
rect 418964 -3964 419284 56679
rect 428344 -3964 428664 56679
rect 429004 -3964 429324 56679
rect 429664 -3964 429984 56679
rect 430324 -3964 430644 56679
rect 430984 -3964 431304 56679
rect 431644 -3964 431964 56679
rect 432304 -3964 432624 56679
rect 432964 -3964 433284 56679
rect 442344 -3964 442664 56679
rect 443004 -3964 443324 56679
rect 443664 -3964 443984 56679
rect 444324 -3964 444644 56679
rect 444984 -3964 445304 56679
rect 445644 -3964 445964 56679
rect 446304 -3964 446624 56679
rect 446964 -3964 447284 56679
rect 456344 -3964 456664 56679
rect 457004 -3964 457324 56679
rect 457664 -3964 457984 56679
rect 458324 -3964 458644 56679
rect 458984 -3964 459304 56679
rect 459644 -3964 459964 56679
rect 460304 -3964 460624 56679
rect 460964 -3964 461284 56679
rect 470344 -3964 470664 56679
rect 471004 -3964 471324 56679
rect 471664 -3964 471984 56679
rect 472324 -3964 472644 56679
rect 472984 -3964 473304 56679
rect 473644 -3964 473964 56679
rect 474304 -3964 474624 56679
rect 474964 -3964 475284 56679
rect 484344 -3964 484664 56679
rect 485004 -3964 485324 56679
rect 485664 -3964 485984 56679
rect 486324 -3964 486644 56679
rect 486984 -3964 487304 56679
rect 487644 -3964 487964 56679
rect 488304 -3964 488624 56679
rect 488964 -3964 489284 56679
rect 498344 -3964 498664 56679
rect 499004 -3964 499324 56679
rect 499664 -3964 499984 56679
rect 500324 -3964 500644 56679
rect 500984 -3964 501304 56679
rect 501644 -3964 501964 56679
rect 502304 -3964 502624 56679
rect 502964 -3964 503284 56679
rect 512344 -3964 512664 56679
rect 513004 -3964 513324 56679
rect 513664 -3964 513984 56679
rect 514324 -3964 514644 56679
rect 514984 -3964 515304 56679
rect 515644 -3964 515964 56679
rect 516304 -3964 516624 56679
rect 516964 -3964 517284 56679
rect 526344 -3964 526664 56679
rect 527004 -3964 527324 56679
rect 527664 -3964 527984 56679
rect 528324 -3964 528644 56679
rect 528984 -3964 529304 56679
rect 529644 -3964 529964 56679
rect 530304 -3964 530624 56679
rect 530964 -3964 531284 56679
rect 540344 -3964 540664 56679
rect 541004 -3964 541324 56679
rect 541664 -3964 541984 56679
rect 542324 -3964 542644 56679
rect 542984 -3964 543304 56679
rect 543644 -3964 543964 56679
rect 544304 -3964 544624 56679
rect 544964 -3964 545284 56679
rect 554344 -3964 554664 56679
rect 555004 -3964 555324 56679
rect 555664 -3964 555984 56679
rect 556324 -3964 556644 56679
rect 556984 -3964 557304 56679
rect 557644 -3964 557964 56679
rect 558304 -3964 558624 56679
rect 558964 -3964 559284 56679
rect 568344 -3964 568664 707900
rect 569004 563740 569324 707900
rect 569664 563740 569984 707900
rect 569004 461468 569324 513828
rect 569664 461468 569984 513828
rect 569004 359740 569324 412100
rect 569664 359740 569984 412100
rect 569004 257468 569324 309828
rect 569664 257468 569984 309828
rect 569004 -3964 569324 208100
rect 569664 -3964 569984 208100
rect 570324 -3964 570644 707900
rect 570984 -3964 571304 707900
rect 571644 -3964 571964 707900
rect 572304 -3964 572624 707900
rect 572964 -3964 573284 707900
rect 578612 54352 578932 649584
rect 582344 -3964 582664 707900
rect 584020 656 584340 703280
rect 584680 -4 585000 703940
rect 585340 -664 585660 704600
rect 586000 -1324 586320 705260
rect 586660 -1984 586980 705920
rect 587320 -2644 587640 706580
rect 587980 -3304 588300 707240
rect 588640 -3964 588960 707900
<< obsm4 >>
rect 3371 649664 8264 700909
rect 3371 54272 4820 649664
rect 5300 54272 8264 649664
rect 3371 3571 8264 54272
rect 8744 3571 8924 700909
rect 9404 3571 9584 700909
rect 10064 3571 10244 700909
rect 10724 3571 10904 700909
rect 11384 3571 11564 700909
rect 12044 3571 12224 700909
rect 12704 3571 12884 700909
rect 13364 646129 22264 700909
rect 22744 646129 22924 700909
rect 23404 646129 23584 700909
rect 24064 646129 24244 700909
rect 24724 646129 24904 700909
rect 25384 646129 25564 700909
rect 26044 646129 26224 700909
rect 26704 646129 26884 700909
rect 27364 646129 36264 700909
rect 36744 646129 36924 700909
rect 37404 646129 37584 700909
rect 38064 646129 38244 700909
rect 38724 646129 38904 700909
rect 39384 646129 39564 700909
rect 40044 646129 40224 700909
rect 40704 646129 40884 700909
rect 41364 646129 50264 700909
rect 50744 646129 50924 700909
rect 51404 646129 51584 700909
rect 52064 646129 52244 700909
rect 52724 646129 52904 700909
rect 53384 646129 53564 700909
rect 54044 646129 54224 700909
rect 54704 646129 54884 700909
rect 55364 646129 64264 700909
rect 64744 646129 64924 700909
rect 65404 646129 65584 700909
rect 66064 646129 66244 700909
rect 66724 646129 66904 700909
rect 67384 646129 67564 700909
rect 68044 646129 68224 700909
rect 68704 646129 68884 700909
rect 69364 646129 78264 700909
rect 78744 646129 78924 700909
rect 79404 646129 79584 700909
rect 80064 646129 80244 700909
rect 80724 646129 80904 700909
rect 81384 646129 81564 700909
rect 82044 646129 82224 700909
rect 82704 646129 82884 700909
rect 83364 646129 92264 700909
rect 92744 646129 92924 700909
rect 93404 646129 93584 700909
rect 94064 646129 94244 700909
rect 94724 646129 94904 700909
rect 95384 646129 95564 700909
rect 96044 646129 96224 700909
rect 96704 646129 96884 700909
rect 97364 646129 106264 700909
rect 106744 646129 106924 700909
rect 107404 646129 107584 700909
rect 108064 646129 108244 700909
rect 108724 646129 108904 700909
rect 109384 646129 109564 700909
rect 110044 646129 110224 700909
rect 110704 646129 110884 700909
rect 111364 646129 120264 700909
rect 120744 646129 120924 700909
rect 121404 646129 121584 700909
rect 122064 646129 122244 700909
rect 122724 646129 122904 700909
rect 123384 646129 123564 700909
rect 124044 646129 124224 700909
rect 124704 646129 124884 700909
rect 125364 646129 134264 700909
rect 134744 646129 134924 700909
rect 135404 646129 135584 700909
rect 136064 646129 136244 700909
rect 136724 646129 136904 700909
rect 137384 646129 137564 700909
rect 138044 646129 138224 700909
rect 138704 646129 138884 700909
rect 139364 646129 148264 700909
rect 148744 646129 148924 700909
rect 149404 646129 149584 700909
rect 150064 646129 150244 700909
rect 150724 646129 150904 700909
rect 151384 646129 151564 700909
rect 152044 646129 152224 700909
rect 152704 646129 152884 700909
rect 153364 646129 162264 700909
rect 162744 646129 162924 700909
rect 163404 646129 163584 700909
rect 164064 646129 164244 700909
rect 164724 646129 164904 700909
rect 165384 646129 165564 700909
rect 166044 646129 166224 700909
rect 166704 646129 166884 700909
rect 167364 646129 176264 700909
rect 176744 646129 176924 700909
rect 177404 646129 177584 700909
rect 178064 646129 178244 700909
rect 178724 646129 178904 700909
rect 179384 646129 179564 700909
rect 180044 646129 180224 700909
rect 180704 646129 180884 700909
rect 181364 646129 190264 700909
rect 190744 646129 190924 700909
rect 191404 646129 191584 700909
rect 192064 646129 192244 700909
rect 192724 646129 192904 700909
rect 193384 646129 193564 700909
rect 194044 646129 194224 700909
rect 194704 646129 194884 700909
rect 195364 646129 204264 700909
rect 204744 646129 204924 700909
rect 205404 646129 205584 700909
rect 206064 646129 206244 700909
rect 206724 646129 206904 700909
rect 207384 646129 207564 700909
rect 208044 646129 208224 700909
rect 208704 646129 208884 700909
rect 209364 646129 218264 700909
rect 218744 646129 218924 700909
rect 219404 646129 219584 700909
rect 220064 646129 220244 700909
rect 220724 646129 220904 700909
rect 221384 646129 221564 700909
rect 222044 646129 222224 700909
rect 222704 646129 222884 700909
rect 223364 646129 232264 700909
rect 232744 646129 232924 700909
rect 233404 646129 233584 700909
rect 234064 646129 234244 700909
rect 234724 646129 234904 700909
rect 235384 646129 235564 700909
rect 236044 646129 236224 700909
rect 236704 646129 236884 700909
rect 237364 646129 246264 700909
rect 246744 646129 246924 700909
rect 247404 646129 247584 700909
rect 248064 646129 248244 700909
rect 248724 646129 248904 700909
rect 249384 646129 249564 700909
rect 250044 646129 250224 700909
rect 250704 646129 250884 700909
rect 251364 646129 260264 700909
rect 260744 646129 260924 700909
rect 261404 646129 261584 700909
rect 262064 646129 262244 700909
rect 262724 646129 262904 700909
rect 263384 646129 263564 700909
rect 264044 646129 264224 700909
rect 264704 646129 264884 700909
rect 265364 646129 274264 700909
rect 274744 646129 274924 700909
rect 275404 646129 275584 700909
rect 276064 646129 276244 700909
rect 276724 646129 276904 700909
rect 277384 646129 277564 700909
rect 278044 646129 278224 700909
rect 278704 646129 278884 700909
rect 279364 646129 288264 700909
rect 288744 646129 288924 700909
rect 289404 646129 289584 700909
rect 290064 646129 290244 700909
rect 290724 646129 290904 700909
rect 291384 646129 291564 700909
rect 292044 646129 292224 700909
rect 292704 646129 292884 700909
rect 293364 646129 302264 700909
rect 302744 646129 302924 700909
rect 303404 646129 303584 700909
rect 304064 646129 304244 700909
rect 304724 646129 304904 700909
rect 305384 646129 305564 700909
rect 306044 646129 306224 700909
rect 306704 646129 306884 700909
rect 307364 646129 316264 700909
rect 316744 646129 316924 700909
rect 317404 646129 317584 700909
rect 318064 646129 318244 700909
rect 318724 646129 318904 700909
rect 319384 646129 319564 700909
rect 320044 646129 320224 700909
rect 320704 646129 320884 700909
rect 321364 646129 330264 700909
rect 330744 646129 330924 700909
rect 331404 646129 331584 700909
rect 332064 646129 332244 700909
rect 332724 646129 332904 700909
rect 333384 646129 333564 700909
rect 334044 646129 334224 700909
rect 334704 646129 334884 700909
rect 335364 646129 344264 700909
rect 344744 646129 344924 700909
rect 345404 646129 345584 700909
rect 346064 646129 346244 700909
rect 346724 646129 346904 700909
rect 347384 646129 347564 700909
rect 348044 646129 348224 700909
rect 348704 646129 348884 700909
rect 349364 646129 358264 700909
rect 358744 646129 358924 700909
rect 359404 646129 359584 700909
rect 360064 646129 360244 700909
rect 360724 646129 360904 700909
rect 361384 646129 361564 700909
rect 362044 646129 362224 700909
rect 362704 646129 362884 700909
rect 363364 646129 372264 700909
rect 372744 646129 372924 700909
rect 373404 646129 373584 700909
rect 374064 646129 374244 700909
rect 374724 646129 374904 700909
rect 375384 646129 375564 700909
rect 376044 646129 376224 700909
rect 376704 646129 376884 700909
rect 377364 646129 386264 700909
rect 386744 646129 386924 700909
rect 387404 646129 387584 700909
rect 388064 646129 388244 700909
rect 388724 646129 388904 700909
rect 389384 646129 389564 700909
rect 390044 646129 390224 700909
rect 390704 646129 390884 700909
rect 391364 646129 400264 700909
rect 400744 646129 400924 700909
rect 401404 646129 401584 700909
rect 402064 646129 402244 700909
rect 402724 646129 402904 700909
rect 403384 646129 403564 700909
rect 404044 646129 404224 700909
rect 404704 646129 404884 700909
rect 405364 646129 414264 700909
rect 414744 646129 414924 700909
rect 415404 646129 415584 700909
rect 416064 646129 416244 700909
rect 416724 646129 416904 700909
rect 417384 646129 417564 700909
rect 418044 646129 418224 700909
rect 418704 646129 418884 700909
rect 419364 646129 428264 700909
rect 428744 646129 428924 700909
rect 429404 646129 429584 700909
rect 430064 646129 430244 700909
rect 430724 646129 430904 700909
rect 431384 646129 431564 700909
rect 432044 646129 432224 700909
rect 432704 646129 432884 700909
rect 433364 646129 442264 700909
rect 442744 646129 442924 700909
rect 443404 646129 443584 700909
rect 444064 646129 444244 700909
rect 444724 646129 444904 700909
rect 445384 646129 445564 700909
rect 446044 646129 446224 700909
rect 446704 646129 446884 700909
rect 447364 646129 456264 700909
rect 456744 646129 456924 700909
rect 457404 646129 457584 700909
rect 458064 646129 458244 700909
rect 458724 646129 458904 700909
rect 459384 646129 459564 700909
rect 460044 646129 460224 700909
rect 460704 646129 460884 700909
rect 461364 646129 470264 700909
rect 470744 646129 470924 700909
rect 471404 646129 471584 700909
rect 472064 646129 472244 700909
rect 472724 646129 472904 700909
rect 473384 646129 473564 700909
rect 474044 646129 474224 700909
rect 474704 646129 474884 700909
rect 475364 646129 484264 700909
rect 484744 646129 484924 700909
rect 485404 646129 485584 700909
rect 486064 646129 486244 700909
rect 486724 646129 486904 700909
rect 487384 646129 487564 700909
rect 488044 646129 488224 700909
rect 488704 646129 488884 700909
rect 489364 646129 498264 700909
rect 498744 646129 498924 700909
rect 499404 646129 499584 700909
rect 500064 646129 500244 700909
rect 500724 646129 500904 700909
rect 501384 646129 501564 700909
rect 502044 646129 502224 700909
rect 502704 646129 502884 700909
rect 503364 646129 512264 700909
rect 512744 646129 512924 700909
rect 513404 646129 513584 700909
rect 514064 646129 514244 700909
rect 514724 646129 514904 700909
rect 515384 646129 515564 700909
rect 516044 646129 516224 700909
rect 516704 646129 516884 700909
rect 517364 646129 526264 700909
rect 526744 646129 526924 700909
rect 527404 646129 527584 700909
rect 528064 646129 528244 700909
rect 528724 646129 528904 700909
rect 529384 646129 529564 700909
rect 530044 646129 530224 700909
rect 530704 646129 530884 700909
rect 531364 646129 540264 700909
rect 540744 646129 540924 700909
rect 541404 646129 541584 700909
rect 542064 646129 542244 700909
rect 542724 646129 542904 700909
rect 543384 646129 543564 700909
rect 544044 646129 544224 700909
rect 544704 646129 544884 700909
rect 545364 646129 554264 700909
rect 554744 646129 554924 700909
rect 555404 646129 555584 700909
rect 556064 646129 556244 700909
rect 556724 646129 556904 700909
rect 557384 646129 557564 700909
rect 558044 646129 558224 700909
rect 558704 646129 558884 700909
rect 559364 646129 568264 700909
rect 13364 56759 568264 646129
rect 13364 3571 22264 56759
rect 22744 3571 22924 56759
rect 23404 3571 23584 56759
rect 24064 3571 24244 56759
rect 24724 3571 24904 56759
rect 25384 3571 25564 56759
rect 26044 3571 26224 56759
rect 26704 3571 26884 56759
rect 27364 3571 36264 56759
rect 36744 3571 36924 56759
rect 37404 3571 37584 56759
rect 38064 3571 38244 56759
rect 38724 3571 38904 56759
rect 39384 3571 39564 56759
rect 40044 3571 40224 56759
rect 40704 3571 40884 56759
rect 41364 3571 50264 56759
rect 50744 3571 50924 56759
rect 51404 3571 51584 56759
rect 52064 3571 52244 56759
rect 52724 3571 52904 56759
rect 53384 3571 53564 56759
rect 54044 3571 54224 56759
rect 54704 3571 54884 56759
rect 55364 3571 64264 56759
rect 64744 3571 64924 56759
rect 65404 3571 65584 56759
rect 66064 3571 66244 56759
rect 66724 3571 66904 56759
rect 67384 3571 67564 56759
rect 68044 3571 68224 56759
rect 68704 3571 68884 56759
rect 69364 3571 78264 56759
rect 78744 3571 78924 56759
rect 79404 3571 79584 56759
rect 80064 3571 80244 56759
rect 80724 3571 80904 56759
rect 81384 3571 81564 56759
rect 82044 3571 82224 56759
rect 82704 3571 82884 56759
rect 83364 3571 92264 56759
rect 92744 3571 92924 56759
rect 93404 3571 93584 56759
rect 94064 3571 94244 56759
rect 94724 3571 94904 56759
rect 95384 3571 95564 56759
rect 96044 3571 96224 56759
rect 96704 3571 96884 56759
rect 97364 3571 106264 56759
rect 106744 3571 106924 56759
rect 107404 3571 107584 56759
rect 108064 3571 108244 56759
rect 108724 3571 108904 56759
rect 109384 3571 109564 56759
rect 110044 3571 110224 56759
rect 110704 3571 110884 56759
rect 111364 3571 120264 56759
rect 120744 3571 120924 56759
rect 121404 3571 121584 56759
rect 122064 3571 122244 56759
rect 122724 3571 122904 56759
rect 123384 3571 123564 56759
rect 124044 3571 124224 56759
rect 124704 3571 124884 56759
rect 125364 3571 134264 56759
rect 134744 3571 134924 56759
rect 135404 3571 135584 56759
rect 136064 3571 136244 56759
rect 136724 3571 136904 56759
rect 137384 3571 137564 56759
rect 138044 3571 138224 56759
rect 138704 3571 138884 56759
rect 139364 3571 148264 56759
rect 148744 3571 148924 56759
rect 149404 3571 149584 56759
rect 150064 3571 150244 56759
rect 150724 3571 150904 56759
rect 151384 3571 151564 56759
rect 152044 3571 152224 56759
rect 152704 3571 152884 56759
rect 153364 3571 162264 56759
rect 162744 3571 162924 56759
rect 163404 3571 163584 56759
rect 164064 3571 164244 56759
rect 164724 3571 164904 56759
rect 165384 3571 165564 56759
rect 166044 3571 166224 56759
rect 166704 3571 166884 56759
rect 167364 3571 176264 56759
rect 176744 3571 176924 56759
rect 177404 3571 177584 56759
rect 178064 3571 178244 56759
rect 178724 3571 178904 56759
rect 179384 3571 179564 56759
rect 180044 3571 180224 56759
rect 180704 3571 180884 56759
rect 181364 3571 190264 56759
rect 190744 3571 190924 56759
rect 191404 3571 191584 56759
rect 192064 3571 192244 56759
rect 192724 3571 192904 56759
rect 193384 3571 193564 56759
rect 194044 3571 194224 56759
rect 194704 3571 194884 56759
rect 195364 3571 204264 56759
rect 204744 3571 204924 56759
rect 205404 3571 205584 56759
rect 206064 3571 206244 56759
rect 206724 3571 206904 56759
rect 207384 3571 207564 56759
rect 208044 3571 208224 56759
rect 208704 3571 208884 56759
rect 209364 3571 218264 56759
rect 218744 3571 218924 56759
rect 219404 3571 219584 56759
rect 220064 3571 220244 56759
rect 220724 3571 220904 56759
rect 221384 3571 221564 56759
rect 222044 3571 222224 56759
rect 222704 3571 222884 56759
rect 223364 3571 232264 56759
rect 232744 3571 232924 56759
rect 233404 3571 233584 56759
rect 234064 3571 234244 56759
rect 234724 3571 234904 56759
rect 235384 3571 235564 56759
rect 236044 3571 236224 56759
rect 236704 3571 236884 56759
rect 237364 3571 246264 56759
rect 246744 3571 246924 56759
rect 247404 3571 247584 56759
rect 248064 3571 248244 56759
rect 248724 3571 248904 56759
rect 249384 3571 249564 56759
rect 250044 3571 250224 56759
rect 250704 3571 250884 56759
rect 251364 3571 260264 56759
rect 260744 3571 260924 56759
rect 261404 3571 261584 56759
rect 262064 3571 262244 56759
rect 262724 3571 262904 56759
rect 263384 3571 263564 56759
rect 264044 3571 264224 56759
rect 264704 3571 264884 56759
rect 265364 3571 274264 56759
rect 274744 3571 274924 56759
rect 275404 3571 275584 56759
rect 276064 3571 276244 56759
rect 276724 3571 276904 56759
rect 277384 3571 277564 56759
rect 278044 3571 278224 56759
rect 278704 3571 278884 56759
rect 279364 3571 288264 56759
rect 288744 3571 288924 56759
rect 289404 3571 289584 56759
rect 290064 3571 290244 56759
rect 290724 3571 290904 56759
rect 291384 3571 291564 56759
rect 292044 3571 292224 56759
rect 292704 3571 292884 56759
rect 293364 3571 302264 56759
rect 302744 3571 302924 56759
rect 303404 3571 303584 56759
rect 304064 3571 304244 56759
rect 304724 3571 304904 56759
rect 305384 3571 305564 56759
rect 306044 3571 306224 56759
rect 306704 3571 306884 56759
rect 307364 3571 316264 56759
rect 316744 3571 316924 56759
rect 317404 3571 317584 56759
rect 318064 3571 318244 56759
rect 318724 3571 318904 56759
rect 319384 3571 319564 56759
rect 320044 3571 320224 56759
rect 320704 3571 320884 56759
rect 321364 3571 330264 56759
rect 330744 3571 330924 56759
rect 331404 3571 331584 56759
rect 332064 3571 332244 56759
rect 332724 3571 332904 56759
rect 333384 3571 333564 56759
rect 334044 3571 334224 56759
rect 334704 3571 334884 56759
rect 335364 3571 344264 56759
rect 344744 3571 344924 56759
rect 345404 3571 345584 56759
rect 346064 3571 346244 56759
rect 346724 3571 346904 56759
rect 347384 3571 347564 56759
rect 348044 3571 348224 56759
rect 348704 3571 348884 56759
rect 349364 3571 358264 56759
rect 358744 3571 358924 56759
rect 359404 3571 359584 56759
rect 360064 3571 360244 56759
rect 360724 3571 360904 56759
rect 361384 3571 361564 56759
rect 362044 3571 362224 56759
rect 362704 3571 362884 56759
rect 363364 3571 372264 56759
rect 372744 3571 372924 56759
rect 373404 3571 373584 56759
rect 374064 3571 374244 56759
rect 374724 3571 374904 56759
rect 375384 3571 375564 56759
rect 376044 3571 376224 56759
rect 376704 3571 376884 56759
rect 377364 3571 386264 56759
rect 386744 3571 386924 56759
rect 387404 3571 387584 56759
rect 388064 3571 388244 56759
rect 388724 3571 388904 56759
rect 389384 3571 389564 56759
rect 390044 3571 390224 56759
rect 390704 3571 390884 56759
rect 391364 3571 400264 56759
rect 400744 3571 400924 56759
rect 401404 3571 401584 56759
rect 402064 3571 402244 56759
rect 402724 3571 402904 56759
rect 403384 3571 403564 56759
rect 404044 3571 404224 56759
rect 404704 3571 404884 56759
rect 405364 3571 414264 56759
rect 414744 3571 414924 56759
rect 415404 3571 415584 56759
rect 416064 3571 416244 56759
rect 416724 3571 416904 56759
rect 417384 3571 417564 56759
rect 418044 3571 418224 56759
rect 418704 3571 418884 56759
rect 419364 3571 428264 56759
rect 428744 3571 428924 56759
rect 429404 3571 429584 56759
rect 430064 3571 430244 56759
rect 430724 3571 430904 56759
rect 431384 3571 431564 56759
rect 432044 3571 432224 56759
rect 432704 3571 432884 56759
rect 433364 3571 442264 56759
rect 442744 3571 442924 56759
rect 443404 3571 443584 56759
rect 444064 3571 444244 56759
rect 444724 3571 444904 56759
rect 445384 3571 445564 56759
rect 446044 3571 446224 56759
rect 446704 3571 446884 56759
rect 447364 3571 456264 56759
rect 456744 3571 456924 56759
rect 457404 3571 457584 56759
rect 458064 3571 458244 56759
rect 458724 3571 458904 56759
rect 459384 3571 459564 56759
rect 460044 3571 460224 56759
rect 460704 3571 460884 56759
rect 461364 3571 470264 56759
rect 470744 3571 470924 56759
rect 471404 3571 471584 56759
rect 472064 3571 472244 56759
rect 472724 3571 472904 56759
rect 473384 3571 473564 56759
rect 474044 3571 474224 56759
rect 474704 3571 474884 56759
rect 475364 3571 484264 56759
rect 484744 3571 484924 56759
rect 485404 3571 485584 56759
rect 486064 3571 486244 56759
rect 486724 3571 486904 56759
rect 487384 3571 487564 56759
rect 488044 3571 488224 56759
rect 488704 3571 488884 56759
rect 489364 3571 498264 56759
rect 498744 3571 498924 56759
rect 499404 3571 499584 56759
rect 500064 3571 500244 56759
rect 500724 3571 500904 56759
rect 501384 3571 501564 56759
rect 502044 3571 502224 56759
rect 502704 3571 502884 56759
rect 503364 3571 512264 56759
rect 512744 3571 512924 56759
rect 513404 3571 513584 56759
rect 514064 3571 514244 56759
rect 514724 3571 514904 56759
rect 515384 3571 515564 56759
rect 516044 3571 516224 56759
rect 516704 3571 516884 56759
rect 517364 3571 526264 56759
rect 526744 3571 526924 56759
rect 527404 3571 527584 56759
rect 528064 3571 528244 56759
rect 528724 3571 528904 56759
rect 529384 3571 529564 56759
rect 530044 3571 530224 56759
rect 530704 3571 530884 56759
rect 531364 3571 540264 56759
rect 540744 3571 540924 56759
rect 541404 3571 541584 56759
rect 542064 3571 542244 56759
rect 542724 3571 542904 56759
rect 543384 3571 543564 56759
rect 544044 3571 544224 56759
rect 544704 3571 544884 56759
rect 545364 3571 554264 56759
rect 554744 3571 554924 56759
rect 555404 3571 555584 56759
rect 556064 3571 556244 56759
rect 556724 3571 556904 56759
rect 557384 3571 557564 56759
rect 558044 3571 558224 56759
rect 558704 3571 558884 56759
rect 559364 3571 568264 56759
rect 568744 563660 568924 700909
rect 569404 563660 569584 700909
rect 570064 563660 570244 700909
rect 568744 513908 570244 563660
rect 568744 461388 568924 513908
rect 569404 461388 569584 513908
rect 570064 461388 570244 513908
rect 568744 412180 570244 461388
rect 568744 359660 568924 412180
rect 569404 359660 569584 412180
rect 570064 359660 570244 412180
rect 568744 309908 570244 359660
rect 568744 257388 568924 309908
rect 569404 257388 569584 309908
rect 570064 257388 570244 309908
rect 568744 208180 570244 257388
rect 568744 3571 568924 208180
rect 569404 3571 569584 208180
rect 570064 3571 570244 208180
rect 570724 3571 570904 700909
rect 571384 3571 571564 700909
rect 572044 3571 572224 700909
rect 572704 3571 572884 700909
rect 573364 3571 574389 700909
<< metal5 >>
rect -5036 707580 588960 707900
rect -4376 706920 588300 707240
rect -3716 706260 587640 706580
rect -3056 705600 586980 705920
rect -2396 704940 586320 705260
rect -1736 704280 585660 704600
rect -1076 703620 585000 703940
rect -416 702960 584340 703280
rect -5036 701396 588960 701716
rect -5036 700736 588960 701056
rect -5036 700076 588960 700396
rect -5036 699416 588960 699736
rect -5036 689036 588960 689356
rect -5036 688376 588960 688696
rect -5036 687716 588960 688036
rect -5036 687056 588960 687376
rect -5036 686396 588960 686716
rect -5036 685736 588960 686056
rect -5036 685076 588960 685396
rect -5036 684416 588960 684736
rect -5036 674036 588960 674356
rect -5036 673376 588960 673696
rect -5036 672716 588960 673036
rect -5036 672056 588960 672376
rect -5036 671396 588960 671716
rect -5036 670736 588960 671056
rect -5036 670076 588960 670396
rect -5036 669416 588960 669736
rect -5036 659036 588960 659356
rect -5036 658376 588960 658696
rect -5036 657716 588960 658036
rect -5036 657056 588960 657376
rect -5036 656396 588960 656716
rect -5036 655736 588960 656056
rect -5036 655076 588960 655396
rect -5036 654416 588960 654736
rect -5036 644036 588960 644356
rect -5036 643376 588960 643696
rect -5036 642716 588960 643036
rect -5036 642056 588960 642376
rect -5036 641396 588960 641716
rect -5036 640736 588960 641056
rect -5036 640076 588960 640396
rect -5036 639416 588960 639736
rect -5036 629036 588960 629356
rect -5036 628376 588960 628696
rect -5036 627716 588960 628036
rect -5036 627056 588960 627376
rect -5036 626396 588960 626716
rect -5036 625736 588960 626056
rect -5036 625076 588960 625396
rect -5036 624416 588960 624736
rect -5036 614036 588960 614356
rect -5036 613376 588960 613696
rect -5036 612716 588960 613036
rect -5036 612056 588960 612376
rect -5036 611396 588960 611716
rect -5036 610736 588960 611056
rect -5036 610076 588960 610396
rect -5036 609416 588960 609736
rect -5036 599036 588960 599356
rect -5036 598376 588960 598696
rect -5036 597716 588960 598036
rect -5036 597056 588960 597376
rect -5036 596396 588960 596716
rect -5036 595736 588960 596056
rect -5036 595076 588960 595396
rect -5036 594416 588960 594736
rect -5036 584036 588960 584356
rect -5036 583376 588960 583696
rect -5036 582716 588960 583036
rect -5036 582056 588960 582376
rect -5036 581396 588960 581716
rect -5036 580736 588960 581056
rect -5036 580076 588960 580396
rect -5036 579416 588960 579736
rect -5036 569036 588960 569356
rect -5036 568376 588960 568696
rect -5036 567716 588960 568036
rect -5036 567056 588960 567376
rect -5036 566396 588960 566716
rect -5036 565736 588960 566056
rect -5036 565076 588960 565396
rect -5036 564416 588960 564736
rect -5036 554036 588960 554356
rect -5036 553376 588960 553696
rect -5036 552716 588960 553036
rect -5036 552056 588960 552376
rect -5036 551396 588960 551716
rect -5036 550736 588960 551056
rect -5036 550076 588960 550396
rect -5036 549416 588960 549736
rect -5036 539036 588960 539356
rect -5036 538376 588960 538696
rect -5036 537716 588960 538036
rect -5036 537056 588960 537376
rect -5036 536396 588960 536716
rect -5036 535736 588960 536056
rect -5036 535076 588960 535396
rect -5036 534416 588960 534736
rect -5036 524036 588960 524356
rect -5036 523376 588960 523696
rect -5036 522716 588960 523036
rect -5036 522056 588960 522376
rect -5036 521396 588960 521716
rect -5036 520736 588960 521056
rect -5036 520076 588960 520396
rect -5036 519416 588960 519736
rect -5036 509036 588960 509356
rect -5036 508376 588960 508696
rect -5036 507716 588960 508036
rect -5036 507056 588960 507376
rect -5036 506396 588960 506716
rect -5036 505736 588960 506056
rect -5036 505076 588960 505396
rect -5036 504416 588960 504736
rect -5036 494036 588960 494356
rect -5036 493376 588960 493696
rect -5036 492716 588960 493036
rect -5036 492056 588960 492376
rect -5036 491396 588960 491716
rect -5036 490736 588960 491056
rect -5036 490076 588960 490396
rect -5036 489416 588960 489736
rect -5036 479036 588960 479356
rect -5036 478376 588960 478696
rect -5036 477716 588960 478036
rect -5036 477056 588960 477376
rect -5036 476396 588960 476716
rect -5036 475736 588960 476056
rect -5036 475076 588960 475396
rect -5036 474416 588960 474736
rect -5036 464036 588960 464356
rect -5036 463376 588960 463696
rect -5036 462716 588960 463036
rect -5036 462056 588960 462376
rect -5036 461396 588960 461716
rect -5036 460736 588960 461056
rect -5036 460076 588960 460396
rect -5036 459416 588960 459736
rect -5036 449036 588960 449356
rect -5036 448376 588960 448696
rect -5036 447716 588960 448036
rect -5036 447056 588960 447376
rect -5036 446396 588960 446716
rect -5036 445736 588960 446056
rect -5036 445076 588960 445396
rect -5036 444416 588960 444736
rect -5036 434036 588960 434356
rect -5036 433376 588960 433696
rect -5036 432716 588960 433036
rect -5036 432056 588960 432376
rect -5036 431396 588960 431716
rect -5036 430736 588960 431056
rect -5036 430076 588960 430396
rect -5036 429416 588960 429736
rect -5036 419036 588960 419356
rect -5036 418376 588960 418696
rect -5036 417716 588960 418036
rect -5036 417056 588960 417376
rect -5036 416396 588960 416716
rect -5036 415736 588960 416056
rect -5036 415076 588960 415396
rect -5036 414416 588960 414736
rect -5036 404036 588960 404356
rect -5036 403376 588960 403696
rect -5036 402716 588960 403036
rect -5036 402056 588960 402376
rect -5036 401396 588960 401716
rect -5036 400736 588960 401056
rect -5036 400076 588960 400396
rect -5036 399416 588960 399736
rect -5036 389036 588960 389356
rect -5036 388376 588960 388696
rect -5036 387716 588960 388036
rect -5036 387056 588960 387376
rect -5036 386396 588960 386716
rect -5036 385736 588960 386056
rect -5036 385076 588960 385396
rect -5036 384416 588960 384736
rect -5036 374036 588960 374356
rect -5036 373376 588960 373696
rect -5036 372716 588960 373036
rect -5036 372056 588960 372376
rect -5036 371396 588960 371716
rect -5036 370736 588960 371056
rect -5036 370076 588960 370396
rect -5036 369416 588960 369736
rect -5036 359036 588960 359356
rect -5036 358376 588960 358696
rect -5036 357716 588960 358036
rect -5036 357056 588960 357376
rect -5036 356396 588960 356716
rect -5036 355736 588960 356056
rect -5036 355076 588960 355396
rect -5036 354416 588960 354736
rect -5036 344036 588960 344356
rect -5036 343376 588960 343696
rect -5036 342716 588960 343036
rect -5036 342056 588960 342376
rect -5036 341396 588960 341716
rect -5036 340736 588960 341056
rect -5036 340076 588960 340396
rect -5036 339416 588960 339736
rect -5036 329036 588960 329356
rect -5036 328376 588960 328696
rect -5036 327716 588960 328036
rect -5036 327056 588960 327376
rect -5036 326396 588960 326716
rect -5036 325736 588960 326056
rect -5036 325076 588960 325396
rect -5036 324416 588960 324736
rect -5036 314036 588960 314356
rect -5036 313376 588960 313696
rect -5036 312716 588960 313036
rect -5036 312056 588960 312376
rect -5036 311396 588960 311716
rect -5036 310736 588960 311056
rect -5036 310076 588960 310396
rect -5036 309416 588960 309736
rect -5036 299036 588960 299356
rect -5036 298376 588960 298696
rect -5036 297716 588960 298036
rect -5036 297056 588960 297376
rect -5036 296396 588960 296716
rect -5036 295736 588960 296056
rect -5036 295076 588960 295396
rect -5036 294416 588960 294736
rect -5036 284036 588960 284356
rect -5036 283376 588960 283696
rect -5036 282716 588960 283036
rect -5036 282056 588960 282376
rect -5036 281396 588960 281716
rect -5036 280736 588960 281056
rect -5036 280076 588960 280396
rect -5036 279416 588960 279736
rect -5036 269036 588960 269356
rect -5036 268376 588960 268696
rect -5036 267716 588960 268036
rect -5036 267056 588960 267376
rect -5036 266396 588960 266716
rect -5036 265736 588960 266056
rect -5036 265076 588960 265396
rect -5036 264416 588960 264736
rect -5036 254036 588960 254356
rect -5036 253376 588960 253696
rect -5036 252716 588960 253036
rect -5036 252056 588960 252376
rect -5036 251396 588960 251716
rect -5036 250736 588960 251056
rect -5036 250076 588960 250396
rect -5036 249416 588960 249736
rect -5036 239036 588960 239356
rect -5036 238376 588960 238696
rect -5036 237716 588960 238036
rect -5036 237056 588960 237376
rect -5036 236396 588960 236716
rect -5036 235736 588960 236056
rect -5036 235076 588960 235396
rect -5036 234416 588960 234736
rect -5036 224036 588960 224356
rect -5036 223376 588960 223696
rect -5036 222716 588960 223036
rect -5036 222056 588960 222376
rect -5036 221396 588960 221716
rect -5036 220736 588960 221056
rect -5036 220076 588960 220396
rect -5036 219416 588960 219736
rect -5036 209036 588960 209356
rect -5036 208376 588960 208696
rect -5036 207716 465010 208036
rect -5036 207056 465010 207376
rect -5036 206396 465010 206716
rect 498630 207716 588960 208036
rect 498630 207056 588960 207376
rect 498630 206396 588960 206716
rect -5036 205736 588960 206056
rect -5036 205076 588960 205396
rect -5036 204416 588960 204736
rect -5036 194036 588960 194356
rect -5036 193376 588960 193696
rect -5036 192716 588960 193036
rect -5036 192056 588960 192376
rect -5036 191396 588960 191716
rect -5036 190736 588960 191056
rect -5036 190076 588960 190396
rect -5036 189416 588960 189736
rect -5036 179036 588960 179356
rect -5036 178376 588960 178696
rect -5036 177716 588960 178036
rect -5036 177056 588960 177376
rect -5036 176396 588960 176716
rect -5036 175736 588960 176056
rect -5036 175076 588960 175396
rect -5036 174416 588960 174736
rect -5036 164036 588960 164356
rect -5036 163376 588960 163696
rect -5036 162716 588960 163036
rect -5036 162056 588960 162376
rect -5036 161396 588960 161716
rect -5036 160736 588960 161056
rect -5036 160076 588960 160396
rect -5036 159416 588960 159736
rect -5036 149036 588960 149356
rect -5036 148376 588960 148696
rect -5036 147716 588960 148036
rect -5036 147056 588960 147376
rect -5036 146396 588960 146716
rect -5036 145736 588960 146056
rect -5036 145076 588960 145396
rect -5036 144416 588960 144736
rect -5036 134036 588960 134356
rect -5036 133376 588960 133696
rect -5036 132716 588960 133036
rect -5036 132056 588960 132376
rect -5036 131396 588960 131716
rect -5036 130736 588960 131056
rect -5036 130076 588960 130396
rect -5036 129416 588960 129736
rect -5036 119036 588960 119356
rect -5036 118376 588960 118696
rect -5036 117716 588960 118036
rect -5036 117056 588960 117376
rect -5036 116396 588960 116716
rect -5036 115736 588960 116056
rect -5036 115076 588960 115396
rect -5036 114416 588960 114736
rect -5036 104036 588960 104356
rect -5036 103376 588960 103696
rect -5036 102716 588960 103036
rect -5036 102056 588960 102376
rect -5036 101396 588960 101716
rect -5036 100736 588960 101056
rect -5036 100076 588960 100396
rect -5036 99416 588960 99736
rect -5036 89036 588960 89356
rect -5036 88376 588960 88696
rect -5036 87716 588960 88036
rect -5036 87056 588960 87376
rect -5036 86396 588960 86716
rect -5036 85736 588960 86056
rect -5036 85076 588960 85396
rect -5036 84416 588960 84736
rect -5036 74036 588960 74356
rect -5036 73376 588960 73696
rect -5036 72716 588960 73036
rect -5036 72056 588960 72376
rect -5036 71396 588960 71716
rect -5036 70736 588960 71056
rect -5036 70076 588960 70396
rect -5036 69416 588960 69736
rect -5036 59036 588960 59356
rect -5036 58376 588960 58696
rect -5036 57716 588960 58036
rect -5036 57056 588960 57376
rect -5036 56396 588960 56716
rect -5036 55736 588960 56056
rect -5036 55076 588960 55396
rect -5036 54416 588960 54736
rect -5036 44036 588960 44356
rect -5036 43376 588960 43696
rect -5036 42716 588960 43036
rect -5036 42056 588960 42376
rect -5036 41396 588960 41716
rect -5036 40736 588960 41056
rect -5036 40076 588960 40396
rect -5036 39416 588960 39736
rect -5036 29036 588960 29356
rect -5036 28376 588960 28696
rect -5036 27716 588960 28036
rect -5036 27056 588960 27376
rect -5036 26396 588960 26716
rect -5036 25736 588960 26056
rect -5036 25076 588960 25396
rect -5036 24416 588960 24736
rect -5036 14036 588960 14356
rect -5036 13376 588960 13696
rect -5036 12716 588960 13036
rect -5036 12056 588960 12376
rect -5036 11396 588960 11716
rect -5036 10736 588960 11056
rect -5036 10076 588960 10396
rect -5036 9416 588960 9736
rect -416 656 584340 976
rect -1076 -4 585000 316
rect -1736 -664 585660 -344
rect -2396 -1324 586320 -1004
rect -3056 -1984 586980 -1664
rect -3716 -2644 587640 -2324
rect -4376 -3304 588300 -2984
rect -5036 -3964 588960 -3644
<< obsm5 >>
rect 12042 629676 571866 637196
rect 12042 614676 571866 624096
rect 12042 599676 571866 609096
rect 12042 584676 571866 594096
rect 12042 569676 571866 579096
rect 12042 554676 571866 564096
rect 12042 539676 571866 549096
rect 12042 524676 571866 534096
rect 12042 509676 571866 519096
rect 12042 494676 571866 504096
rect 12042 479676 571866 489096
rect 12042 464676 571866 474096
rect 12042 449676 571866 459096
rect 12042 434676 571866 444096
rect 12042 419676 571866 429096
rect 12042 404676 571866 414096
rect 12042 389676 571866 399096
rect 12042 374676 571866 384096
rect 12042 359676 571866 369096
rect 12042 344676 571866 354096
rect 12042 329676 571866 339096
rect 12042 314676 571866 324096
rect 12042 299676 571866 309096
rect 12042 284676 571866 294096
rect 12042 269676 571866 279096
rect 12042 254676 571866 264096
rect 12042 239676 571866 249096
rect 12042 224676 571866 234096
rect 12042 209676 571866 219096
rect 465330 206376 498310 208056
rect 12042 194676 571866 204096
rect 12042 179676 571866 189096
rect 12042 164676 571866 174096
rect 12042 149676 571866 159096
rect 12042 134676 571866 144096
rect 12042 119676 571866 129096
rect 12042 104676 571866 114096
rect 12042 89676 571866 99096
rect 12042 74676 571866 84096
rect 12042 66216 571866 69096
<< labels >>
rlabel metal2 s 373538 703200 373594 703800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 583200 656208 583800 656328 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583200 299888 583800 300008 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 164882 200 164938 800 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 498474 200 498530 800 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 420550 703200 420606 703800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 583200 175448 583800 175568 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 129462 200 129518 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 78586 200 78642 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 583200 63248 583800 63368 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 583200 590248 583800 590368 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 318798 703200 318854 703800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 200 128528 800 128648 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 583200 233248 583800 233368 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 377402 703200 377458 703800 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 204166 200 204222 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 515218 703200 515274 703800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 251178 200 251234 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 583200 639888 583800 640008 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 583200 701768 583800 701888 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 200 609288 800 609408 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 169390 703200 169446 703800 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 200 443368 800 443488 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 244094 703200 244150 703800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 200 522248 800 522368 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 200 451528 800 451648 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583200 187688 583800 187808 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal3 s 200 82968 800 83088 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 583200 586168 583800 586288 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583200 602488 583800 602608 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 200 41488 800 41608 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583200 312128 583800 312248 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 452106 703200 452162 703800 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 122378 703200 122434 703800 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 130106 703200 130162 703800 6 io_in[14]
port 35 nsew signal input
rlabel metal3 s 200 700408 800 700528 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 200 617448 800 617568 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 153290 703200 153346 703800 6 io_in[17]
port 38 nsew signal input
rlabel metal3 s 200 464448 800 464568 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 157798 703200 157854 703800 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 200 675928 800 676048 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 423770 200 423826 800 6 io_in[20]
port 42 nsew signal input
rlabel metal3 s 583200 561008 583800 561128 6 io_in[21]
port 43 nsew signal input
rlabel metal3 s 583200 199928 583800 200048 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 227350 200 227406 800 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 259550 703200 259606 703800 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 583200 125128 583800 125248 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 200 8168 800 8288 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 200 348168 800 348288 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 566094 703200 566150 703800 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 583200 179528 583800 179648 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 200 555568 800 555688 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 569958 703200 570014 703800 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 43810 703200 43866 703800 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 583200 229168 583800 229288 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 583200 46928 583800 47048 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 200 646688 800 646808 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 381266 703200 381322 703800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 184846 703200 184902 703800 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 583200 162528 583800 162648 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 499118 703200 499174 703800 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 200 588888 800 589008 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 419906 200 419962 800 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 200 306688 800 306808 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583200 697688 583800 697808 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 502338 200 502394 800 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 483018 200 483074 800 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 550638 703200 550694 703800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 152646 200 152702 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 117870 200 117926 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583200 42168 583800 42288 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583200 357688 583800 357808 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583200 573248 583800 573368 6 io_oeb[14]
port 73 nsew signal output
rlabel metal3 s 200 460368 800 460488 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 522302 200 522358 800 6 io_oeb[16]
port 75 nsew signal output
rlabel metal3 s 583200 88408 583800 88528 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 8390 703200 8446 703800 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 538402 703200 538458 703800 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 200 597048 800 597168 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 200 20408 800 20528 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 357438 200 357494 800 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 479154 200 479210 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 200 281528 800 281648 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 583200 544688 583800 544808 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 200 207408 800 207528 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 583200 333208 583800 333328 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 55402 703200 55458 703800 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 200 174088 800 174208 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 200 488928 800 489048 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 200 634448 800 634568 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 583200 635808 583800 635928 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 522946 703200 523002 703800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 583200 142128 583800 142248 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 279514 703200 279570 703800 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 79230 703200 79286 703800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 305918 200 305974 800 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 200 592968 800 593088 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 200 692248 800 692368 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583200 594328 583800 594448 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 408958 703200 409014 703800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 200 476688 800 476808 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 282734 200 282790 800 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 54758 200 54814 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583200 25848 583800 25968 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 240230 703200 240286 703800 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 561586 200 561642 800 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 200 91128 800 91248 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 200 431128 800 431248 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 200 654848 800 654968 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583200 515448 583800 515568 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 455970 703200 456026 703800 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 58622 200 58678 800 6 io_out[16]
port 113 nsew signal output
rlabel metal3 s 200 385568 800 385688 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 200 211488 800 211608 6 io_out[18]
port 115 nsew signal output
rlabel metal3 s 583200 395088 583800 395208 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 200 389648 800 389768 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 94042 200 94098 800 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 12254 703200 12310 703800 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 30930 200 30986 800 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 266634 200 266690 800 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 583200 511368 583800 511488 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 180982 703200 181038 703800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 271786 703200 271842 703800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 459190 200 459246 800 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 141698 703200 141754 703800 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 583200 171368 583800 171488 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583200 499128 583800 499248 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 82450 200 82506 800 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 247314 200 247370 800 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 583200 486208 583800 486328 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 583200 349528 583800 349648 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 443734 200 443790 800 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 97906 200 97962 800 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 463698 703200 463754 703800 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 161018 200 161074 800 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 157154 200 157210 800 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 39302 200 39358 800 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 397366 703200 397422 703800 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 200 198568 800 198688 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583200 465808 583800 465928 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 318154 200 318210 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583200 262488 583800 262608 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 200 422968 800 423088 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 145562 703200 145618 703800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 224130 703200 224186 703800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 137834 703200 137890 703800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal3 s 583200 665048 583800 665168 6 la_data_in[103]
port 148 nsew signal input
rlabel metal3 s 583200 320288 583800 320408 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 200 186328 800 186448 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 200 658928 800 659048 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 200 323008 800 323128 6 la_data_in[107]
port 152 nsew signal input
rlabel metal3 s 200 547408 800 547528 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 126242 703200 126298 703800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 200 684088 800 684208 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 286598 200 286654 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 314934 703200 314990 703800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 200 32648 800 32768 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 109498 200 109554 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal3 s 200 447448 800 447568 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 404450 200 404506 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 583200 673208 583800 673328 6 la_data_in[116]
port 162 nsew signal input
rlabel metal3 s 583200 337288 583800 337408 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 365166 200 365222 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 583200 482128 583800 482248 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 200 360408 800 360528 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 212538 703200 212594 703800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal3 s 583200 535848 583800 535968 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 193218 703200 193274 703800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal3 s 583200 469888 583800 470008 6 la_data_in[123]
port 170 nsew signal input
rlabel metal3 s 583200 316208 583800 316328 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 451462 200 451518 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 428922 703200 428978 703800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal3 s 583200 121048 583800 121168 6 la_data_in[127]
port 174 nsew signal input
rlabel metal3 s 200 257048 800 257168 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 583200 490288 583800 490408 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 495254 703200 495310 703800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 177118 703200 177174 703800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 583200 556928 583800 557048 6 la_data_in[16]
port 179 nsew signal input
rlabel metal3 s 583200 59168 583800 59288 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 583200 51008 583800 51128 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 311070 703200 311126 703800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 200 551488 800 551608 6 la_data_in[1]
port 183 nsew signal input
rlabel metal3 s 200 136688 800 136808 6 la_data_in[20]
port 184 nsew signal input
rlabel metal3 s 583200 129888 583800 130008 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 200 393728 800 393848 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 200 688168 800 688288 6 la_data_in[23]
port 187 nsew signal input
rlabel metal3 s 200 240048 800 240168 6 la_data_in[24]
port 188 nsew signal input
rlabel metal3 s 200 57808 800 57928 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 200946 703200 201002 703800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 275006 200 275062 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 583200 374688 583800 374808 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 86958 703200 87014 703800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal3 s 200 190408 800 190528 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 200 119688 800 119808 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235722 200 235778 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 275650 703200 275706 703800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 200 534488 800 534608 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 200 493008 800 493128 6 la_data_in[34]
port 199 nsew signal input
rlabel metal3 s 583200 245488 583800 245608 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 510710 200 510766 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 290462 200 290518 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 4526 703200 4582 703800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal3 s 200 638528 800 638648 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 583200 386928 583800 387048 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 204810 703200 204866 703800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 102414 703200 102470 703800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal3 s 583200 270648 583800 270768 6 la_data_in[43]
port 209 nsew signal input
rlabel metal3 s 200 53728 800 53848 6 la_data_in[44]
port 210 nsew signal input
rlabel metal3 s 583200 416168 583800 416288 6 la_data_in[45]
port 211 nsew signal input
rlabel metal3 s 200 223728 800 223848 6 la_data_in[46]
port 212 nsew signal input
rlabel metal3 s 583200 436568 583800 436688 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 200 356328 800 356448 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 47674 703200 47730 703800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 408314 200 408370 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 573822 703200 573878 703800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 200 427048 800 427168 6 la_data_in[51]
port 218 nsew signal input
rlabel metal3 s 200 642608 800 642728 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 200 70048 800 70168 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 3882 200 3938 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal3 s 583200 478048 583800 478168 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 200 480768 800 480888 6 la_data_in[56]
port 223 nsew signal input
rlabel metal3 s 583200 631728 583800 631848 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 86314 200 86370 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal3 s 583200 411408 583800 411528 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 341982 703200 342038 703800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 518438 200 518494 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal3 s 583200 461728 583800 461848 6 la_data_in[61]
port 229 nsew signal input
rlabel metal3 s 583200 17688 583800 17808 6 la_data_in[62]
port 230 nsew signal input
rlabel metal3 s 583200 382848 583800 382968 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 361946 703200 362002 703800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal3 s 200 435208 800 435328 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 546774 703200 546830 703800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal3 s 200 352248 800 352368 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 200 501848 800 501968 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 583200 13608 583800 13728 6 la_data_in[69]
port 237 nsew signal input
rlabel metal3 s 583200 258408 583800 258528 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 583200 577328 583800 577448 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 583200 614728 583800 614848 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 436650 703200 436706 703800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal3 s 200 65968 800 66088 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 583200 282888 583800 283008 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 133970 703200 134026 703800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal3 s 583200 116968 583800 117088 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 491390 703200 491446 703800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 337474 200 337530 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 583200 565088 583800 565208 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 329746 200 329802 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal3 s 200 78208 800 78328 6 la_data_in[80]
port 250 nsew signal input
rlabel metal3 s 583200 38088 583800 38208 6 la_data_in[81]
port 251 nsew signal input
rlabel metal3 s 583200 303968 583800 304088 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 526810 703200 526866 703800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 553858 200 553914 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 173254 703200 173310 703800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal3 s 583200 407328 583800 407448 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 424414 703200 424470 703800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 149426 703200 149482 703800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 345846 703200 345902 703800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal3 s 200 335928 800 336048 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 541622 200 541678 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal3 s 200 381488 800 381608 6 la_data_in[91]
port 262 nsew signal input
rlabel metal3 s 583200 548768 583800 548888 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 232502 703200 232558 703800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 200 294448 800 294568 6 la_data_in[94]
port 265 nsew signal input
rlabel metal3 s 583200 648048 583800 648168 6 la_data_in[95]
port 266 nsew signal input
rlabel metal3 s 200 472608 800 472728 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 393502 703200 393558 703800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 270498 200 270554 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 200 514088 800 514208 6 la_data_in[99]
port 270 nsew signal input
rlabel metal3 s 583200 365848 583800 365968 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 334254 703200 334310 703800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal3 s 583200 428408 583800 428528 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 223486 200 223542 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 121734 200 121790 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 583200 221008 583800 221128 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 507490 703200 507546 703800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 583200 158448 583800 158568 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 148782 200 148838 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal3 s 583200 353608 583800 353728 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 583200 473968 583800 474088 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 416686 703200 416742 703800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 427634 200 427690 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 200 277448 800 277568 6 la_data_out[110]
port 284 nsew signal output
rlabel metal3 s 583200 195848 583800 195968 6 la_data_out[111]
port 285 nsew signal output
rlabel metal3 s 200 202648 800 202768 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 196438 200 196494 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 662 703200 718 703800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 583200 154368 583800 154488 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 396722 200 396778 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 19982 703200 20038 703800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal3 s 583200 361768 583800 361888 6 la_data_out[118]
port 292 nsew signal output
rlabel metal3 s 583200 5448 583800 5568 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 583200 249568 583800 249688 6 la_data_out[11]
port 294 nsew signal output
rlabel metal3 s 200 148928 800 149048 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 255042 200 255098 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 200 28568 800 28688 6 la_data_out[122]
port 297 nsew signal output
rlabel metal3 s 583200 643968 583800 644088 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 534538 703200 534594 703800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal3 s 200 667768 800 667888 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 74722 703200 74778 703800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 59266 703200 59322 703800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 219622 200 219678 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal3 s 583200 21768 583800 21888 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 200 613368 800 613488 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 200 468528 800 468648 6 la_data_out[15]
port 306 nsew signal output
rlabel metal3 s 583200 444728 583800 444848 6 la_data_out[16]
port 307 nsew signal output
rlabel metal3 s 583200 399168 583800 399288 6 la_data_out[17]
port 308 nsew signal output
rlabel metal3 s 200 182248 800 182368 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 66994 703200 67050 703800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal3 s 583200 71408 583800 71528 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 294970 703200 295026 703800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal3 s 583200 204008 583800 204128 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 200 539248 800 539368 6 la_data_out[22]
port 314 nsew signal output
rlabel metal3 s 583200 208088 583800 208208 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 580906 200 580962 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 511354 703200 511410 703800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 200 377408 800 377528 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 90822 703200 90878 703800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 302054 200 302110 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 298190 200 298246 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 466918 200 466974 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 287242 703200 287298 703800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 200 244128 800 244248 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 200 298528 800 298648 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 350354 703200 350410 703800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 309782 200 309838 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 583200 133968 583800 134088 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 51538 703200 51594 703800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 577042 200 577098 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal3 s 583200 55088 583800 55208 6 la_data_out[38]
port 331 nsew signal output
rlabel metal3 s 583200 112888 583800 113008 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 188710 703200 188766 703800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal3 s 583200 324368 583800 324488 6 la_data_out[40]
port 334 nsew signal output
rlabel metal3 s 200 95208 800 95328 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 200 680008 800 680128 6 la_data_out[42]
port 336 nsew signal output
rlabel metal3 s 200 61888 800 62008 6 la_data_out[43]
port 337 nsew signal output
rlabel metal3 s 200 331848 800 331968 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 369030 200 369086 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 106278 703200 106334 703800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 66350 200 66406 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 291106 703200 291162 703800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 200 650768 800 650888 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 519082 703200 519138 703800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 200 248888 800 249008 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 361302 200 361358 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 200 87048 800 87168 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 389638 703200 389694 703800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 200 410048 800 410168 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 200302 200 200358 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 412178 200 412234 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 197082 703200 197138 703800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 39946 703200 40002 703800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 200 327088 800 327208 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 349066 200 349122 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 341338 200 341394 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 487526 703200 487582 703800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 200 124448 800 124568 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 468206 703200 468262 703800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 200 418888 800 419008 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 514574 200 514630 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 573178 200 573234 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 583200 440648 583800 440768 6 la_data_out[67]
port 363 nsew signal output
rlabel metal3 s 583200 225088 583800 225208 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 98550 703200 98606 703800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 314290 200 314346 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 463054 200 463110 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 239586 200 239642 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal3 s 200 622208 800 622328 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 353574 200 353630 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 490746 200 490802 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 392858 200 392914 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 172610 200 172666 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 31574 703200 31630 703800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 325882 200 325938 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal3 s 200 103368 800 103488 6 la_data_out[79]
port 376 nsew signal output
rlabel metal3 s 583200 34008 583800 34128 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 583200 216928 583800 217048 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 110142 703200 110198 703800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal3 s 200 49648 800 49768 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 200 575968 800 576088 6 la_data_out[83]
port 381 nsew signal output
rlabel metal3 s 200 219648 800 219768 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 542266 703200 542322 703800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 530030 200 530086 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 583200 685448 583800 685568 6 la_data_out[87]
port 385 nsew signal output
rlabel metal3 s 200 115608 800 115728 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 583200 67328 583800 67448 6 la_data_out[89]
port 387 nsew signal output
rlabel metal3 s 583200 424328 583800 424448 6 la_data_out[8]
port 388 nsew signal output
rlabel metal3 s 200 559648 800 559768 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 161662 703200 161718 703800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 236366 703200 236422 703800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal3 s 200 626288 800 626408 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 486882 200 486938 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 549994 200 550050 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 267278 703200 267334 703800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 188066 200 188122 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 577686 703200 577742 703800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 200 314848 800 314968 6 la_data_out[99]
port 398 nsew signal output
rlabel metal3 s 200 285608 800 285728 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 448242 703200 448298 703800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 432786 703200 432842 703800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 583200 75488 583800 75608 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 294326 200 294382 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal3 s 200 663688 800 663808 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 558366 703200 558422 703800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 583200 150288 583800 150408 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 444378 703200 444434 703800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 168746 200 168802 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal3 s 200 153008 800 153128 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 475290 200 475346 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 530674 703200 530730 703800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal3 s 200 518168 800 518288 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 200 584808 800 584928 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 405094 703200 405150 703800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 258906 200 258962 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 583200 582088 583800 582208 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 471426 200 471482 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 583200 420248 583800 420368 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 125598 200 125654 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 283378 703200 283434 703800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 376758 200 376814 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 333610 200 333666 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal3 s 200 290368 800 290488 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 583200 328448 583800 328568 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 200 696328 800 696448 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 583200 448808 583800 448928 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 70858 703200 70914 703800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 231214 200 231270 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 306562 703200 306618 703800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal3 s 200 227808 800 227928 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 583200 291728 583800 291848 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 583200 391008 583800 391128 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 533894 200 533950 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 583200 237328 583800 237448 6 la_oenb[15]
port 434 nsew signal input
rlabel metal3 s 583200 527688 583800 527808 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 302698 703200 302754 703800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 200 157088 800 157208 6 la_oenb[18]
port 437 nsew signal input
rlabel metal3 s 200 74128 800 74248 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 184202 200 184258 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 583200 183608 583800 183728 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 43166 200 43222 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 191930 200 191986 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal3 s 583200 166608 583800 166728 6 la_oenb[23]
port 443 nsew signal input
rlabel metal3 s 583200 689528 583800 689648 6 la_oenb[24]
port 444 nsew signal input
rlabel metal3 s 583200 345448 583800 345568 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 70214 200 70270 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal3 s 583200 295808 583800 295928 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 447598 200 447654 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 475934 703200 475990 703800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 416042 200 416098 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal3 s 583200 432488 583800 432608 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 554502 703200 554558 703800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 200 235968 800 236088 6 la_oenb[32]
port 453 nsew signal input
rlabel metal3 s 200 505928 800 506048 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 562230 703200 562286 703800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal3 s 200 99288 800 99408 6 la_oenb[35]
port 456 nsew signal input
rlabel metal3 s 200 310768 800 310888 6 la_oenb[36]
port 457 nsew signal input
rlabel metal3 s 583200 108808 583800 108928 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 200 194488 800 194608 6 la_oenb[38]
port 459 nsew signal input
rlabel metal3 s 200 265208 800 265328 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 227994 703200 228050 703800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 494610 200 494666 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal3 s 200 401888 800 402008 6 la_oenb[41]
port 463 nsew signal input
rlabel metal3 s 200 344088 800 344208 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 200 340008 800 340128 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 583200 669128 583800 669248 6 la_oenb[44]
port 466 nsew signal input
rlabel metal3 s 583200 9528 583800 9648 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 200 165928 800 166048 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 569314 200 569370 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal3 s 200 161168 800 161288 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 113362 200 113418 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 176474 200 176530 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 583200 29928 583800 30048 6 la_oenb[50]
port 473 nsew signal input
rlabel metal3 s 583200 266568 583800 266688 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 583200 610648 583800 610768 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 247958 703200 248014 703800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 220266 703200 220322 703800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 200 497768 800 497888 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 215758 200 215814 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 583200 677288 583800 677408 6 la_oenb[57]
port 480 nsew signal input
rlabel metal3 s 200 302608 800 302728 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 83094 703200 83150 703800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 137190 200 137246 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal3 s 583200 598408 583800 598528 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 200 132608 800 132728 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 326526 703200 326582 703800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 440514 703200 440570 703800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 472070 703200 472126 703800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 479798 703200 479854 703800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal3 s 200 45568 800 45688 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 263414 703200 263470 703800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 23202 200 23258 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 7746 200 7802 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 565450 200 565506 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal3 s 200 107448 800 107568 6 la_oenb[70]
port 495 nsew signal input
rlabel metal3 s 583200 191768 583800 191888 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 200 456288 800 456408 6 la_oenb[72]
port 497 nsew signal input
rlabel metal3 s 200 439288 800 439408 6 la_oenb[73]
port 498 nsew signal input
rlabel metal3 s 200 530408 800 530528 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 200 273368 800 273488 6 la_oenb[75]
port 500 nsew signal input
rlabel metal3 s 200 231888 800 232008 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 200 178168 800 178288 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 251822 703200 251878 703800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 583200 688 583800 808 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 278870 200 278926 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 200 510008 800 510128 6 la_oenb[80]
port 506 nsew signal input
rlabel metal3 s 583200 523608 583800 523728 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 583200 660288 583800 660408 6 la_oenb[82]
port 508 nsew signal input
rlabel metal3 s 200 368568 800 368688 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 200 24488 800 24608 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 583200 138048 583800 138168 6 la_oenb[85]
port 511 nsew signal input
rlabel metal3 s 583200 627648 583800 627768 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 165526 703200 165582 703800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 583200 531768 583800 531888 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 545486 200 545542 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 322662 703200 322718 703800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal3 s 583200 212848 583800 212968 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 118514 703200 118570 703800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal3 s 583200 79568 583800 79688 6 la_oenb[92]
port 519 nsew signal input
rlabel metal3 s 200 571888 800 572008 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 90178 200 90234 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 583200 507288 583800 507408 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 400586 200 400642 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 583200 618808 583800 618928 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 180338 200 180394 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal3 s 583200 92488 583800 92608 6 la_oenb[99]
port 526 nsew signal input
rlabel metal3 s 200 630368 800 630488 6 la_oenb[9]
port 527 nsew signal input
rlabel metal3 s 200 318928 800 319048 6 user_clock2
port 528 nsew signal input
rlabel metal3 s 200 144848 800 144968 6 user_irq[0]
port 529 nsew signal output
rlabel metal3 s 200 605208 800 605328 6 user_irq[1]
port 530 nsew signal output
rlabel metal3 s 200 671848 800 671968 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -416 656 -96 703280 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -416 656 584340 976 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -416 702960 584340 703280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 584020 656 584340 703280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 8344 -3964 8664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 22344 -3964 22664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 22344 646209 22664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 36344 -3964 36664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 36344 646209 36664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 50344 -3964 50664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 50344 646209 50664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 64344 -3964 64664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 64344 646209 64664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 78344 -3964 78664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 78344 646209 78664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 92344 -3964 92664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 92344 646209 92664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 106344 -3964 106664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 106344 646209 106664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 120344 -3964 120664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 120344 646209 120664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 134344 -3964 134664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 134344 646209 134664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148344 -3964 148664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148344 646209 148664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 162344 -3964 162664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 162344 646209 162664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 176344 -3964 176664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 176344 646209 176664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 190344 -3964 190664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 190344 646209 190664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 204344 -3964 204664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 204344 646209 204664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 218344 -3964 218664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 218344 646209 218664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 232344 -3964 232664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 232344 646209 232664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 246344 -3964 246664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 246344 646209 246664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 260344 -3964 260664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 260344 646209 260664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 274344 -3964 274664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 274344 646209 274664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 288344 -3964 288664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 288344 646209 288664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 302344 -3964 302664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 302344 646209 302664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 316344 -3964 316664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 316344 646209 316664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 330344 -3964 330664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 330344 646209 330664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 344344 -3964 344664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 344344 646209 344664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 358344 -3964 358664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 358344 646209 358664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 372344 -3964 372664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 372344 646209 372664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 386344 -3964 386664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 386344 646209 386664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400344 -3964 400664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400344 646209 400664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 414344 -3964 414664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 414344 646209 414664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 428344 -3964 428664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 428344 646209 428664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442344 -3964 442664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442344 646209 442664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 456344 -3964 456664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 456344 646209 456664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 470344 -3964 470664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 470344 646209 470664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 484344 -3964 484664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 484344 646209 484664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 498344 -3964 498664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 498344 646209 498664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 512344 -3964 512664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 512344 646209 512664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 526344 -3964 526664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 526344 646209 526664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 540344 -3964 540664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 540344 646209 540664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 554344 -3964 554664 56679 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 554344 646209 554664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 568344 -3964 568664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 582344 -3964 582664 707900 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 9416 588960 9736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 24416 588960 24736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 39416 588960 39736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 54416 588960 54736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 69416 588960 69736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 84416 588960 84736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 99416 588960 99736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 114416 588960 114736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 129416 588960 129736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 144416 588960 144736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 159416 588960 159736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 174416 588960 174736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 189416 588960 189736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 204416 588960 204736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 219416 588960 219736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 234416 588960 234736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 249416 588960 249736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 264416 588960 264736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 279416 588960 279736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 294416 588960 294736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 309416 588960 309736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 324416 588960 324736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 339416 588960 339736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 354416 588960 354736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 369416 588960 369736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 384416 588960 384736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 399416 588960 399736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 414416 588960 414736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 429416 588960 429736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 444416 588960 444736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 459416 588960 459736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 474416 588960 474736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 489416 588960 489736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 504416 588960 504736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 519416 588960 519736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 534416 588960 534736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 549416 588960 549736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 564416 588960 564736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 579416 588960 579736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 594416 588960 594736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 609416 588960 609736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 624416 588960 624736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 639416 588960 639736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 654416 588960 654736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 669416 588960 669736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 684416 588960 684736 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -5036 699416 588960 699736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -1736 -664 -1416 704600 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -1736 -664 585660 -344 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -1736 704280 585660 704600 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 585340 -664 585660 704600 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 9664 -3964 9984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 23664 -3964 23984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 23664 646209 23984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 37664 -3964 37984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 37664 646209 37984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 51664 -3964 51984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 51664 646209 51984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 65664 -3964 65984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 65664 646209 65984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 79664 -3964 79984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 79664 646209 79984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 93664 -3964 93984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 93664 646209 93984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 107664 -3964 107984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 107664 646209 107984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 121664 -3964 121984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 121664 646209 121984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 135664 -3964 135984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 135664 646209 135984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149664 -3964 149984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149664 646209 149984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 163664 -3964 163984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 163664 646209 163984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 177664 -3964 177984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 177664 646209 177984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 191664 -3964 191984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 191664 646209 191984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 205664 -3964 205984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 205664 646209 205984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219664 -3964 219984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219664 646209 219984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 233664 -3964 233984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 233664 646209 233984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 247664 -3964 247984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 247664 646209 247984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 261664 -3964 261984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 261664 646209 261984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 275664 -3964 275984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 275664 646209 275984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 289664 -3964 289984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 289664 646209 289984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 303664 -3964 303984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 303664 646209 303984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 317664 -3964 317984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 317664 646209 317984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 331664 -3964 331984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 331664 646209 331984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 345664 -3964 345984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 345664 646209 345984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 359664 -3964 359984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 359664 646209 359984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 373664 -3964 373984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 373664 646209 373984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 387664 -3964 387984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 387664 646209 387984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401664 -3964 401984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401664 646209 401984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 415664 -3964 415984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 415664 646209 415984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 429664 -3964 429984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 429664 646209 429984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 443664 -3964 443984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 443664 646209 443984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 457664 -3964 457984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 457664 646209 457984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 471664 -3964 471984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 471664 646209 471984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 485664 -3964 485984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 485664 646209 485984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 499664 -3964 499984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 499664 646209 499984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 513664 -3964 513984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 513664 646209 513984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 527664 -3964 527984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 527664 646209 527984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 541664 -3964 541984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 541664 646209 541984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 555664 -3964 555984 56679 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 555664 646209 555984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 569664 -3964 569984 208100 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 569664 257468 569984 309828 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 569664 359740 569984 412100 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 569664 461468 569984 513828 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 569664 563740 569984 707900 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 10736 588960 11056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 25736 588960 26056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 40736 588960 41056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 55736 588960 56056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 70736 588960 71056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 85736 588960 86056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 100736 588960 101056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 115736 588960 116056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 130736 588960 131056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 145736 588960 146056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 160736 588960 161056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 175736 588960 176056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 190736 588960 191056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 205736 588960 206056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 220736 588960 221056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 235736 588960 236056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 250736 588960 251056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 265736 588960 266056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 280736 588960 281056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 295736 588960 296056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 310736 588960 311056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 325736 588960 326056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 340736 588960 341056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 355736 588960 356056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 370736 588960 371056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 385736 588960 386056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 400736 588960 401056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 415736 588960 416056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 430736 588960 431056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 445736 588960 446056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 460736 588960 461056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 475736 588960 476056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 490736 588960 491056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 505736 588960 506056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 520736 588960 521056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 535736 588960 536056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 550736 588960 551056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 565736 588960 566056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 580736 588960 581056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 595736 588960 596056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 610736 588960 611056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 625736 588960 626056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 640736 588960 641056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 655736 588960 656056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 670736 588960 671056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 685736 588960 686056 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -5036 700736 588960 701056 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -3056 -1984 -2736 705920 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -3056 -1984 586980 -1664 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -3056 705600 586980 705920 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 586660 -1984 586980 705920 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 10984 -3964 11304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 24984 -3964 25304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 24984 646209 25304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 38984 -3964 39304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 38984 646209 39304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 52984 -3964 53304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 52984 646209 53304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 66984 -3964 67304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 66984 646209 67304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 80984 -3964 81304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 80984 646209 81304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 94984 -3964 95304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 94984 646209 95304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 108984 -3964 109304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 108984 646209 109304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 122984 -3964 123304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 122984 646209 123304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136984 -3964 137304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136984 646209 137304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 150984 -3964 151304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 150984 646209 151304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 164984 -3964 165304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 164984 646209 165304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 178984 -3964 179304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 178984 646209 179304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 192984 -3964 193304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 192984 646209 193304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 206984 -3964 207304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 206984 646209 207304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 220984 -3964 221304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 220984 646209 221304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 234984 -3964 235304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 234984 646209 235304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 248984 -3964 249304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 248984 646209 249304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 262984 -3964 263304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 262984 646209 263304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 276984 -3964 277304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 276984 646209 277304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 290984 -3964 291304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 290984 646209 291304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 304984 -3964 305304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 304984 646209 305304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 318984 -3964 319304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 318984 646209 319304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 332984 -3964 333304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 332984 646209 333304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 346984 -3964 347304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 346984 646209 347304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 360984 -3964 361304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 360984 646209 361304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 374984 -3964 375304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 374984 646209 375304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 388984 -3964 389304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 388984 646209 389304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 402984 -3964 403304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 402984 646209 403304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 416984 -3964 417304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 416984 646209 417304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 430984 -3964 431304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 430984 646209 431304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 444984 -3964 445304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 444984 646209 445304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 458984 -3964 459304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 458984 646209 459304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 472984 -3964 473304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 472984 646209 473304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 486984 -3964 487304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 486984 646209 487304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 500984 -3964 501304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 500984 646209 501304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 514984 -3964 515304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 514984 646209 515304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 528984 -3964 529304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 528984 646209 529304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 542984 -3964 543304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 542984 646209 543304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556984 -3964 557304 56679 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556984 646209 557304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 570984 -3964 571304 707900 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 12056 588960 12376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 27056 588960 27376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 42056 588960 42376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 57056 588960 57376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 72056 588960 72376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 87056 588960 87376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 102056 588960 102376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 117056 588960 117376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 132056 588960 132376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 147056 588960 147376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 162056 588960 162376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 177056 588960 177376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 192056 588960 192376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 207056 465010 207376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 222056 588960 222376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 237056 588960 237376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 252056 588960 252376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 267056 588960 267376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 282056 588960 282376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 297056 588960 297376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 312056 588960 312376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 327056 588960 327376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 342056 588960 342376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 357056 588960 357376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 372056 588960 372376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 387056 588960 387376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 402056 588960 402376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 417056 588960 417376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 432056 588960 432376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 447056 588960 447376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 462056 588960 462376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 477056 588960 477376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 492056 588960 492376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 507056 588960 507376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 522056 588960 522376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 537056 588960 537376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 552056 588960 552376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 567056 588960 567376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 582056 588960 582376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 597056 588960 597376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 612056 588960 612376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 627056 588960 627376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 642056 588960 642376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 657056 588960 657376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 672056 588960 672376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5036 687056 588960 687376 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 498630 207056 588960 207376 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -4376 -3304 -4056 707240 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4376 -3304 588300 -2984 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -4376 706920 588300 707240 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 587980 -3304 588300 707240 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 12304 -3964 12624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 26304 -3964 26624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 26304 646209 26624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 40304 -3964 40624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 40304 646209 40624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54304 -3964 54624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54304 646209 54624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 68304 -3964 68624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 68304 646209 68624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 82304 -3964 82624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 82304 646209 82624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96304 -3964 96624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96304 646209 96624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 110304 -3964 110624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 110304 646209 110624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 124304 -3964 124624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 124304 646209 124624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 138304 -3964 138624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 138304 646209 138624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 152304 -3964 152624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 152304 646209 152624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 166304 -3964 166624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 166304 646209 166624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 180304 -3964 180624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 180304 646209 180624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 194304 -3964 194624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 194304 646209 194624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 208304 -3964 208624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 208304 646209 208624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 222304 -3964 222624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 222304 646209 222624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 236304 -3964 236624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 236304 646209 236624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 250304 -3964 250624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 250304 646209 250624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 264304 -3964 264624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 264304 646209 264624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 278304 -3964 278624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 278304 646209 278624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 292304 -3964 292624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 292304 646209 292624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 306304 -3964 306624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 306304 646209 306624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 320304 -3964 320624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 320304 646209 320624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 334304 -3964 334624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 334304 646209 334624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 348304 -3964 348624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 348304 646209 348624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 362304 -3964 362624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 362304 646209 362624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 376304 -3964 376624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 376304 646209 376624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 390304 -3964 390624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 390304 646209 390624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 404304 -3964 404624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 404304 646209 404624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 418304 -3964 418624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 418304 646209 418624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 432304 -3964 432624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 432304 646209 432624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 446304 -3964 446624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 446304 646209 446624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 460304 -3964 460624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 460304 646209 460624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474304 -3964 474624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474304 646209 474624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 488304 -3964 488624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 488304 646209 488624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 502304 -3964 502624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 502304 646209 502624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 516304 -3964 516624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 516304 646209 516624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 530304 -3964 530624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 530304 646209 530624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 544304 -3964 544624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 544304 646209 544624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 558304 -3964 558624 56679 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 558304 646209 558624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 572304 -3964 572624 707900 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 13376 588960 13696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 28376 588960 28696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 43376 588960 43696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 58376 588960 58696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 73376 588960 73696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 88376 588960 88696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 103376 588960 103696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 118376 588960 118696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 133376 588960 133696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 148376 588960 148696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 163376 588960 163696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 178376 588960 178696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 193376 588960 193696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 208376 588960 208696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 223376 588960 223696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 238376 588960 238696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 253376 588960 253696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 268376 588960 268696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 283376 588960 283696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 298376 588960 298696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 313376 588960 313696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 328376 588960 328696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 343376 588960 343696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 358376 588960 358696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 373376 588960 373696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 388376 588960 388696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 403376 588960 403696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 418376 588960 418696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 433376 588960 433696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 448376 588960 448696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 463376 588960 463696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 478376 588960 478696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 493376 588960 493696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 508376 588960 508696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 523376 588960 523696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 538376 588960 538696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 553376 588960 553696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 568376 588960 568696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 583376 588960 583696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 598376 588960 598696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 613376 588960 613696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 628376 588960 628696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 643376 588960 643696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 658376 588960 658696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 673376 588960 673696 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -5036 688376 588960 688696 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -3716 -2644 -3396 706580 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -3716 -2644 587640 -2324 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -3716 706260 587640 706580 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 587320 -2644 587640 706580 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 11644 -3964 11964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 25644 -3964 25964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 25644 646209 25964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 39644 -3964 39964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 39644 646209 39964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 53644 -3964 53964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 53644 646209 53964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 67644 -3964 67964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 67644 646209 67964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 81644 -3964 81964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 81644 646209 81964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 95644 -3964 95964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 95644 646209 95964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 109644 -3964 109964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 109644 646209 109964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 123644 -3964 123964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 123644 646209 123964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 137644 -3964 137964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 137644 646209 137964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 151644 -3964 151964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 151644 646209 151964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 165644 -3964 165964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 165644 646209 165964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 179644 -3964 179964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 179644 646209 179964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 193644 -3964 193964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 193644 646209 193964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 207644 -3964 207964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 207644 646209 207964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 221644 -3964 221964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 221644 646209 221964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 235644 -3964 235964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 235644 646209 235964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 249644 -3964 249964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 249644 646209 249964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 263644 -3964 263964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 263644 646209 263964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 277644 -3964 277964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 277644 646209 277964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 291644 -3964 291964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 291644 646209 291964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 305644 -3964 305964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 305644 646209 305964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 319644 -3964 319964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 319644 646209 319964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 333644 -3964 333964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 333644 646209 333964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 347644 -3964 347964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 347644 646209 347964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 361644 -3964 361964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 361644 646209 361964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 375644 -3964 375964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 375644 646209 375964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 389644 -3964 389964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 389644 646209 389964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 403644 -3964 403964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 403644 646209 403964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 417644 -3964 417964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 417644 646209 417964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 431644 -3964 431964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 431644 646209 431964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 445644 -3964 445964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 445644 646209 445964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 459644 -3964 459964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 459644 646209 459964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 473644 -3964 473964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 473644 646209 473964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 487644 -3964 487964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 487644 646209 487964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 501644 -3964 501964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 501644 646209 501964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 515644 -3964 515964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 515644 646209 515964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 529644 -3964 529964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 529644 646209 529964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 543644 -3964 543964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 543644 646209 543964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 557644 -3964 557964 56679 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 557644 646209 557964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 571644 -3964 571964 707900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 12716 588960 13036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 27716 588960 28036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 42716 588960 43036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 57716 588960 58036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 72716 588960 73036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 87716 588960 88036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 102716 588960 103036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 117716 588960 118036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 132716 588960 133036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 147716 588960 148036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 162716 588960 163036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 177716 588960 178036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 192716 588960 193036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 207716 465010 208036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 222716 588960 223036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 237716 588960 238036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 252716 588960 253036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 267716 588960 268036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 282716 588960 283036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 297716 588960 298036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 312716 588960 313036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 327716 588960 328036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 342716 588960 343036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 357716 588960 358036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 372716 588960 373036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 387716 588960 388036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 402716 588960 403036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 417716 588960 418036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 432716 588960 433036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 447716 588960 448036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 462716 588960 463036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 477716 588960 478036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 492716 588960 493036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 507716 588960 508036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 522716 588960 523036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 537716 588960 538036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 552716 588960 553036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 567716 588960 568036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 582716 588960 583036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 597716 588960 598036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 612716 588960 613036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 627716 588960 628036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 642716 588960 643036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 657716 588960 658036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 672716 588960 673036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -5036 687716 588960 688036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 498630 207716 588960 208036 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -5036 -3964 -4716 707900 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 -3964 588960 -3644 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 707580 588960 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 588640 -3964 588960 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 12964 -3964 13284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 26964 -3964 27284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 26964 646209 27284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 40964 -3964 41284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 40964 646209 41284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 54964 -3964 55284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 54964 646209 55284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 68964 -3964 69284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 68964 646209 69284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 82964 -3964 83284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 82964 646209 83284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 96964 -3964 97284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 96964 646209 97284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 110964 -3964 111284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 110964 646209 111284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 124964 -3964 125284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 124964 646209 125284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 138964 -3964 139284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 138964 646209 139284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 152964 -3964 153284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 152964 646209 153284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 166964 -3964 167284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 166964 646209 167284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 180964 -3964 181284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 180964 646209 181284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 194964 -3964 195284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 194964 646209 195284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 208964 -3964 209284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 208964 646209 209284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 222964 -3964 223284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 222964 646209 223284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 236964 -3964 237284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 236964 646209 237284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 250964 -3964 251284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 250964 646209 251284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 264964 -3964 265284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 264964 646209 265284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 278964 -3964 279284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 278964 646209 279284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 292964 -3964 293284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 292964 646209 293284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 306964 -3964 307284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 306964 646209 307284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 320964 -3964 321284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 320964 646209 321284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 334964 -3964 335284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 334964 646209 335284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 348964 -3964 349284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 348964 646209 349284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 362964 -3964 363284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 362964 646209 363284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 376964 -3964 377284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 376964 646209 377284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 390964 -3964 391284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 390964 646209 391284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 404964 -3964 405284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 404964 646209 405284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 418964 -3964 419284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 418964 646209 419284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 432964 -3964 433284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 432964 646209 433284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 446964 -3964 447284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 446964 646209 447284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 460964 -3964 461284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 460964 646209 461284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 474964 -3964 475284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 474964 646209 475284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 488964 -3964 489284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 488964 646209 489284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 502964 -3964 503284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 502964 646209 503284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 516964 -3964 517284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 516964 646209 517284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 530964 -3964 531284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 530964 646209 531284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 544964 -3964 545284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 544964 646209 545284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 558964 -3964 559284 56679 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 558964 646209 559284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 572964 -3964 573284 707900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 14036 588960 14356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 29036 588960 29356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 44036 588960 44356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 59036 588960 59356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 74036 588960 74356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 89036 588960 89356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 104036 588960 104356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 119036 588960 119356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 134036 588960 134356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 149036 588960 149356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 164036 588960 164356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 179036 588960 179356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 194036 588960 194356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 209036 588960 209356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 224036 588960 224356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 239036 588960 239356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 254036 588960 254356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 269036 588960 269356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 284036 588960 284356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 299036 588960 299356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 314036 588960 314356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 329036 588960 329356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 344036 588960 344356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 359036 588960 359356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 374036 588960 374356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 389036 588960 389356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 404036 588960 404356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 419036 588960 419356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 434036 588960 434356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 449036 588960 449356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 464036 588960 464356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 479036 588960 479356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 494036 588960 494356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 509036 588960 509356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 524036 588960 524356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 539036 588960 539356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 554036 588960 554356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 569036 588960 569356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 584036 588960 584356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 599036 588960 599356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 614036 588960 614356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 629036 588960 629356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 644036 588960 644356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 659036 588960 659356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 674036 588960 674356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -5036 689036 588960 689356 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -1076 -4 -756 703940 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -1076 -4 585000 316 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -1076 703620 585000 703940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 584680 -4 585000 703940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 9004 -3964 9324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 23004 -3964 23324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 23004 646209 23324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 37004 -3964 37324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 37004 646209 37324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 51004 -3964 51324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 51004 646209 51324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65004 -3964 65324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65004 646209 65324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 79004 -3964 79324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 79004 646209 79324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 93004 -3964 93324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 93004 646209 93324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 107004 -3964 107324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 107004 646209 107324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 121004 -3964 121324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 121004 646209 121324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 135004 -3964 135324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 135004 646209 135324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149004 -3964 149324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149004 646209 149324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 163004 -3964 163324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 163004 646209 163324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 177004 -3964 177324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 177004 646209 177324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 191004 -3964 191324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 191004 646209 191324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 205004 -3964 205324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 205004 646209 205324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219004 -3964 219324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219004 646209 219324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 233004 -3964 233324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 233004 646209 233324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 247004 -3964 247324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 247004 646209 247324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 261004 -3964 261324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 261004 646209 261324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 275004 -3964 275324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 275004 646209 275324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 289004 -3964 289324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 289004 646209 289324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 303004 -3964 303324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 303004 646209 303324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 317004 -3964 317324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 317004 646209 317324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 331004 -3964 331324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 331004 646209 331324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 345004 -3964 345324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 345004 646209 345324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 359004 -3964 359324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 359004 646209 359324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 373004 -3964 373324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 373004 646209 373324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387004 -3964 387324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387004 646209 387324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401004 -3964 401324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401004 646209 401324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 415004 -3964 415324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 415004 646209 415324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 429004 -3964 429324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 429004 646209 429324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 443004 -3964 443324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 443004 646209 443324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 457004 -3964 457324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 457004 646209 457324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 471004 -3964 471324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 471004 646209 471324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485004 -3964 485324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485004 646209 485324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 499004 -3964 499324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 499004 646209 499324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 513004 -3964 513324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 513004 646209 513324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 527004 -3964 527324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 527004 646209 527324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 541004 -3964 541324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 541004 646209 541324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 555004 -3964 555324 56679 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 555004 646209 555324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 569004 -3964 569324 208100 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 569004 257468 569324 309828 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 569004 359740 569324 412100 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 569004 461468 569324 513828 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 569004 563740 569324 707900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 10076 588960 10396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 25076 588960 25396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 40076 588960 40396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 55076 588960 55396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 70076 588960 70396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 85076 588960 85396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 100076 588960 100396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 115076 588960 115396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 130076 588960 130396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 145076 588960 145396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 160076 588960 160396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 175076 588960 175396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 190076 588960 190396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 205076 588960 205396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 220076 588960 220396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 235076 588960 235396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 250076 588960 250396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 265076 588960 265396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 280076 588960 280396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 295076 588960 295396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 310076 588960 310396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 325076 588960 325396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 340076 588960 340396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 355076 588960 355396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 370076 588960 370396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 385076 588960 385396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 400076 588960 400396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 415076 588960 415396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 430076 588960 430396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 445076 588960 445396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 460076 588960 460396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 475076 588960 475396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 490076 588960 490396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 505076 588960 505396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 520076 588960 520396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 535076 588960 535396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 550076 588960 550396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 565076 588960 565396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 580076 588960 580396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 595076 588960 595396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 610076 588960 610396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 625076 588960 625396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 640076 588960 640396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 655076 588960 655396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 670076 588960 670396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 685076 588960 685396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -5036 700076 588960 700396 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 4900 54352 5220 649584 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 578612 54352 578932 649584 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -2396 -1324 -2076 705260 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -2396 -1324 586320 -1004 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -2396 704940 586320 705260 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 586000 -1324 586320 705260 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 10324 -3964 10644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 24324 -3964 24644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 24324 646209 24644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 38324 -3964 38644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 38324 646209 38644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 52324 -3964 52644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 52324 646209 52644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 66324 -3964 66644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 66324 646209 66644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 80324 -3964 80644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 80324 646209 80644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 94324 -3964 94644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 94324 646209 94644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 108324 -3964 108644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 108324 646209 108644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 122324 -3964 122644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 122324 646209 122644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 136324 -3964 136644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 136324 646209 136644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 150324 -3964 150644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 150324 646209 150644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 164324 -3964 164644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 164324 646209 164644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 178324 -3964 178644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 178324 646209 178644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192324 -3964 192644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192324 646209 192644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 206324 -3964 206644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 206324 646209 206644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 220324 -3964 220644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 220324 646209 220644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 234324 -3964 234644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 234324 646209 234644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 248324 -3964 248644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 248324 646209 248644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 262324 -3964 262644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 262324 646209 262644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 276324 -3964 276644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 276324 646209 276644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 290324 -3964 290644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 290324 646209 290644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 304324 -3964 304644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 304324 646209 304644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 318324 -3964 318644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 318324 646209 318644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 332324 -3964 332644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 332324 646209 332644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 346324 -3964 346644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 346324 646209 346644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 360324 -3964 360644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 360324 646209 360644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 374324 -3964 374644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 374324 646209 374644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 388324 -3964 388644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 388324 646209 388644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 402324 -3964 402644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 402324 646209 402644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 416324 -3964 416644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 416324 646209 416644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 430324 -3964 430644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 430324 646209 430644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444324 -3964 444644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444324 646209 444644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 458324 -3964 458644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 458324 646209 458644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 472324 -3964 472644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 472324 646209 472644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 486324 -3964 486644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 486324 646209 486644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 500324 -3964 500644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 500324 646209 500644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 514324 -3964 514644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 514324 646209 514644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 528324 -3964 528644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 528324 646209 528644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 542324 -3964 542644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 542324 646209 542644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 556324 -3964 556644 56679 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 556324 646209 556644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 570324 -3964 570644 707900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 11396 588960 11716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 26396 588960 26716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 41396 588960 41716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 56396 588960 56716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 71396 588960 71716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 86396 588960 86716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 101396 588960 101716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 116396 588960 116716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 131396 588960 131716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 146396 588960 146716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 161396 588960 161716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 176396 588960 176716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 191396 588960 191716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 206396 465010 206716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 221396 588960 221716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 236396 588960 236716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 251396 588960 251716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 266396 588960 266716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 281396 588960 281716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 296396 588960 296716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 311396 588960 311716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 326396 588960 326716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 341396 588960 341716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 356396 588960 356716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 371396 588960 371716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 386396 588960 386716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 401396 588960 401716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 416396 588960 416716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 431396 588960 431716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 446396 588960 446716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 461396 588960 461716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 476396 588960 476716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 491396 588960 491716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 506396 588960 506716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 521396 588960 521716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 536396 588960 536716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 551396 588960 551716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 566396 588960 566716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 581396 588960 581716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 596396 588960 596716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 611396 588960 611716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 626396 588960 626716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 641396 588960 641716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 656396 588960 656716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 671396 588960 671716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 686396 588960 686716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5036 701396 588960 701716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 498630 206396 588960 206716 6 vssd2
port 539 nsew ground bidirectional
rlabel metal3 s 583200 254328 583800 254448 6 wb_clk_i
port 540 nsew signal input
rlabel metal3 s 200 567808 800 567928 6 wb_rst_i
port 541 nsew signal input
rlabel metal3 s 583200 378768 583800 378888 6 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 208674 703200 208730 703800 6 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 63130 703200 63186 703800 6 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal3 s 200 484848 800 484968 6 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 62486 200 62542 800 6 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal3 s 200 373328 800 373448 6 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal3 s 583200 652128 583800 652248 6 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal3 s 583200 606568 583800 606688 6 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 439870 200 439926 800 6 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal3 s 583200 552848 583800 552968 6 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal3 s 583200 341368 583800 341488 6 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal3 s 583200 83648 583800 83768 6 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 216402 703200 216458 703800 6 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal3 s 200 215568 800 215688 6 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 388350 200 388406 800 6 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 557722 200 557778 800 6 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal3 s 583200 274728 583800 274848 6 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal3 s 200 563728 800 563848 6 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 372894 200 372950 800 6 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 74078 200 74134 800 6 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 23846 703200 23902 703800 6 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal3 s 583200 519528 583800 519648 6 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 502982 703200 503038 703800 6 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 262770 200 262826 800 6 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 338118 703200 338174 703800 6 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal3 s 583200 403248 583800 403368 6 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 526166 200 526222 800 6 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 330390 703200 330446 703800 6 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal3 s 200 111528 800 111648 6 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 211894 200 211950 800 6 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 34794 200 34850 800 6 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal3 s 583200 96568 583800 96688 6 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal3 s 583200 286968 583800 287088 6 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 35438 703200 35494 703800 6 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 581550 703200 581606 703800 6 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal3 s 200 364488 800 364608 6 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal3 s 200 414808 800 414928 6 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal3 s 200 397808 800 397928 6 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 27066 200 27122 800 6 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 144918 200 144974 800 6 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal3 s 583200 452888 583800 453008 6 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal3 s 200 36728 800 36848 6 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 298834 703200 298890 703800 6 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 459834 703200 459890 703800 6 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal3 s 200 580728 800 580848 6 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 101770 200 101826 800 6 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal3 s 583200 503208 583800 503328 6 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 483662 703200 483718 703800 6 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal3 s 200 269288 800 269408 6 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal3 s 583200 623568 583800 623688 6 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal3 s 583200 308048 583800 308168 6 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal3 s 200 16328 800 16448 6 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 412822 703200 412878 703800 6 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 27710 703200 27766 703800 6 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 208030 200 208086 800 6 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal3 s 583200 494368 583800 494488 6 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 537758 200 537814 800 6 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal3 s 583200 278808 583800 278928 6 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal3 s 200 252968 800 253088 6 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal3 s 583200 100648 583800 100768 6 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 105634 200 105690 800 6 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 322018 200 322074 800 6 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal3 s 200 4088 800 4208 6 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 401230 703200 401286 703800 6 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal3 s 583200 681368 583800 681488 6 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal3 s 583200 104728 583800 104848 6 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 50894 200 50950 800 6 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal3 s 583200 457648 583800 457768 6 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 15474 200 15530 800 6 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal3 s 583200 693608 583800 693728 6 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 385130 703200 385186 703800 6 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal3 s 583200 146208 583800 146328 6 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 365810 703200 365866 703800 6 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 436006 200 436062 800 6 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal3 s 200 12248 800 12368 6 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 432142 200 432198 800 6 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 18 200 74 800 6 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 506202 200 506258 800 6 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal3 s 200 261128 800 261248 6 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal3 s 200 526328 800 526448 6 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 94686 703200 94742 703800 6 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal3 s 200 170008 800 170128 6 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 133326 200 133382 800 6 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 47030 200 47086 800 6 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 255686 703200 255742 703800 6 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 114006 703200 114062 703800 6 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 345202 200 345258 800 6 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 369674 703200 369730 703800 6 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal3 s 583200 241408 583800 241528 6 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal3 s 200 405968 800 406088 6 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal3 s 583200 569168 583800 569288 6 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 141054 200 141110 800 6 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 243450 200 243506 800 6 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 380622 200 380678 800 6 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal3 s 583200 540608 583800 540728 6 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 384486 200 384542 800 6 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 358082 703200 358138 703800 6 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 354218 703200 354274 703800 6 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal3 s 200 601128 800 601248 6 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 16118 703200 16174 703800 6 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 455326 200 455382 800 6 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal3 s 200 140768 800 140888 6 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal3 s 200 543328 800 543448 6 wbs_stb_i
port 644 nsew signal input
rlabel metal3 s 583200 369928 583800 370048 6 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 122267766
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/user_project_wrapper/runs/23_01_01_14_20/results/signoff/user_project_wrapper.magic.gds
string GDS_START 95819546
<< end >>

